// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 12 2017 08:25:46

// File Generated:     Sep 12 2019 18:03:59

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "TinyFPGA_B" view "INTERFACE"

module TinyFPGA_B (
    USBPU,
    PIN_9,
    PIN_8,
    PIN_7,
    PIN_6,
    PIN_5,
    PIN_4,
    PIN_3,
    PIN_24,
    PIN_23,
    PIN_22,
    PIN_21,
    PIN_20,
    PIN_2,
    PIN_19,
    PIN_18,
    PIN_17,
    PIN_16,
    PIN_15,
    PIN_14,
    PIN_13,
    PIN_12,
    PIN_11,
    PIN_10,
    PIN_1,
    LED,
    CLK);

    output USBPU;
    input PIN_9;
    input PIN_8;
    input PIN_7;
    input PIN_6;
    input PIN_5;
    input PIN_4;
    inout PIN_3;
    input PIN_24;
    input PIN_23;
    input PIN_22;
    input PIN_21;
    input PIN_20;
    inout PIN_2;
    input PIN_19;
    input PIN_18;
    input PIN_17;
    input PIN_16;
    input PIN_15;
    input PIN_14;
    input PIN_13;
    input PIN_12;
    input PIN_11;
    input PIN_10;
    inout PIN_1;
    output LED;
    input CLK;

    wire N__50526;
    wire N__50525;
    wire N__50524;
    wire N__50517;
    wire N__50516;
    wire N__50515;
    wire N__50508;
    wire N__50507;
    wire N__50506;
    wire N__50499;
    wire N__50498;
    wire N__50497;
    wire N__50490;
    wire N__50489;
    wire N__50488;
    wire N__50481;
    wire N__50480;
    wire N__50479;
    wire N__50462;
    wire N__50459;
    wire N__50456;
    wire N__50453;
    wire N__50450;
    wire N__50447;
    wire N__50446;
    wire N__50443;
    wire N__50440;
    wire N__50435;
    wire N__50434;
    wire N__50433;
    wire N__50432;
    wire N__50431;
    wire N__50430;
    wire N__50429;
    wire N__50428;
    wire N__50427;
    wire N__50426;
    wire N__50425;
    wire N__50424;
    wire N__50423;
    wire N__50422;
    wire N__50421;
    wire N__50420;
    wire N__50419;
    wire N__50418;
    wire N__50417;
    wire N__50416;
    wire N__50415;
    wire N__50414;
    wire N__50413;
    wire N__50412;
    wire N__50411;
    wire N__50410;
    wire N__50409;
    wire N__50408;
    wire N__50407;
    wire N__50406;
    wire N__50405;
    wire N__50404;
    wire N__50403;
    wire N__50402;
    wire N__50401;
    wire N__50400;
    wire N__50399;
    wire N__50398;
    wire N__50397;
    wire N__50396;
    wire N__50395;
    wire N__50394;
    wire N__50393;
    wire N__50392;
    wire N__50391;
    wire N__50390;
    wire N__50389;
    wire N__50388;
    wire N__50387;
    wire N__50386;
    wire N__50385;
    wire N__50384;
    wire N__50383;
    wire N__50382;
    wire N__50381;
    wire N__50380;
    wire N__50379;
    wire N__50378;
    wire N__50377;
    wire N__50376;
    wire N__50375;
    wire N__50374;
    wire N__50373;
    wire N__50372;
    wire N__50371;
    wire N__50370;
    wire N__50369;
    wire N__50368;
    wire N__50367;
    wire N__50366;
    wire N__50365;
    wire N__50364;
    wire N__50363;
    wire N__50362;
    wire N__50361;
    wire N__50360;
    wire N__50359;
    wire N__50358;
    wire N__50357;
    wire N__50356;
    wire N__50355;
    wire N__50354;
    wire N__50353;
    wire N__50352;
    wire N__50351;
    wire N__50350;
    wire N__50349;
    wire N__50348;
    wire N__50347;
    wire N__50346;
    wire N__50345;
    wire N__50344;
    wire N__50343;
    wire N__50342;
    wire N__50341;
    wire N__50340;
    wire N__50339;
    wire N__50338;
    wire N__50337;
    wire N__50336;
    wire N__50335;
    wire N__50334;
    wire N__50333;
    wire N__50332;
    wire N__50331;
    wire N__50330;
    wire N__50329;
    wire N__50328;
    wire N__50327;
    wire N__50326;
    wire N__50325;
    wire N__50324;
    wire N__50323;
    wire N__50322;
    wire N__50321;
    wire N__50320;
    wire N__50319;
    wire N__50318;
    wire N__50317;
    wire N__50316;
    wire N__50315;
    wire N__50314;
    wire N__50313;
    wire N__50312;
    wire N__50311;
    wire N__50310;
    wire N__50309;
    wire N__50308;
    wire N__50307;
    wire N__50306;
    wire N__50305;
    wire N__50304;
    wire N__50303;
    wire N__50302;
    wire N__50301;
    wire N__50300;
    wire N__50299;
    wire N__50298;
    wire N__50297;
    wire N__50296;
    wire N__50295;
    wire N__50294;
    wire N__50293;
    wire N__50292;
    wire N__50291;
    wire N__50290;
    wire N__50289;
    wire N__50288;
    wire N__50287;
    wire N__50286;
    wire N__50285;
    wire N__50284;
    wire N__50283;
    wire N__50282;
    wire N__50281;
    wire N__50280;
    wire N__50279;
    wire N__50278;
    wire N__50277;
    wire N__50276;
    wire N__50275;
    wire N__50274;
    wire N__50273;
    wire N__50272;
    wire N__50271;
    wire N__50270;
    wire N__50269;
    wire N__50268;
    wire N__50267;
    wire N__50266;
    wire N__50265;
    wire N__50264;
    wire N__50263;
    wire N__50262;
    wire N__50261;
    wire N__50260;
    wire N__50259;
    wire N__50258;
    wire N__50257;
    wire N__50256;
    wire N__50255;
    wire N__50254;
    wire N__50253;
    wire N__50252;
    wire N__50251;
    wire N__49880;
    wire N__49877;
    wire N__49874;
    wire N__49873;
    wire N__49872;
    wire N__49869;
    wire N__49868;
    wire N__49867;
    wire N__49866;
    wire N__49863;
    wire N__49860;
    wire N__49857;
    wire N__49854;
    wire N__49853;
    wire N__49850;
    wire N__49847;
    wire N__49846;
    wire N__49843;
    wire N__49836;
    wire N__49833;
    wire N__49830;
    wire N__49827;
    wire N__49824;
    wire N__49819;
    wire N__49808;
    wire N__49807;
    wire N__49804;
    wire N__49801;
    wire N__49798;
    wire N__49793;
    wire N__49792;
    wire N__49791;
    wire N__49790;
    wire N__49787;
    wire N__49784;
    wire N__49783;
    wire N__49780;
    wire N__49777;
    wire N__49774;
    wire N__49771;
    wire N__49768;
    wire N__49763;
    wire N__49760;
    wire N__49755;
    wire N__49748;
    wire N__49745;
    wire N__49744;
    wire N__49741;
    wire N__49738;
    wire N__49733;
    wire N__49730;
    wire N__49727;
    wire N__49724;
    wire N__49721;
    wire N__49718;
    wire N__49715;
    wire N__49712;
    wire N__49709;
    wire N__49708;
    wire N__49707;
    wire N__49706;
    wire N__49703;
    wire N__49698;
    wire N__49697;
    wire N__49694;
    wire N__49691;
    wire N__49688;
    wire N__49685;
    wire N__49682;
    wire N__49679;
    wire N__49676;
    wire N__49667;
    wire N__49664;
    wire N__49663;
    wire N__49660;
    wire N__49657;
    wire N__49652;
    wire N__49651;
    wire N__49648;
    wire N__49645;
    wire N__49642;
    wire N__49637;
    wire N__49634;
    wire N__49633;
    wire N__49630;
    wire N__49627;
    wire N__49624;
    wire N__49621;
    wire N__49616;
    wire N__49615;
    wire N__49612;
    wire N__49611;
    wire N__49610;
    wire N__49607;
    wire N__49604;
    wire N__49603;
    wire N__49598;
    wire N__49595;
    wire N__49592;
    wire N__49589;
    wire N__49586;
    wire N__49581;
    wire N__49574;
    wire N__49571;
    wire N__49568;
    wire N__49567;
    wire N__49566;
    wire N__49565;
    wire N__49562;
    wire N__49555;
    wire N__49550;
    wire N__49549;
    wire N__49546;
    wire N__49543;
    wire N__49540;
    wire N__49537;
    wire N__49534;
    wire N__49531;
    wire N__49526;
    wire N__49523;
    wire N__49520;
    wire N__49519;
    wire N__49516;
    wire N__49513;
    wire N__49510;
    wire N__49505;
    wire N__49504;
    wire N__49501;
    wire N__49498;
    wire N__49493;
    wire N__49490;
    wire N__49487;
    wire N__49486;
    wire N__49483;
    wire N__49480;
    wire N__49477;
    wire N__49476;
    wire N__49473;
    wire N__49470;
    wire N__49467;
    wire N__49464;
    wire N__49461;
    wire N__49456;
    wire N__49451;
    wire N__49450;
    wire N__49449;
    wire N__49448;
    wire N__49447;
    wire N__49446;
    wire N__49445;
    wire N__49444;
    wire N__49443;
    wire N__49442;
    wire N__49437;
    wire N__49436;
    wire N__49435;
    wire N__49432;
    wire N__49427;
    wire N__49424;
    wire N__49423;
    wire N__49422;
    wire N__49421;
    wire N__49420;
    wire N__49419;
    wire N__49418;
    wire N__49417;
    wire N__49416;
    wire N__49415;
    wire N__49414;
    wire N__49411;
    wire N__49404;
    wire N__49401;
    wire N__49398;
    wire N__49397;
    wire N__49392;
    wire N__49389;
    wire N__49386;
    wire N__49385;
    wire N__49384;
    wire N__49383;
    wire N__49378;
    wire N__49371;
    wire N__49368;
    wire N__49365;
    wire N__49364;
    wire N__49363;
    wire N__49356;
    wire N__49353;
    wire N__49350;
    wire N__49347;
    wire N__49344;
    wire N__49341;
    wire N__49334;
    wire N__49329;
    wire N__49328;
    wire N__49327;
    wire N__49326;
    wire N__49325;
    wire N__49324;
    wire N__49323;
    wire N__49322;
    wire N__49321;
    wire N__49318;
    wire N__49309;
    wire N__49308;
    wire N__49305;
    wire N__49304;
    wire N__49301;
    wire N__49298;
    wire N__49295;
    wire N__49292;
    wire N__49291;
    wire N__49290;
    wire N__49289;
    wire N__49282;
    wire N__49277;
    wire N__49272;
    wire N__49267;
    wire N__49264;
    wire N__49257;
    wire N__49256;
    wire N__49255;
    wire N__49254;
    wire N__49253;
    wire N__49248;
    wire N__49245;
    wire N__49244;
    wire N__49237;
    wire N__49230;
    wire N__49223;
    wire N__49218;
    wire N__49209;
    wire N__49204;
    wire N__49199;
    wire N__49196;
    wire N__49191;
    wire N__49184;
    wire N__49181;
    wire N__49176;
    wire N__49163;
    wire N__49160;
    wire N__49157;
    wire N__49154;
    wire N__49151;
    wire N__49148;
    wire N__49145;
    wire N__49142;
    wire N__49139;
    wire N__49136;
    wire N__49133;
    wire N__49130;
    wire N__49127;
    wire N__49124;
    wire N__49121;
    wire N__49118;
    wire N__49115;
    wire N__49112;
    wire N__49111;
    wire N__49108;
    wire N__49103;
    wire N__49102;
    wire N__49099;
    wire N__49096;
    wire N__49091;
    wire N__49088;
    wire N__49087;
    wire N__49082;
    wire N__49079;
    wire N__49078;
    wire N__49075;
    wire N__49072;
    wire N__49067;
    wire N__49064;
    wire N__49063;
    wire N__49058;
    wire N__49057;
    wire N__49054;
    wire N__49051;
    wire N__49046;
    wire N__49043;
    wire N__49040;
    wire N__49039;
    wire N__49034;
    wire N__49031;
    wire N__49028;
    wire N__49025;
    wire N__49024;
    wire N__49021;
    wire N__49018;
    wire N__49013;
    wire N__49010;
    wire N__49007;
    wire N__49004;
    wire N__49001;
    wire N__48998;
    wire N__48995;
    wire N__48992;
    wire N__48989;
    wire N__48986;
    wire N__48983;
    wire N__48980;
    wire N__48977;
    wire N__48974;
    wire N__48971;
    wire N__48968;
    wire N__48965;
    wire N__48962;
    wire N__48959;
    wire N__48956;
    wire N__48953;
    wire N__48950;
    wire N__48947;
    wire N__48944;
    wire N__48941;
    wire N__48938;
    wire N__48935;
    wire N__48932;
    wire N__48929;
    wire N__48926;
    wire N__48923;
    wire N__48920;
    wire N__48917;
    wire N__48914;
    wire N__48911;
    wire N__48908;
    wire N__48905;
    wire N__48902;
    wire N__48899;
    wire N__48896;
    wire N__48893;
    wire N__48890;
    wire N__48887;
    wire N__48884;
    wire N__48881;
    wire N__48878;
    wire N__48875;
    wire N__48872;
    wire N__48869;
    wire N__48866;
    wire N__48863;
    wire N__48860;
    wire N__48857;
    wire N__48854;
    wire N__48851;
    wire N__48848;
    wire N__48845;
    wire N__48844;
    wire N__48841;
    wire N__48840;
    wire N__48839;
    wire N__48838;
    wire N__48837;
    wire N__48834;
    wire N__48833;
    wire N__48830;
    wire N__48825;
    wire N__48822;
    wire N__48819;
    wire N__48816;
    wire N__48815;
    wire N__48812;
    wire N__48811;
    wire N__48808;
    wire N__48805;
    wire N__48804;
    wire N__48801;
    wire N__48798;
    wire N__48795;
    wire N__48792;
    wire N__48787;
    wire N__48782;
    wire N__48779;
    wire N__48764;
    wire N__48761;
    wire N__48760;
    wire N__48759;
    wire N__48756;
    wire N__48755;
    wire N__48754;
    wire N__48751;
    wire N__48748;
    wire N__48745;
    wire N__48742;
    wire N__48739;
    wire N__48738;
    wire N__48737;
    wire N__48736;
    wire N__48733;
    wire N__48730;
    wire N__48725;
    wire N__48724;
    wire N__48721;
    wire N__48720;
    wire N__48717;
    wire N__48712;
    wire N__48705;
    wire N__48702;
    wire N__48699;
    wire N__48696;
    wire N__48683;
    wire N__48682;
    wire N__48679;
    wire N__48676;
    wire N__48675;
    wire N__48674;
    wire N__48671;
    wire N__48668;
    wire N__48665;
    wire N__48662;
    wire N__48661;
    wire N__48660;
    wire N__48657;
    wire N__48652;
    wire N__48649;
    wire N__48648;
    wire N__48643;
    wire N__48642;
    wire N__48635;
    wire N__48632;
    wire N__48629;
    wire N__48626;
    wire N__48617;
    wire N__48614;
    wire N__48611;
    wire N__48608;
    wire N__48607;
    wire N__48604;
    wire N__48601;
    wire N__48598;
    wire N__48593;
    wire N__48592;
    wire N__48591;
    wire N__48590;
    wire N__48589;
    wire N__48586;
    wire N__48583;
    wire N__48580;
    wire N__48577;
    wire N__48574;
    wire N__48571;
    wire N__48570;
    wire N__48569;
    wire N__48564;
    wire N__48561;
    wire N__48556;
    wire N__48553;
    wire N__48550;
    wire N__48547;
    wire N__48542;
    wire N__48533;
    wire N__48530;
    wire N__48527;
    wire N__48526;
    wire N__48523;
    wire N__48522;
    wire N__48519;
    wire N__48516;
    wire N__48513;
    wire N__48510;
    wire N__48507;
    wire N__48504;
    wire N__48503;
    wire N__48502;
    wire N__48501;
    wire N__48496;
    wire N__48493;
    wire N__48486;
    wire N__48479;
    wire N__48476;
    wire N__48473;
    wire N__48470;
    wire N__48469;
    wire N__48468;
    wire N__48467;
    wire N__48466;
    wire N__48465;
    wire N__48464;
    wire N__48463;
    wire N__48462;
    wire N__48461;
    wire N__48460;
    wire N__48459;
    wire N__48458;
    wire N__48457;
    wire N__48454;
    wire N__48447;
    wire N__48440;
    wire N__48433;
    wire N__48432;
    wire N__48431;
    wire N__48430;
    wire N__48429;
    wire N__48428;
    wire N__48427;
    wire N__48426;
    wire N__48425;
    wire N__48422;
    wire N__48421;
    wire N__48420;
    wire N__48419;
    wire N__48418;
    wire N__48417;
    wire N__48416;
    wire N__48415;
    wire N__48414;
    wire N__48413;
    wire N__48412;
    wire N__48411;
    wire N__48404;
    wire N__48403;
    wire N__48402;
    wire N__48401;
    wire N__48400;
    wire N__48399;
    wire N__48398;
    wire N__48397;
    wire N__48396;
    wire N__48395;
    wire N__48394;
    wire N__48385;
    wire N__48378;
    wire N__48377;
    wire N__48376;
    wire N__48373;
    wire N__48368;
    wire N__48365;
    wire N__48362;
    wire N__48359;
    wire N__48354;
    wire N__48349;
    wire N__48344;
    wire N__48333;
    wire N__48330;
    wire N__48325;
    wire N__48318;
    wire N__48315;
    wire N__48314;
    wire N__48313;
    wire N__48312;
    wire N__48307;
    wire N__48306;
    wire N__48303;
    wire N__48300;
    wire N__48295;
    wire N__48292;
    wire N__48289;
    wire N__48284;
    wire N__48281;
    wire N__48274;
    wire N__48261;
    wire N__48258;
    wire N__48255;
    wire N__48250;
    wire N__48247;
    wire N__48244;
    wire N__48237;
    wire N__48222;
    wire N__48209;
    wire N__48208;
    wire N__48205;
    wire N__48202;
    wire N__48199;
    wire N__48198;
    wire N__48195;
    wire N__48192;
    wire N__48189;
    wire N__48182;
    wire N__48179;
    wire N__48176;
    wire N__48173;
    wire N__48170;
    wire N__48167;
    wire N__48164;
    wire N__48163;
    wire N__48160;
    wire N__48159;
    wire N__48158;
    wire N__48157;
    wire N__48156;
    wire N__48155;
    wire N__48152;
    wire N__48151;
    wire N__48150;
    wire N__48149;
    wire N__48148;
    wire N__48145;
    wire N__48140;
    wire N__48137;
    wire N__48136;
    wire N__48135;
    wire N__48134;
    wire N__48133;
    wire N__48130;
    wire N__48129;
    wire N__48126;
    wire N__48123;
    wire N__48116;
    wire N__48113;
    wire N__48112;
    wire N__48111;
    wire N__48110;
    wire N__48109;
    wire N__48108;
    wire N__48107;
    wire N__48106;
    wire N__48103;
    wire N__48100;
    wire N__48097;
    wire N__48092;
    wire N__48089;
    wire N__48082;
    wire N__48081;
    wire N__48080;
    wire N__48077;
    wire N__48072;
    wire N__48069;
    wire N__48066;
    wire N__48061;
    wire N__48056;
    wire N__48051;
    wire N__48038;
    wire N__48033;
    wire N__48024;
    wire N__48021;
    wire N__48018;
    wire N__48013;
    wire N__48008;
    wire N__47999;
    wire N__47996;
    wire N__47993;
    wire N__47990;
    wire N__47987;
    wire N__47986;
    wire N__47985;
    wire N__47984;
    wire N__47983;
    wire N__47982;
    wire N__47981;
    wire N__47978;
    wire N__47975;
    wire N__47974;
    wire N__47973;
    wire N__47972;
    wire N__47971;
    wire N__47970;
    wire N__47969;
    wire N__47968;
    wire N__47967;
    wire N__47964;
    wire N__47961;
    wire N__47958;
    wire N__47957;
    wire N__47956;
    wire N__47953;
    wire N__47950;
    wire N__47947;
    wire N__47944;
    wire N__47941;
    wire N__47934;
    wire N__47931;
    wire N__47930;
    wire N__47927;
    wire N__47922;
    wire N__47919;
    wire N__47916;
    wire N__47913;
    wire N__47908;
    wire N__47903;
    wire N__47894;
    wire N__47891;
    wire N__47890;
    wire N__47887;
    wire N__47884;
    wire N__47881;
    wire N__47876;
    wire N__47871;
    wire N__47864;
    wire N__47861;
    wire N__47846;
    wire N__47843;
    wire N__47840;
    wire N__47837;
    wire N__47834;
    wire N__47833;
    wire N__47830;
    wire N__47827;
    wire N__47826;
    wire N__47825;
    wire N__47822;
    wire N__47819;
    wire N__47814;
    wire N__47807;
    wire N__47804;
    wire N__47801;
    wire N__47800;
    wire N__47799;
    wire N__47796;
    wire N__47793;
    wire N__47790;
    wire N__47783;
    wire N__47780;
    wire N__47779;
    wire N__47774;
    wire N__47771;
    wire N__47770;
    wire N__47769;
    wire N__47768;
    wire N__47767;
    wire N__47766;
    wire N__47763;
    wire N__47760;
    wire N__47757;
    wire N__47754;
    wire N__47753;
    wire N__47750;
    wire N__47747;
    wire N__47744;
    wire N__47741;
    wire N__47736;
    wire N__47733;
    wire N__47730;
    wire N__47723;
    wire N__47720;
    wire N__47711;
    wire N__47708;
    wire N__47705;
    wire N__47704;
    wire N__47703;
    wire N__47700;
    wire N__47697;
    wire N__47696;
    wire N__47695;
    wire N__47692;
    wire N__47687;
    wire N__47684;
    wire N__47681;
    wire N__47674;
    wire N__47671;
    wire N__47670;
    wire N__47669;
    wire N__47664;
    wire N__47661;
    wire N__47658;
    wire N__47655;
    wire N__47648;
    wire N__47645;
    wire N__47644;
    wire N__47641;
    wire N__47640;
    wire N__47637;
    wire N__47636;
    wire N__47635;
    wire N__47632;
    wire N__47629;
    wire N__47626;
    wire N__47623;
    wire N__47620;
    wire N__47619;
    wire N__47616;
    wire N__47613;
    wire N__47610;
    wire N__47605;
    wire N__47602;
    wire N__47599;
    wire N__47596;
    wire N__47591;
    wire N__47584;
    wire N__47579;
    wire N__47578;
    wire N__47577;
    wire N__47574;
    wire N__47571;
    wire N__47568;
    wire N__47565;
    wire N__47562;
    wire N__47561;
    wire N__47558;
    wire N__47553;
    wire N__47550;
    wire N__47547;
    wire N__47544;
    wire N__47537;
    wire N__47534;
    wire N__47533;
    wire N__47530;
    wire N__47529;
    wire N__47526;
    wire N__47523;
    wire N__47520;
    wire N__47513;
    wire N__47510;
    wire N__47507;
    wire N__47504;
    wire N__47501;
    wire N__47498;
    wire N__47495;
    wire N__47494;
    wire N__47489;
    wire N__47488;
    wire N__47485;
    wire N__47482;
    wire N__47477;
    wire N__47476;
    wire N__47473;
    wire N__47470;
    wire N__47465;
    wire N__47462;
    wire N__47461;
    wire N__47458;
    wire N__47455;
    wire N__47454;
    wire N__47453;
    wire N__47452;
    wire N__47451;
    wire N__47450;
    wire N__47449;
    wire N__47448;
    wire N__47447;
    wire N__47446;
    wire N__47445;
    wire N__47444;
    wire N__47443;
    wire N__47442;
    wire N__47441;
    wire N__47440;
    wire N__47439;
    wire N__47438;
    wire N__47437;
    wire N__47436;
    wire N__47435;
    wire N__47434;
    wire N__47431;
    wire N__47428;
    wire N__47421;
    wire N__47416;
    wire N__47415;
    wire N__47414;
    wire N__47413;
    wire N__47412;
    wire N__47411;
    wire N__47410;
    wire N__47409;
    wire N__47406;
    wire N__47405;
    wire N__47404;
    wire N__47403;
    wire N__47402;
    wire N__47401;
    wire N__47400;
    wire N__47399;
    wire N__47398;
    wire N__47397;
    wire N__47386;
    wire N__47375;
    wire N__47368;
    wire N__47363;
    wire N__47356;
    wire N__47353;
    wire N__47348;
    wire N__47343;
    wire N__47342;
    wire N__47341;
    wire N__47338;
    wire N__47333;
    wire N__47330;
    wire N__47327;
    wire N__47322;
    wire N__47317;
    wire N__47312;
    wire N__47307;
    wire N__47302;
    wire N__47301;
    wire N__47300;
    wire N__47299;
    wire N__47298;
    wire N__47297;
    wire N__47296;
    wire N__47295;
    wire N__47284;
    wire N__47283;
    wire N__47280;
    wire N__47277;
    wire N__47276;
    wire N__47275;
    wire N__47272;
    wire N__47259;
    wire N__47252;
    wire N__47243;
    wire N__47242;
    wire N__47241;
    wire N__47240;
    wire N__47237;
    wire N__47236;
    wire N__47235;
    wire N__47230;
    wire N__47229;
    wire N__47226;
    wire N__47223;
    wire N__47220;
    wire N__47217;
    wire N__47212;
    wire N__47203;
    wire N__47200;
    wire N__47197;
    wire N__47194;
    wire N__47191;
    wire N__47188;
    wire N__47185;
    wire N__47182;
    wire N__47179;
    wire N__47170;
    wire N__47163;
    wire N__47144;
    wire N__47143;
    wire N__47142;
    wire N__47141;
    wire N__47138;
    wire N__47137;
    wire N__47136;
    wire N__47135;
    wire N__47134;
    wire N__47131;
    wire N__47128;
    wire N__47127;
    wire N__47126;
    wire N__47123;
    wire N__47122;
    wire N__47119;
    wire N__47112;
    wire N__47111;
    wire N__47110;
    wire N__47107;
    wire N__47106;
    wire N__47103;
    wire N__47100;
    wire N__47097;
    wire N__47094;
    wire N__47089;
    wire N__47086;
    wire N__47083;
    wire N__47080;
    wire N__47079;
    wire N__47078;
    wire N__47077;
    wire N__47074;
    wire N__47071;
    wire N__47068;
    wire N__47065;
    wire N__47062;
    wire N__47059;
    wire N__47054;
    wire N__47049;
    wire N__47044;
    wire N__47041;
    wire N__47040;
    wire N__47039;
    wire N__47036;
    wire N__47033;
    wire N__47030;
    wire N__47027;
    wire N__47022;
    wire N__47019;
    wire N__47016;
    wire N__47011;
    wire N__47004;
    wire N__47001;
    wire N__46992;
    wire N__46979;
    wire N__46978;
    wire N__46977;
    wire N__46976;
    wire N__46973;
    wire N__46970;
    wire N__46965;
    wire N__46962;
    wire N__46955;
    wire N__46954;
    wire N__46951;
    wire N__46950;
    wire N__46949;
    wire N__46946;
    wire N__46943;
    wire N__46940;
    wire N__46937;
    wire N__46934;
    wire N__46931;
    wire N__46928;
    wire N__46919;
    wire N__46918;
    wire N__46917;
    wire N__46916;
    wire N__46915;
    wire N__46914;
    wire N__46911;
    wire N__46908;
    wire N__46907;
    wire N__46904;
    wire N__46903;
    wire N__46902;
    wire N__46901;
    wire N__46900;
    wire N__46899;
    wire N__46898;
    wire N__46897;
    wire N__46896;
    wire N__46895;
    wire N__46894;
    wire N__46893;
    wire N__46892;
    wire N__46891;
    wire N__46890;
    wire N__46889;
    wire N__46888;
    wire N__46885;
    wire N__46884;
    wire N__46883;
    wire N__46882;
    wire N__46881;
    wire N__46880;
    wire N__46879;
    wire N__46878;
    wire N__46877;
    wire N__46874;
    wire N__46873;
    wire N__46872;
    wire N__46871;
    wire N__46870;
    wire N__46869;
    wire N__46866;
    wire N__46863;
    wire N__46858;
    wire N__46855;
    wire N__46848;
    wire N__46845;
    wire N__46842;
    wire N__46837;
    wire N__46830;
    wire N__46825;
    wire N__46820;
    wire N__46815;
    wire N__46812;
    wire N__46805;
    wire N__46804;
    wire N__46801;
    wire N__46800;
    wire N__46799;
    wire N__46796;
    wire N__46795;
    wire N__46794;
    wire N__46793;
    wire N__46790;
    wire N__46789;
    wire N__46788;
    wire N__46787;
    wire N__46786;
    wire N__46785;
    wire N__46780;
    wire N__46773;
    wire N__46766;
    wire N__46759;
    wire N__46756;
    wire N__46753;
    wire N__46744;
    wire N__46733;
    wire N__46730;
    wire N__46725;
    wire N__46724;
    wire N__46723;
    wire N__46720;
    wire N__46717;
    wire N__46714;
    wire N__46711;
    wire N__46706;
    wire N__46703;
    wire N__46698;
    wire N__46697;
    wire N__46696;
    wire N__46695;
    wire N__46694;
    wire N__46691;
    wire N__46688;
    wire N__46673;
    wire N__46672;
    wire N__46671;
    wire N__46670;
    wire N__46667;
    wire N__46662;
    wire N__46657;
    wire N__46654;
    wire N__46647;
    wire N__46646;
    wire N__46645;
    wire N__46642;
    wire N__46637;
    wire N__46628;
    wire N__46627;
    wire N__46624;
    wire N__46621;
    wire N__46618;
    wire N__46611;
    wire N__46606;
    wire N__46599;
    wire N__46594;
    wire N__46587;
    wire N__46584;
    wire N__46565;
    wire N__46564;
    wire N__46561;
    wire N__46558;
    wire N__46557;
    wire N__46554;
    wire N__46551;
    wire N__46548;
    wire N__46547;
    wire N__46546;
    wire N__46539;
    wire N__46538;
    wire N__46535;
    wire N__46532;
    wire N__46531;
    wire N__46528;
    wire N__46525;
    wire N__46524;
    wire N__46523;
    wire N__46520;
    wire N__46517;
    wire N__46516;
    wire N__46513;
    wire N__46508;
    wire N__46503;
    wire N__46502;
    wire N__46499;
    wire N__46496;
    wire N__46493;
    wire N__46490;
    wire N__46485;
    wire N__46484;
    wire N__46481;
    wire N__46478;
    wire N__46475;
    wire N__46472;
    wire N__46467;
    wire N__46462;
    wire N__46451;
    wire N__46450;
    wire N__46449;
    wire N__46448;
    wire N__46447;
    wire N__46442;
    wire N__46441;
    wire N__46440;
    wire N__46435;
    wire N__46432;
    wire N__46429;
    wire N__46426;
    wire N__46423;
    wire N__46416;
    wire N__46413;
    wire N__46412;
    wire N__46409;
    wire N__46406;
    wire N__46403;
    wire N__46400;
    wire N__46397;
    wire N__46394;
    wire N__46391;
    wire N__46382;
    wire N__46379;
    wire N__46378;
    wire N__46375;
    wire N__46372;
    wire N__46367;
    wire N__46366;
    wire N__46365;
    wire N__46364;
    wire N__46361;
    wire N__46358;
    wire N__46355;
    wire N__46352;
    wire N__46349;
    wire N__46346;
    wire N__46343;
    wire N__46340;
    wire N__46335;
    wire N__46328;
    wire N__46325;
    wire N__46322;
    wire N__46319;
    wire N__46316;
    wire N__46313;
    wire N__46310;
    wire N__46309;
    wire N__46306;
    wire N__46303;
    wire N__46302;
    wire N__46297;
    wire N__46294;
    wire N__46291;
    wire N__46286;
    wire N__46283;
    wire N__46280;
    wire N__46279;
    wire N__46276;
    wire N__46275;
    wire N__46272;
    wire N__46269;
    wire N__46266;
    wire N__46261;
    wire N__46256;
    wire N__46255;
    wire N__46252;
    wire N__46249;
    wire N__46244;
    wire N__46241;
    wire N__46238;
    wire N__46235;
    wire N__46232;
    wire N__46229;
    wire N__46226;
    wire N__46223;
    wire N__46220;
    wire N__46219;
    wire N__46216;
    wire N__46213;
    wire N__46210;
    wire N__46207;
    wire N__46204;
    wire N__46199;
    wire N__46198;
    wire N__46195;
    wire N__46192;
    wire N__46189;
    wire N__46184;
    wire N__46183;
    wire N__46180;
    wire N__46177;
    wire N__46174;
    wire N__46169;
    wire N__46166;
    wire N__46163;
    wire N__46160;
    wire N__46157;
    wire N__46154;
    wire N__46151;
    wire N__46150;
    wire N__46149;
    wire N__46148;
    wire N__46143;
    wire N__46138;
    wire N__46135;
    wire N__46134;
    wire N__46131;
    wire N__46128;
    wire N__46125;
    wire N__46122;
    wire N__46119;
    wire N__46112;
    wire N__46109;
    wire N__46106;
    wire N__46105;
    wire N__46102;
    wire N__46099;
    wire N__46094;
    wire N__46091;
    wire N__46088;
    wire N__46087;
    wire N__46086;
    wire N__46083;
    wire N__46080;
    wire N__46079;
    wire N__46076;
    wire N__46073;
    wire N__46070;
    wire N__46067;
    wire N__46064;
    wire N__46057;
    wire N__46054;
    wire N__46049;
    wire N__46048;
    wire N__46047;
    wire N__46042;
    wire N__46041;
    wire N__46038;
    wire N__46037;
    wire N__46036;
    wire N__46035;
    wire N__46034;
    wire N__46033;
    wire N__46032;
    wire N__46031;
    wire N__46030;
    wire N__46029;
    wire N__46026;
    wire N__46023;
    wire N__46022;
    wire N__46019;
    wire N__46016;
    wire N__46015;
    wire N__46012;
    wire N__46009;
    wire N__46008;
    wire N__46005;
    wire N__46002;
    wire N__45995;
    wire N__45992;
    wire N__45987;
    wire N__45984;
    wire N__45981;
    wire N__45978;
    wire N__45975;
    wire N__45970;
    wire N__45967;
    wire N__45964;
    wire N__45959;
    wire N__45952;
    wire N__45949;
    wire N__45942;
    wire N__45939;
    wire N__45934;
    wire N__45931;
    wire N__45920;
    wire N__45917;
    wire N__45914;
    wire N__45913;
    wire N__45912;
    wire N__45911;
    wire N__45908;
    wire N__45905;
    wire N__45900;
    wire N__45899;
    wire N__45896;
    wire N__45891;
    wire N__45888;
    wire N__45883;
    wire N__45878;
    wire N__45875;
    wire N__45872;
    wire N__45869;
    wire N__45866;
    wire N__45863;
    wire N__45860;
    wire N__45857;
    wire N__45854;
    wire N__45851;
    wire N__45848;
    wire N__45845;
    wire N__45842;
    wire N__45839;
    wire N__45838;
    wire N__45835;
    wire N__45834;
    wire N__45831;
    wire N__45828;
    wire N__45825;
    wire N__45820;
    wire N__45817;
    wire N__45814;
    wire N__45811;
    wire N__45808;
    wire N__45803;
    wire N__45800;
    wire N__45797;
    wire N__45794;
    wire N__45791;
    wire N__45788;
    wire N__45785;
    wire N__45782;
    wire N__45779;
    wire N__45778;
    wire N__45775;
    wire N__45772;
    wire N__45769;
    wire N__45766;
    wire N__45763;
    wire N__45758;
    wire N__45755;
    wire N__45752;
    wire N__45749;
    wire N__45746;
    wire N__45745;
    wire N__45742;
    wire N__45739;
    wire N__45736;
    wire N__45733;
    wire N__45728;
    wire N__45725;
    wire N__45722;
    wire N__45721;
    wire N__45718;
    wire N__45717;
    wire N__45714;
    wire N__45713;
    wire N__45710;
    wire N__45707;
    wire N__45704;
    wire N__45701;
    wire N__45696;
    wire N__45691;
    wire N__45688;
    wire N__45685;
    wire N__45680;
    wire N__45677;
    wire N__45674;
    wire N__45671;
    wire N__45668;
    wire N__45665;
    wire N__45662;
    wire N__45659;
    wire N__45658;
    wire N__45657;
    wire N__45656;
    wire N__45655;
    wire N__45654;
    wire N__45653;
    wire N__45650;
    wire N__45647;
    wire N__45640;
    wire N__45635;
    wire N__45632;
    wire N__45629;
    wire N__45626;
    wire N__45625;
    wire N__45622;
    wire N__45619;
    wire N__45614;
    wire N__45611;
    wire N__45606;
    wire N__45599;
    wire N__45598;
    wire N__45597;
    wire N__45596;
    wire N__45591;
    wire N__45590;
    wire N__45587;
    wire N__45584;
    wire N__45581;
    wire N__45578;
    wire N__45575;
    wire N__45572;
    wire N__45565;
    wire N__45562;
    wire N__45557;
    wire N__45554;
    wire N__45551;
    wire N__45548;
    wire N__45545;
    wire N__45542;
    wire N__45539;
    wire N__45536;
    wire N__45533;
    wire N__45530;
    wire N__45527;
    wire N__45524;
    wire N__45521;
    wire N__45518;
    wire N__45515;
    wire N__45512;
    wire N__45511;
    wire N__45506;
    wire N__45505;
    wire N__45504;
    wire N__45503;
    wire N__45502;
    wire N__45501;
    wire N__45498;
    wire N__45497;
    wire N__45496;
    wire N__45495;
    wire N__45494;
    wire N__45493;
    wire N__45490;
    wire N__45489;
    wire N__45488;
    wire N__45487;
    wire N__45486;
    wire N__45485;
    wire N__45484;
    wire N__45483;
    wire N__45482;
    wire N__45481;
    wire N__45478;
    wire N__45475;
    wire N__45474;
    wire N__45469;
    wire N__45466;
    wire N__45461;
    wire N__45460;
    wire N__45457;
    wire N__45456;
    wire N__45455;
    wire N__45454;
    wire N__45453;
    wire N__45452;
    wire N__45451;
    wire N__45448;
    wire N__45447;
    wire N__45446;
    wire N__45445;
    wire N__45434;
    wire N__45433;
    wire N__45432;
    wire N__45431;
    wire N__45430;
    wire N__45429;
    wire N__45426;
    wire N__45423;
    wire N__45420;
    wire N__45419;
    wire N__45418;
    wire N__45417;
    wire N__45416;
    wire N__45415;
    wire N__45412;
    wire N__45411;
    wire N__45410;
    wire N__45409;
    wire N__45406;
    wire N__45403;
    wire N__45396;
    wire N__45389;
    wire N__45386;
    wire N__45385;
    wire N__45382;
    wire N__45375;
    wire N__45360;
    wire N__45357;
    wire N__45354;
    wire N__45353;
    wire N__45352;
    wire N__45351;
    wire N__45350;
    wire N__45349;
    wire N__45348;
    wire N__45347;
    wire N__45346;
    wire N__45345;
    wire N__45344;
    wire N__45343;
    wire N__45342;
    wire N__45341;
    wire N__45340;
    wire N__45331;
    wire N__45330;
    wire N__45329;
    wire N__45324;
    wire N__45317;
    wire N__45302;
    wire N__45299;
    wire N__45296;
    wire N__45295;
    wire N__45294;
    wire N__45293;
    wire N__45292;
    wire N__45291;
    wire N__45284;
    wire N__45281;
    wire N__45280;
    wire N__45277;
    wire N__45270;
    wire N__45267;
    wire N__45264;
    wire N__45255;
    wire N__45254;
    wire N__45253;
    wire N__45252;
    wire N__45251;
    wire N__45250;
    wire N__45249;
    wire N__45248;
    wire N__45247;
    wire N__45246;
    wire N__45245;
    wire N__45242;
    wire N__45239;
    wire N__45238;
    wire N__45235;
    wire N__45234;
    wire N__45233;
    wire N__45232;
    wire N__45231;
    wire N__45228;
    wire N__45227;
    wire N__45226;
    wire N__45223;
    wire N__45220;
    wire N__45217;
    wire N__45214;
    wire N__45213;
    wire N__45212;
    wire N__45211;
    wire N__45210;
    wire N__45209;
    wire N__45208;
    wire N__45207;
    wire N__45206;
    wire N__45205;
    wire N__45204;
    wire N__45203;
    wire N__45202;
    wire N__45201;
    wire N__45200;
    wire N__45199;
    wire N__45198;
    wire N__45197;
    wire N__45196;
    wire N__45193;
    wire N__45190;
    wire N__45185;
    wire N__45178;
    wire N__45173;
    wire N__45168;
    wire N__45165;
    wire N__45164;
    wire N__45163;
    wire N__45162;
    wire N__45161;
    wire N__45160;
    wire N__45159;
    wire N__45158;
    wire N__45157;
    wire N__45156;
    wire N__45155;
    wire N__45154;
    wire N__45153;
    wire N__45152;
    wire N__45149;
    wire N__45146;
    wire N__45143;
    wire N__45142;
    wire N__45141;
    wire N__45140;
    wire N__45137;
    wire N__45134;
    wire N__45123;
    wire N__45118;
    wire N__45117;
    wire N__45116;
    wire N__45115;
    wire N__45114;
    wire N__45113;
    wire N__45112;
    wire N__45111;
    wire N__45110;
    wire N__45107;
    wire N__45106;
    wire N__45105;
    wire N__45100;
    wire N__45093;
    wire N__45088;
    wire N__45081;
    wire N__45078;
    wire N__45077;
    wire N__45072;
    wire N__45069;
    wire N__45068;
    wire N__45067;
    wire N__45066;
    wire N__45057;
    wire N__45056;
    wire N__45055;
    wire N__45054;
    wire N__45053;
    wire N__45052;
    wire N__45051;
    wire N__45050;
    wire N__45047;
    wire N__45032;
    wire N__45029;
    wire N__45020;
    wire N__45017;
    wire N__45014;
    wire N__45007;
    wire N__45000;
    wire N__44997;
    wire N__44984;
    wire N__44981;
    wire N__44978;
    wire N__44969;
    wire N__44968;
    wire N__44963;
    wire N__44960;
    wire N__44953;
    wire N__44952;
    wire N__44951;
    wire N__44950;
    wire N__44949;
    wire N__44948;
    wire N__44947;
    wire N__44946;
    wire N__44945;
    wire N__44944;
    wire N__44941;
    wire N__44938;
    wire N__44937;
    wire N__44936;
    wire N__44935;
    wire N__44934;
    wire N__44929;
    wire N__44926;
    wire N__44923;
    wire N__44918;
    wire N__44913;
    wire N__44908;
    wire N__44903;
    wire N__44902;
    wire N__44899;
    wire N__44894;
    wire N__44891;
    wire N__44890;
    wire N__44889;
    wire N__44888;
    wire N__44885;
    wire N__44876;
    wire N__44867;
    wire N__44866;
    wire N__44865;
    wire N__44862;
    wire N__44859;
    wire N__44854;
    wire N__44847;
    wire N__44844;
    wire N__44839;
    wire N__44836;
    wire N__44827;
    wire N__44824;
    wire N__44817;
    wire N__44812;
    wire N__44801;
    wire N__44796;
    wire N__44793;
    wire N__44792;
    wire N__44791;
    wire N__44786;
    wire N__44783;
    wire N__44776;
    wire N__44769;
    wire N__44768;
    wire N__44767;
    wire N__44762;
    wire N__44759;
    wire N__44746;
    wire N__44741;
    wire N__44730;
    wire N__44727;
    wire N__44722;
    wire N__44713;
    wire N__44710;
    wire N__44705;
    wire N__44700;
    wire N__44689;
    wire N__44672;
    wire N__44665;
    wire N__44656;
    wire N__44653;
    wire N__44652;
    wire N__44651;
    wire N__44650;
    wire N__44649;
    wire N__44648;
    wire N__44645;
    wire N__44640;
    wire N__44637;
    wire N__44632;
    wire N__44625;
    wire N__44614;
    wire N__44609;
    wire N__44606;
    wire N__44601;
    wire N__44594;
    wire N__44589;
    wire N__44584;
    wire N__44579;
    wire N__44576;
    wire N__44561;
    wire N__44558;
    wire N__44555;
    wire N__44552;
    wire N__44551;
    wire N__44548;
    wire N__44545;
    wire N__44540;
    wire N__44537;
    wire N__44534;
    wire N__44533;
    wire N__44530;
    wire N__44527;
    wire N__44522;
    wire N__44519;
    wire N__44516;
    wire N__44513;
    wire N__44512;
    wire N__44509;
    wire N__44506;
    wire N__44503;
    wire N__44500;
    wire N__44495;
    wire N__44492;
    wire N__44489;
    wire N__44488;
    wire N__44485;
    wire N__44482;
    wire N__44481;
    wire N__44478;
    wire N__44475;
    wire N__44474;
    wire N__44471;
    wire N__44468;
    wire N__44465;
    wire N__44462;
    wire N__44453;
    wire N__44450;
    wire N__44447;
    wire N__44444;
    wire N__44441;
    wire N__44438;
    wire N__44435;
    wire N__44432;
    wire N__44429;
    wire N__44426;
    wire N__44423;
    wire N__44420;
    wire N__44419;
    wire N__44416;
    wire N__44413;
    wire N__44410;
    wire N__44407;
    wire N__44402;
    wire N__44399;
    wire N__44396;
    wire N__44395;
    wire N__44392;
    wire N__44389;
    wire N__44388;
    wire N__44383;
    wire N__44380;
    wire N__44375;
    wire N__44372;
    wire N__44369;
    wire N__44368;
    wire N__44365;
    wire N__44362;
    wire N__44359;
    wire N__44354;
    wire N__44351;
    wire N__44348;
    wire N__44345;
    wire N__44342;
    wire N__44339;
    wire N__44336;
    wire N__44333;
    wire N__44330;
    wire N__44327;
    wire N__44324;
    wire N__44321;
    wire N__44318;
    wire N__44315;
    wire N__44312;
    wire N__44309;
    wire N__44306;
    wire N__44303;
    wire N__44300;
    wire N__44297;
    wire N__44294;
    wire N__44291;
    wire N__44288;
    wire N__44285;
    wire N__44282;
    wire N__44279;
    wire N__44276;
    wire N__44273;
    wire N__44272;
    wire N__44269;
    wire N__44268;
    wire N__44265;
    wire N__44264;
    wire N__44261;
    wire N__44258;
    wire N__44255;
    wire N__44252;
    wire N__44247;
    wire N__44240;
    wire N__44237;
    wire N__44234;
    wire N__44231;
    wire N__44228;
    wire N__44225;
    wire N__44222;
    wire N__44219;
    wire N__44216;
    wire N__44213;
    wire N__44210;
    wire N__44209;
    wire N__44206;
    wire N__44203;
    wire N__44200;
    wire N__44197;
    wire N__44192;
    wire N__44189;
    wire N__44188;
    wire N__44187;
    wire N__44186;
    wire N__44183;
    wire N__44180;
    wire N__44177;
    wire N__44174;
    wire N__44173;
    wire N__44168;
    wire N__44165;
    wire N__44162;
    wire N__44159;
    wire N__44156;
    wire N__44153;
    wire N__44148;
    wire N__44141;
    wire N__44140;
    wire N__44139;
    wire N__44138;
    wire N__44135;
    wire N__44132;
    wire N__44129;
    wire N__44128;
    wire N__44125;
    wire N__44124;
    wire N__44123;
    wire N__44120;
    wire N__44115;
    wire N__44112;
    wire N__44109;
    wire N__44106;
    wire N__44103;
    wire N__44100;
    wire N__44095;
    wire N__44084;
    wire N__44081;
    wire N__44080;
    wire N__44077;
    wire N__44074;
    wire N__44069;
    wire N__44066;
    wire N__44063;
    wire N__44060;
    wire N__44057;
    wire N__44054;
    wire N__44051;
    wire N__44050;
    wire N__44047;
    wire N__44046;
    wire N__44043;
    wire N__44040;
    wire N__44037;
    wire N__44034;
    wire N__44029;
    wire N__44026;
    wire N__44023;
    wire N__44020;
    wire N__44015;
    wire N__44014;
    wire N__44013;
    wire N__44010;
    wire N__44005;
    wire N__44002;
    wire N__44001;
    wire N__44000;
    wire N__43995;
    wire N__43994;
    wire N__43991;
    wire N__43988;
    wire N__43985;
    wire N__43980;
    wire N__43973;
    wire N__43970;
    wire N__43967;
    wire N__43964;
    wire N__43961;
    wire N__43958;
    wire N__43955;
    wire N__43952;
    wire N__43949;
    wire N__43948;
    wire N__43947;
    wire N__43946;
    wire N__43945;
    wire N__43944;
    wire N__43941;
    wire N__43940;
    wire N__43937;
    wire N__43934;
    wire N__43931;
    wire N__43926;
    wire N__43923;
    wire N__43920;
    wire N__43917;
    wire N__43914;
    wire N__43911;
    wire N__43906;
    wire N__43901;
    wire N__43898;
    wire N__43889;
    wire N__43886;
    wire N__43883;
    wire N__43880;
    wire N__43879;
    wire N__43876;
    wire N__43873;
    wire N__43868;
    wire N__43865;
    wire N__43862;
    wire N__43859;
    wire N__43858;
    wire N__43855;
    wire N__43852;
    wire N__43849;
    wire N__43846;
    wire N__43841;
    wire N__43838;
    wire N__43835;
    wire N__43832;
    wire N__43829;
    wire N__43826;
    wire N__43825;
    wire N__43820;
    wire N__43817;
    wire N__43814;
    wire N__43811;
    wire N__43810;
    wire N__43807;
    wire N__43804;
    wire N__43803;
    wire N__43798;
    wire N__43797;
    wire N__43796;
    wire N__43793;
    wire N__43790;
    wire N__43787;
    wire N__43784;
    wire N__43777;
    wire N__43772;
    wire N__43771;
    wire N__43770;
    wire N__43769;
    wire N__43766;
    wire N__43763;
    wire N__43760;
    wire N__43757;
    wire N__43754;
    wire N__43751;
    wire N__43750;
    wire N__43749;
    wire N__43746;
    wire N__43743;
    wire N__43738;
    wire N__43733;
    wire N__43726;
    wire N__43721;
    wire N__43718;
    wire N__43715;
    wire N__43712;
    wire N__43709;
    wire N__43708;
    wire N__43705;
    wire N__43702;
    wire N__43699;
    wire N__43696;
    wire N__43693;
    wire N__43690;
    wire N__43687;
    wire N__43682;
    wire N__43679;
    wire N__43676;
    wire N__43673;
    wire N__43672;
    wire N__43669;
    wire N__43666;
    wire N__43661;
    wire N__43658;
    wire N__43655;
    wire N__43652;
    wire N__43651;
    wire N__43650;
    wire N__43649;
    wire N__43648;
    wire N__43647;
    wire N__43646;
    wire N__43643;
    wire N__43640;
    wire N__43637;
    wire N__43634;
    wire N__43631;
    wire N__43628;
    wire N__43625;
    wire N__43620;
    wire N__43617;
    wire N__43614;
    wire N__43607;
    wire N__43604;
    wire N__43601;
    wire N__43592;
    wire N__43589;
    wire N__43588;
    wire N__43585;
    wire N__43584;
    wire N__43581;
    wire N__43580;
    wire N__43577;
    wire N__43574;
    wire N__43571;
    wire N__43568;
    wire N__43563;
    wire N__43562;
    wire N__43561;
    wire N__43558;
    wire N__43555;
    wire N__43552;
    wire N__43549;
    wire N__43546;
    wire N__43543;
    wire N__43532;
    wire N__43529;
    wire N__43528;
    wire N__43527;
    wire N__43524;
    wire N__43521;
    wire N__43518;
    wire N__43515;
    wire N__43512;
    wire N__43509;
    wire N__43502;
    wire N__43499;
    wire N__43496;
    wire N__43493;
    wire N__43490;
    wire N__43487;
    wire N__43486;
    wire N__43483;
    wire N__43480;
    wire N__43475;
    wire N__43472;
    wire N__43469;
    wire N__43466;
    wire N__43465;
    wire N__43462;
    wire N__43461;
    wire N__43458;
    wire N__43455;
    wire N__43452;
    wire N__43449;
    wire N__43446;
    wire N__43439;
    wire N__43436;
    wire N__43433;
    wire N__43430;
    wire N__43427;
    wire N__43424;
    wire N__43421;
    wire N__43420;
    wire N__43417;
    wire N__43414;
    wire N__43413;
    wire N__43410;
    wire N__43409;
    wire N__43408;
    wire N__43407;
    wire N__43404;
    wire N__43401;
    wire N__43398;
    wire N__43395;
    wire N__43394;
    wire N__43391;
    wire N__43388;
    wire N__43385;
    wire N__43380;
    wire N__43375;
    wire N__43370;
    wire N__43361;
    wire N__43358;
    wire N__43355;
    wire N__43352;
    wire N__43351;
    wire N__43348;
    wire N__43345;
    wire N__43342;
    wire N__43339;
    wire N__43334;
    wire N__43333;
    wire N__43332;
    wire N__43329;
    wire N__43328;
    wire N__43325;
    wire N__43322;
    wire N__43319;
    wire N__43316;
    wire N__43313;
    wire N__43308;
    wire N__43301;
    wire N__43300;
    wire N__43297;
    wire N__43294;
    wire N__43291;
    wire N__43288;
    wire N__43285;
    wire N__43280;
    wire N__43277;
    wire N__43274;
    wire N__43271;
    wire N__43270;
    wire N__43269;
    wire N__43266;
    wire N__43263;
    wire N__43260;
    wire N__43257;
    wire N__43254;
    wire N__43251;
    wire N__43248;
    wire N__43245;
    wire N__43242;
    wire N__43235;
    wire N__43232;
    wire N__43231;
    wire N__43230;
    wire N__43227;
    wire N__43226;
    wire N__43223;
    wire N__43220;
    wire N__43217;
    wire N__43214;
    wire N__43211;
    wire N__43202;
    wire N__43199;
    wire N__43196;
    wire N__43193;
    wire N__43190;
    wire N__43187;
    wire N__43184;
    wire N__43181;
    wire N__43180;
    wire N__43177;
    wire N__43174;
    wire N__43171;
    wire N__43166;
    wire N__43163;
    wire N__43160;
    wire N__43157;
    wire N__43154;
    wire N__43151;
    wire N__43148;
    wire N__43145;
    wire N__43142;
    wire N__43139;
    wire N__43136;
    wire N__43133;
    wire N__43132;
    wire N__43129;
    wire N__43126;
    wire N__43121;
    wire N__43118;
    wire N__43115;
    wire N__43112;
    wire N__43109;
    wire N__43106;
    wire N__43103;
    wire N__43100;
    wire N__43097;
    wire N__43094;
    wire N__43091;
    wire N__43088;
    wire N__43085;
    wire N__43082;
    wire N__43079;
    wire N__43076;
    wire N__43073;
    wire N__43070;
    wire N__43069;
    wire N__43068;
    wire N__43065;
    wire N__43062;
    wire N__43059;
    wire N__43052;
    wire N__43051;
    wire N__43050;
    wire N__43047;
    wire N__43044;
    wire N__43041;
    wire N__43034;
    wire N__43031;
    wire N__43028;
    wire N__43027;
    wire N__43026;
    wire N__43023;
    wire N__43020;
    wire N__43017;
    wire N__43010;
    wire N__43007;
    wire N__43006;
    wire N__43003;
    wire N__43002;
    wire N__42999;
    wire N__42996;
    wire N__42993;
    wire N__42986;
    wire N__42985;
    wire N__42984;
    wire N__42983;
    wire N__42980;
    wire N__42979;
    wire N__42976;
    wire N__42971;
    wire N__42968;
    wire N__42965;
    wire N__42962;
    wire N__42959;
    wire N__42956;
    wire N__42951;
    wire N__42950;
    wire N__42947;
    wire N__42942;
    wire N__42939;
    wire N__42932;
    wire N__42931;
    wire N__42930;
    wire N__42927;
    wire N__42924;
    wire N__42921;
    wire N__42916;
    wire N__42915;
    wire N__42914;
    wire N__42913;
    wire N__42910;
    wire N__42907;
    wire N__42900;
    wire N__42893;
    wire N__42892;
    wire N__42889;
    wire N__42888;
    wire N__42885;
    wire N__42884;
    wire N__42881;
    wire N__42878;
    wire N__42875;
    wire N__42874;
    wire N__42871;
    wire N__42870;
    wire N__42867;
    wire N__42862;
    wire N__42859;
    wire N__42856;
    wire N__42853;
    wire N__42848;
    wire N__42839;
    wire N__42838;
    wire N__42837;
    wire N__42836;
    wire N__42833;
    wire N__42830;
    wire N__42829;
    wire N__42828;
    wire N__42827;
    wire N__42824;
    wire N__42821;
    wire N__42818;
    wire N__42815;
    wire N__42808;
    wire N__42797;
    wire N__42794;
    wire N__42793;
    wire N__42790;
    wire N__42787;
    wire N__42784;
    wire N__42779;
    wire N__42778;
    wire N__42775;
    wire N__42772;
    wire N__42769;
    wire N__42764;
    wire N__42761;
    wire N__42758;
    wire N__42755;
    wire N__42752;
    wire N__42749;
    wire N__42746;
    wire N__42745;
    wire N__42744;
    wire N__42741;
    wire N__42736;
    wire N__42731;
    wire N__42730;
    wire N__42729;
    wire N__42726;
    wire N__42723;
    wire N__42720;
    wire N__42713;
    wire N__42712;
    wire N__42709;
    wire N__42708;
    wire N__42707;
    wire N__42706;
    wire N__42701;
    wire N__42698;
    wire N__42697;
    wire N__42696;
    wire N__42693;
    wire N__42692;
    wire N__42689;
    wire N__42686;
    wire N__42683;
    wire N__42678;
    wire N__42675;
    wire N__42672;
    wire N__42669;
    wire N__42660;
    wire N__42657;
    wire N__42656;
    wire N__42653;
    wire N__42650;
    wire N__42647;
    wire N__42644;
    wire N__42635;
    wire N__42632;
    wire N__42629;
    wire N__42628;
    wire N__42625;
    wire N__42622;
    wire N__42617;
    wire N__42616;
    wire N__42613;
    wire N__42610;
    wire N__42607;
    wire N__42602;
    wire N__42601;
    wire N__42598;
    wire N__42595;
    wire N__42590;
    wire N__42587;
    wire N__42584;
    wire N__42581;
    wire N__42580;
    wire N__42579;
    wire N__42576;
    wire N__42575;
    wire N__42574;
    wire N__42573;
    wire N__42572;
    wire N__42571;
    wire N__42570;
    wire N__42569;
    wire N__42568;
    wire N__42567;
    wire N__42566;
    wire N__42563;
    wire N__42562;
    wire N__42561;
    wire N__42556;
    wire N__42555;
    wire N__42554;
    wire N__42553;
    wire N__42552;
    wire N__42551;
    wire N__42546;
    wire N__42541;
    wire N__42538;
    wire N__42535;
    wire N__42532;
    wire N__42529;
    wire N__42526;
    wire N__42521;
    wire N__42516;
    wire N__42513;
    wire N__42510;
    wire N__42507;
    wire N__42504;
    wire N__42499;
    wire N__42496;
    wire N__42493;
    wire N__42488;
    wire N__42461;
    wire N__42458;
    wire N__42455;
    wire N__42452;
    wire N__42449;
    wire N__42448;
    wire N__42445;
    wire N__42442;
    wire N__42439;
    wire N__42438;
    wire N__42437;
    wire N__42436;
    wire N__42435;
    wire N__42434;
    wire N__42433;
    wire N__42432;
    wire N__42431;
    wire N__42430;
    wire N__42429;
    wire N__42428;
    wire N__42427;
    wire N__42424;
    wire N__42421;
    wire N__42416;
    wire N__42407;
    wire N__42400;
    wire N__42393;
    wire N__42380;
    wire N__42379;
    wire N__42376;
    wire N__42375;
    wire N__42374;
    wire N__42371;
    wire N__42368;
    wire N__42363;
    wire N__42356;
    wire N__42355;
    wire N__42354;
    wire N__42353;
    wire N__42350;
    wire N__42347;
    wire N__42342;
    wire N__42335;
    wire N__42334;
    wire N__42333;
    wire N__42330;
    wire N__42329;
    wire N__42326;
    wire N__42323;
    wire N__42320;
    wire N__42315;
    wire N__42312;
    wire N__42309;
    wire N__42302;
    wire N__42301;
    wire N__42300;
    wire N__42297;
    wire N__42296;
    wire N__42293;
    wire N__42290;
    wire N__42287;
    wire N__42284;
    wire N__42275;
    wire N__42272;
    wire N__42269;
    wire N__42266;
    wire N__42263;
    wire N__42260;
    wire N__42257;
    wire N__42254;
    wire N__42251;
    wire N__42248;
    wire N__42245;
    wire N__42242;
    wire N__42241;
    wire N__42240;
    wire N__42237;
    wire N__42234;
    wire N__42231;
    wire N__42224;
    wire N__42221;
    wire N__42218;
    wire N__42215;
    wire N__42212;
    wire N__42209;
    wire N__42206;
    wire N__42205;
    wire N__42202;
    wire N__42199;
    wire N__42196;
    wire N__42191;
    wire N__42188;
    wire N__42185;
    wire N__42184;
    wire N__42183;
    wire N__42180;
    wire N__42177;
    wire N__42176;
    wire N__42175;
    wire N__42172;
    wire N__42167;
    wire N__42162;
    wire N__42155;
    wire N__42154;
    wire N__42151;
    wire N__42148;
    wire N__42143;
    wire N__42142;
    wire N__42139;
    wire N__42136;
    wire N__42131;
    wire N__42128;
    wire N__42127;
    wire N__42126;
    wire N__42123;
    wire N__42120;
    wire N__42117;
    wire N__42110;
    wire N__42109;
    wire N__42108;
    wire N__42103;
    wire N__42100;
    wire N__42095;
    wire N__42092;
    wire N__42089;
    wire N__42086;
    wire N__42083;
    wire N__42082;
    wire N__42081;
    wire N__42078;
    wire N__42075;
    wire N__42072;
    wire N__42069;
    wire N__42066;
    wire N__42065;
    wire N__42058;
    wire N__42055;
    wire N__42050;
    wire N__42049;
    wire N__42048;
    wire N__42047;
    wire N__42044;
    wire N__42041;
    wire N__42038;
    wire N__42035;
    wire N__42032;
    wire N__42029;
    wire N__42026;
    wire N__42023;
    wire N__42014;
    wire N__42011;
    wire N__42008;
    wire N__42005;
    wire N__42004;
    wire N__42003;
    wire N__42000;
    wire N__41995;
    wire N__41990;
    wire N__41989;
    wire N__41988;
    wire N__41985;
    wire N__41980;
    wire N__41975;
    wire N__41974;
    wire N__41971;
    wire N__41968;
    wire N__41965;
    wire N__41964;
    wire N__41961;
    wire N__41960;
    wire N__41957;
    wire N__41954;
    wire N__41951;
    wire N__41948;
    wire N__41945;
    wire N__41936;
    wire N__41935;
    wire N__41932;
    wire N__41931;
    wire N__41928;
    wire N__41927;
    wire N__41924;
    wire N__41921;
    wire N__41918;
    wire N__41915;
    wire N__41910;
    wire N__41907;
    wire N__41900;
    wire N__41897;
    wire N__41894;
    wire N__41891;
    wire N__41888;
    wire N__41885;
    wire N__41882;
    wire N__41881;
    wire N__41878;
    wire N__41875;
    wire N__41872;
    wire N__41869;
    wire N__41864;
    wire N__41861;
    wire N__41858;
    wire N__41855;
    wire N__41852;
    wire N__41849;
    wire N__41846;
    wire N__41845;
    wire N__41842;
    wire N__41839;
    wire N__41836;
    wire N__41833;
    wire N__41828;
    wire N__41825;
    wire N__41822;
    wire N__41821;
    wire N__41818;
    wire N__41815;
    wire N__41810;
    wire N__41807;
    wire N__41804;
    wire N__41801;
    wire N__41798;
    wire N__41797;
    wire N__41794;
    wire N__41793;
    wire N__41792;
    wire N__41789;
    wire N__41786;
    wire N__41783;
    wire N__41780;
    wire N__41775;
    wire N__41772;
    wire N__41769;
    wire N__41766;
    wire N__41759;
    wire N__41756;
    wire N__41755;
    wire N__41752;
    wire N__41749;
    wire N__41744;
    wire N__41743;
    wire N__41740;
    wire N__41739;
    wire N__41738;
    wire N__41735;
    wire N__41732;
    wire N__41727;
    wire N__41722;
    wire N__41717;
    wire N__41716;
    wire N__41713;
    wire N__41710;
    wire N__41707;
    wire N__41704;
    wire N__41699;
    wire N__41696;
    wire N__41693;
    wire N__41690;
    wire N__41689;
    wire N__41686;
    wire N__41683;
    wire N__41678;
    wire N__41675;
    wire N__41672;
    wire N__41669;
    wire N__41668;
    wire N__41665;
    wire N__41662;
    wire N__41657;
    wire N__41656;
    wire N__41653;
    wire N__41650;
    wire N__41649;
    wire N__41648;
    wire N__41645;
    wire N__41642;
    wire N__41637;
    wire N__41634;
    wire N__41631;
    wire N__41624;
    wire N__41623;
    wire N__41622;
    wire N__41621;
    wire N__41616;
    wire N__41615;
    wire N__41614;
    wire N__41611;
    wire N__41608;
    wire N__41605;
    wire N__41600;
    wire N__41591;
    wire N__41588;
    wire N__41587;
    wire N__41584;
    wire N__41581;
    wire N__41578;
    wire N__41575;
    wire N__41570;
    wire N__41567;
    wire N__41564;
    wire N__41561;
    wire N__41558;
    wire N__41555;
    wire N__41552;
    wire N__41549;
    wire N__41546;
    wire N__41545;
    wire N__41542;
    wire N__41541;
    wire N__41538;
    wire N__41535;
    wire N__41532;
    wire N__41525;
    wire N__41522;
    wire N__41519;
    wire N__41516;
    wire N__41513;
    wire N__41510;
    wire N__41507;
    wire N__41504;
    wire N__41501;
    wire N__41500;
    wire N__41497;
    wire N__41494;
    wire N__41491;
    wire N__41488;
    wire N__41483;
    wire N__41480;
    wire N__41477;
    wire N__41476;
    wire N__41473;
    wire N__41470;
    wire N__41467;
    wire N__41464;
    wire N__41461;
    wire N__41458;
    wire N__41453;
    wire N__41450;
    wire N__41447;
    wire N__41444;
    wire N__41441;
    wire N__41438;
    wire N__41435;
    wire N__41432;
    wire N__41429;
    wire N__41426;
    wire N__41423;
    wire N__41420;
    wire N__41417;
    wire N__41414;
    wire N__41411;
    wire N__41410;
    wire N__41407;
    wire N__41404;
    wire N__41401;
    wire N__41398;
    wire N__41393;
    wire N__41390;
    wire N__41387;
    wire N__41384;
    wire N__41381;
    wire N__41378;
    wire N__41375;
    wire N__41372;
    wire N__41369;
    wire N__41366;
    wire N__41363;
    wire N__41360;
    wire N__41357;
    wire N__41354;
    wire N__41351;
    wire N__41348;
    wire N__41345;
    wire N__41342;
    wire N__41339;
    wire N__41336;
    wire N__41333;
    wire N__41330;
    wire N__41327;
    wire N__41324;
    wire N__41321;
    wire N__41320;
    wire N__41317;
    wire N__41314;
    wire N__41311;
    wire N__41306;
    wire N__41303;
    wire N__41300;
    wire N__41299;
    wire N__41296;
    wire N__41293;
    wire N__41288;
    wire N__41285;
    wire N__41282;
    wire N__41281;
    wire N__41278;
    wire N__41275;
    wire N__41270;
    wire N__41267;
    wire N__41266;
    wire N__41263;
    wire N__41260;
    wire N__41255;
    wire N__41254;
    wire N__41251;
    wire N__41248;
    wire N__41245;
    wire N__41244;
    wire N__41241;
    wire N__41238;
    wire N__41237;
    wire N__41234;
    wire N__41231;
    wire N__41228;
    wire N__41225;
    wire N__41216;
    wire N__41213;
    wire N__41210;
    wire N__41209;
    wire N__41206;
    wire N__41203;
    wire N__41200;
    wire N__41195;
    wire N__41192;
    wire N__41189;
    wire N__41186;
    wire N__41183;
    wire N__41180;
    wire N__41177;
    wire N__41174;
    wire N__41171;
    wire N__41168;
    wire N__41165;
    wire N__41162;
    wire N__41159;
    wire N__41156;
    wire N__41153;
    wire N__41150;
    wire N__41147;
    wire N__41144;
    wire N__41141;
    wire N__41138;
    wire N__41135;
    wire N__41132;
    wire N__41129;
    wire N__41126;
    wire N__41123;
    wire N__41122;
    wire N__41121;
    wire N__41118;
    wire N__41115;
    wire N__41112;
    wire N__41107;
    wire N__41102;
    wire N__41101;
    wire N__41100;
    wire N__41097;
    wire N__41092;
    wire N__41087;
    wire N__41086;
    wire N__41085;
    wire N__41082;
    wire N__41079;
    wire N__41076;
    wire N__41073;
    wire N__41066;
    wire N__41065;
    wire N__41064;
    wire N__41061;
    wire N__41058;
    wire N__41055;
    wire N__41048;
    wire N__41047;
    wire N__41044;
    wire N__41043;
    wire N__41040;
    wire N__41037;
    wire N__41036;
    wire N__41033;
    wire N__41028;
    wire N__41025;
    wire N__41018;
    wire N__41015;
    wire N__41012;
    wire N__41011;
    wire N__41010;
    wire N__41009;
    wire N__41006;
    wire N__41003;
    wire N__41000;
    wire N__40997;
    wire N__40994;
    wire N__40989;
    wire N__40982;
    wire N__40981;
    wire N__40978;
    wire N__40975;
    wire N__40974;
    wire N__40969;
    wire N__40968;
    wire N__40965;
    wire N__40962;
    wire N__40959;
    wire N__40952;
    wire N__40949;
    wire N__40946;
    wire N__40943;
    wire N__40942;
    wire N__40939;
    wire N__40936;
    wire N__40931;
    wire N__40928;
    wire N__40925;
    wire N__40922;
    wire N__40919;
    wire N__40916;
    wire N__40913;
    wire N__40910;
    wire N__40907;
    wire N__40904;
    wire N__40901;
    wire N__40898;
    wire N__40895;
    wire N__40892;
    wire N__40889;
    wire N__40886;
    wire N__40883;
    wire N__40880;
    wire N__40877;
    wire N__40874;
    wire N__40871;
    wire N__40868;
    wire N__40865;
    wire N__40862;
    wire N__40859;
    wire N__40856;
    wire N__40853;
    wire N__40850;
    wire N__40849;
    wire N__40848;
    wire N__40847;
    wire N__40846;
    wire N__40843;
    wire N__40838;
    wire N__40835;
    wire N__40832;
    wire N__40831;
    wire N__40824;
    wire N__40819;
    wire N__40814;
    wire N__40811;
    wire N__40808;
    wire N__40807;
    wire N__40804;
    wire N__40801;
    wire N__40796;
    wire N__40793;
    wire N__40792;
    wire N__40789;
    wire N__40786;
    wire N__40783;
    wire N__40780;
    wire N__40777;
    wire N__40772;
    wire N__40769;
    wire N__40766;
    wire N__40765;
    wire N__40762;
    wire N__40759;
    wire N__40756;
    wire N__40753;
    wire N__40748;
    wire N__40745;
    wire N__40744;
    wire N__40743;
    wire N__40742;
    wire N__40741;
    wire N__40740;
    wire N__40733;
    wire N__40730;
    wire N__40729;
    wire N__40728;
    wire N__40725;
    wire N__40722;
    wire N__40717;
    wire N__40712;
    wire N__40703;
    wire N__40702;
    wire N__40701;
    wire N__40698;
    wire N__40697;
    wire N__40694;
    wire N__40693;
    wire N__40690;
    wire N__40687;
    wire N__40686;
    wire N__40683;
    wire N__40680;
    wire N__40677;
    wire N__40674;
    wire N__40671;
    wire N__40666;
    wire N__40655;
    wire N__40652;
    wire N__40649;
    wire N__40646;
    wire N__40643;
    wire N__40640;
    wire N__40637;
    wire N__40634;
    wire N__40631;
    wire N__40628;
    wire N__40625;
    wire N__40622;
    wire N__40619;
    wire N__40616;
    wire N__40615;
    wire N__40612;
    wire N__40609;
    wire N__40606;
    wire N__40603;
    wire N__40598;
    wire N__40595;
    wire N__40592;
    wire N__40589;
    wire N__40588;
    wire N__40585;
    wire N__40582;
    wire N__40579;
    wire N__40576;
    wire N__40571;
    wire N__40568;
    wire N__40565;
    wire N__40562;
    wire N__40561;
    wire N__40558;
    wire N__40555;
    wire N__40550;
    wire N__40547;
    wire N__40544;
    wire N__40541;
    wire N__40538;
    wire N__40535;
    wire N__40532;
    wire N__40529;
    wire N__40526;
    wire N__40523;
    wire N__40520;
    wire N__40517;
    wire N__40514;
    wire N__40511;
    wire N__40508;
    wire N__40505;
    wire N__40502;
    wire N__40501;
    wire N__40498;
    wire N__40497;
    wire N__40496;
    wire N__40493;
    wire N__40490;
    wire N__40485;
    wire N__40482;
    wire N__40477;
    wire N__40472;
    wire N__40471;
    wire N__40468;
    wire N__40465;
    wire N__40460;
    wire N__40459;
    wire N__40456;
    wire N__40453;
    wire N__40452;
    wire N__40451;
    wire N__40446;
    wire N__40445;
    wire N__40444;
    wire N__40441;
    wire N__40438;
    wire N__40435;
    wire N__40430;
    wire N__40427;
    wire N__40418;
    wire N__40415;
    wire N__40414;
    wire N__40413;
    wire N__40408;
    wire N__40405;
    wire N__40404;
    wire N__40403;
    wire N__40402;
    wire N__40397;
    wire N__40394;
    wire N__40389;
    wire N__40386;
    wire N__40379;
    wire N__40376;
    wire N__40375;
    wire N__40374;
    wire N__40373;
    wire N__40372;
    wire N__40371;
    wire N__40370;
    wire N__40369;
    wire N__40366;
    wire N__40363;
    wire N__40354;
    wire N__40351;
    wire N__40350;
    wire N__40347;
    wire N__40346;
    wire N__40343;
    wire N__40340;
    wire N__40339;
    wire N__40338;
    wire N__40337;
    wire N__40334;
    wire N__40329;
    wire N__40326;
    wire N__40325;
    wire N__40324;
    wire N__40321;
    wire N__40316;
    wire N__40313;
    wire N__40308;
    wire N__40305;
    wire N__40302;
    wire N__40299;
    wire N__40294;
    wire N__40293;
    wire N__40292;
    wire N__40291;
    wire N__40290;
    wire N__40289;
    wire N__40288;
    wire N__40281;
    wire N__40278;
    wire N__40273;
    wire N__40268;
    wire N__40259;
    wire N__40254;
    wire N__40241;
    wire N__40240;
    wire N__40239;
    wire N__40238;
    wire N__40237;
    wire N__40234;
    wire N__40231;
    wire N__40226;
    wire N__40223;
    wire N__40222;
    wire N__40221;
    wire N__40216;
    wire N__40215;
    wire N__40214;
    wire N__40213;
    wire N__40210;
    wire N__40207;
    wire N__40206;
    wire N__40203;
    wire N__40200;
    wire N__40197;
    wire N__40194;
    wire N__40191;
    wire N__40188;
    wire N__40183;
    wire N__40178;
    wire N__40163;
    wire N__40162;
    wire N__40161;
    wire N__40160;
    wire N__40159;
    wire N__40156;
    wire N__40155;
    wire N__40154;
    wire N__40153;
    wire N__40150;
    wire N__40147;
    wire N__40146;
    wire N__40145;
    wire N__40142;
    wire N__40137;
    wire N__40134;
    wire N__40133;
    wire N__40130;
    wire N__40123;
    wire N__40120;
    wire N__40117;
    wire N__40112;
    wire N__40109;
    wire N__40108;
    wire N__40107;
    wire N__40104;
    wire N__40103;
    wire N__40102;
    wire N__40101;
    wire N__40096;
    wire N__40091;
    wire N__40086;
    wire N__40077;
    wire N__40072;
    wire N__40061;
    wire N__40058;
    wire N__40055;
    wire N__40054;
    wire N__40051;
    wire N__40048;
    wire N__40043;
    wire N__40040;
    wire N__40037;
    wire N__40034;
    wire N__40031;
    wire N__40028;
    wire N__40025;
    wire N__40022;
    wire N__40019;
    wire N__40016;
    wire N__40013;
    wire N__40010;
    wire N__40007;
    wire N__40004;
    wire N__40001;
    wire N__39998;
    wire N__39995;
    wire N__39992;
    wire N__39989;
    wire N__39986;
    wire N__39983;
    wire N__39980;
    wire N__39977;
    wire N__39974;
    wire N__39971;
    wire N__39968;
    wire N__39965;
    wire N__39962;
    wire N__39959;
    wire N__39956;
    wire N__39953;
    wire N__39950;
    wire N__39947;
    wire N__39944;
    wire N__39941;
    wire N__39938;
    wire N__39935;
    wire N__39932;
    wire N__39931;
    wire N__39928;
    wire N__39925;
    wire N__39922;
    wire N__39919;
    wire N__39918;
    wire N__39915;
    wire N__39912;
    wire N__39909;
    wire N__39906;
    wire N__39899;
    wire N__39896;
    wire N__39893;
    wire N__39892;
    wire N__39889;
    wire N__39886;
    wire N__39885;
    wire N__39882;
    wire N__39879;
    wire N__39878;
    wire N__39875;
    wire N__39872;
    wire N__39869;
    wire N__39866;
    wire N__39863;
    wire N__39858;
    wire N__39853;
    wire N__39850;
    wire N__39845;
    wire N__39844;
    wire N__39841;
    wire N__39838;
    wire N__39835;
    wire N__39834;
    wire N__39831;
    wire N__39828;
    wire N__39825;
    wire N__39822;
    wire N__39819;
    wire N__39812;
    wire N__39811;
    wire N__39808;
    wire N__39805;
    wire N__39800;
    wire N__39797;
    wire N__39794;
    wire N__39791;
    wire N__39788;
    wire N__39785;
    wire N__39782;
    wire N__39779;
    wire N__39778;
    wire N__39775;
    wire N__39774;
    wire N__39773;
    wire N__39772;
    wire N__39771;
    wire N__39768;
    wire N__39765;
    wire N__39758;
    wire N__39755;
    wire N__39754;
    wire N__39753;
    wire N__39752;
    wire N__39749;
    wire N__39744;
    wire N__39735;
    wire N__39732;
    wire N__39729;
    wire N__39726;
    wire N__39719;
    wire N__39718;
    wire N__39717;
    wire N__39714;
    wire N__39713;
    wire N__39712;
    wire N__39711;
    wire N__39710;
    wire N__39707;
    wire N__39704;
    wire N__39697;
    wire N__39694;
    wire N__39691;
    wire N__39690;
    wire N__39689;
    wire N__39688;
    wire N__39687;
    wire N__39684;
    wire N__39675;
    wire N__39666;
    wire N__39661;
    wire N__39656;
    wire N__39655;
    wire N__39654;
    wire N__39651;
    wire N__39650;
    wire N__39645;
    wire N__39642;
    wire N__39641;
    wire N__39638;
    wire N__39635;
    wire N__39632;
    wire N__39631;
    wire N__39626;
    wire N__39623;
    wire N__39620;
    wire N__39617;
    wire N__39608;
    wire N__39605;
    wire N__39602;
    wire N__39599;
    wire N__39596;
    wire N__39593;
    wire N__39590;
    wire N__39589;
    wire N__39588;
    wire N__39587;
    wire N__39586;
    wire N__39585;
    wire N__39584;
    wire N__39581;
    wire N__39572;
    wire N__39571;
    wire N__39566;
    wire N__39565;
    wire N__39560;
    wire N__39557;
    wire N__39556;
    wire N__39553;
    wire N__39550;
    wire N__39547;
    wire N__39544;
    wire N__39541;
    wire N__39536;
    wire N__39533;
    wire N__39528;
    wire N__39521;
    wire N__39518;
    wire N__39515;
    wire N__39512;
    wire N__39509;
    wire N__39506;
    wire N__39505;
    wire N__39502;
    wire N__39499;
    wire N__39496;
    wire N__39493;
    wire N__39488;
    wire N__39485;
    wire N__39484;
    wire N__39481;
    wire N__39478;
    wire N__39475;
    wire N__39470;
    wire N__39467;
    wire N__39464;
    wire N__39463;
    wire N__39460;
    wire N__39457;
    wire N__39454;
    wire N__39451;
    wire N__39446;
    wire N__39443;
    wire N__39440;
    wire N__39437;
    wire N__39436;
    wire N__39433;
    wire N__39430;
    wire N__39427;
    wire N__39424;
    wire N__39419;
    wire N__39416;
    wire N__39413;
    wire N__39412;
    wire N__39409;
    wire N__39406;
    wire N__39403;
    wire N__39400;
    wire N__39395;
    wire N__39392;
    wire N__39389;
    wire N__39386;
    wire N__39383;
    wire N__39380;
    wire N__39377;
    wire N__39374;
    wire N__39371;
    wire N__39368;
    wire N__39367;
    wire N__39364;
    wire N__39361;
    wire N__39358;
    wire N__39353;
    wire N__39350;
    wire N__39349;
    wire N__39346;
    wire N__39343;
    wire N__39340;
    wire N__39335;
    wire N__39332;
    wire N__39331;
    wire N__39328;
    wire N__39325;
    wire N__39320;
    wire N__39317;
    wire N__39314;
    wire N__39313;
    wire N__39308;
    wire N__39307;
    wire N__39304;
    wire N__39301;
    wire N__39300;
    wire N__39297;
    wire N__39294;
    wire N__39291;
    wire N__39290;
    wire N__39287;
    wire N__39286;
    wire N__39285;
    wire N__39282;
    wire N__39279;
    wire N__39276;
    wire N__39273;
    wire N__39270;
    wire N__39267;
    wire N__39262;
    wire N__39251;
    wire N__39248;
    wire N__39245;
    wire N__39242;
    wire N__39241;
    wire N__39240;
    wire N__39237;
    wire N__39236;
    wire N__39231;
    wire N__39230;
    wire N__39229;
    wire N__39228;
    wire N__39225;
    wire N__39222;
    wire N__39219;
    wire N__39216;
    wire N__39211;
    wire N__39206;
    wire N__39203;
    wire N__39194;
    wire N__39191;
    wire N__39190;
    wire N__39187;
    wire N__39184;
    wire N__39179;
    wire N__39176;
    wire N__39175;
    wire N__39172;
    wire N__39169;
    wire N__39164;
    wire N__39161;
    wire N__39160;
    wire N__39157;
    wire N__39154;
    wire N__39151;
    wire N__39148;
    wire N__39143;
    wire N__39140;
    wire N__39137;
    wire N__39134;
    wire N__39131;
    wire N__39130;
    wire N__39127;
    wire N__39126;
    wire N__39125;
    wire N__39124;
    wire N__39123;
    wire N__39122;
    wire N__39119;
    wire N__39116;
    wire N__39113;
    wire N__39108;
    wire N__39107;
    wire N__39104;
    wire N__39101;
    wire N__39096;
    wire N__39091;
    wire N__39086;
    wire N__39077;
    wire N__39074;
    wire N__39071;
    wire N__39068;
    wire N__39065;
    wire N__39064;
    wire N__39061;
    wire N__39058;
    wire N__39053;
    wire N__39052;
    wire N__39049;
    wire N__39046;
    wire N__39041;
    wire N__39040;
    wire N__39037;
    wire N__39034;
    wire N__39029;
    wire N__39028;
    wire N__39023;
    wire N__39020;
    wire N__39019;
    wire N__39016;
    wire N__39013;
    wire N__39008;
    wire N__39007;
    wire N__39002;
    wire N__38999;
    wire N__38996;
    wire N__38993;
    wire N__38990;
    wire N__38987;
    wire N__38984;
    wire N__38983;
    wire N__38980;
    wire N__38977;
    wire N__38972;
    wire N__38969;
    wire N__38966;
    wire N__38965;
    wire N__38962;
    wire N__38959;
    wire N__38954;
    wire N__38951;
    wire N__38950;
    wire N__38947;
    wire N__38944;
    wire N__38943;
    wire N__38940;
    wire N__38937;
    wire N__38934;
    wire N__38927;
    wire N__38926;
    wire N__38925;
    wire N__38922;
    wire N__38919;
    wire N__38918;
    wire N__38915;
    wire N__38912;
    wire N__38907;
    wire N__38906;
    wire N__38905;
    wire N__38902;
    wire N__38899;
    wire N__38896;
    wire N__38893;
    wire N__38890;
    wire N__38887;
    wire N__38880;
    wire N__38873;
    wire N__38872;
    wire N__38869;
    wire N__38866;
    wire N__38861;
    wire N__38860;
    wire N__38855;
    wire N__38852;
    wire N__38851;
    wire N__38846;
    wire N__38843;
    wire N__38842;
    wire N__38839;
    wire N__38836;
    wire N__38833;
    wire N__38828;
    wire N__38825;
    wire N__38824;
    wire N__38821;
    wire N__38818;
    wire N__38813;
    wire N__38810;
    wire N__38807;
    wire N__38804;
    wire N__38801;
    wire N__38800;
    wire N__38797;
    wire N__38794;
    wire N__38791;
    wire N__38790;
    wire N__38787;
    wire N__38784;
    wire N__38781;
    wire N__38778;
    wire N__38775;
    wire N__38768;
    wire N__38765;
    wire N__38762;
    wire N__38761;
    wire N__38758;
    wire N__38755;
    wire N__38752;
    wire N__38749;
    wire N__38744;
    wire N__38743;
    wire N__38740;
    wire N__38737;
    wire N__38732;
    wire N__38729;
    wire N__38726;
    wire N__38725;
    wire N__38722;
    wire N__38719;
    wire N__38714;
    wire N__38713;
    wire N__38710;
    wire N__38707;
    wire N__38702;
    wire N__38701;
    wire N__38696;
    wire N__38693;
    wire N__38690;
    wire N__38687;
    wire N__38684;
    wire N__38681;
    wire N__38678;
    wire N__38675;
    wire N__38672;
    wire N__38671;
    wire N__38668;
    wire N__38665;
    wire N__38660;
    wire N__38657;
    wire N__38654;
    wire N__38651;
    wire N__38648;
    wire N__38645;
    wire N__38642;
    wire N__38639;
    wire N__38636;
    wire N__38633;
    wire N__38630;
    wire N__38627;
    wire N__38626;
    wire N__38623;
    wire N__38620;
    wire N__38615;
    wire N__38612;
    wire N__38609;
    wire N__38608;
    wire N__38605;
    wire N__38602;
    wire N__38597;
    wire N__38596;
    wire N__38591;
    wire N__38588;
    wire N__38587;
    wire N__38582;
    wire N__38579;
    wire N__38578;
    wire N__38573;
    wire N__38570;
    wire N__38569;
    wire N__38566;
    wire N__38563;
    wire N__38558;
    wire N__38557;
    wire N__38554;
    wire N__38551;
    wire N__38546;
    wire N__38543;
    wire N__38540;
    wire N__38537;
    wire N__38536;
    wire N__38533;
    wire N__38530;
    wire N__38525;
    wire N__38524;
    wire N__38521;
    wire N__38518;
    wire N__38513;
    wire N__38510;
    wire N__38507;
    wire N__38506;
    wire N__38503;
    wire N__38500;
    wire N__38497;
    wire N__38494;
    wire N__38493;
    wire N__38490;
    wire N__38487;
    wire N__38484;
    wire N__38477;
    wire N__38474;
    wire N__38471;
    wire N__38468;
    wire N__38465;
    wire N__38464;
    wire N__38461;
    wire N__38458;
    wire N__38453;
    wire N__38450;
    wire N__38447;
    wire N__38444;
    wire N__38443;
    wire N__38440;
    wire N__38437;
    wire N__38432;
    wire N__38431;
    wire N__38426;
    wire N__38423;
    wire N__38422;
    wire N__38417;
    wire N__38414;
    wire N__38413;
    wire N__38408;
    wire N__38405;
    wire N__38402;
    wire N__38399;
    wire N__38398;
    wire N__38395;
    wire N__38392;
    wire N__38389;
    wire N__38384;
    wire N__38381;
    wire N__38378;
    wire N__38377;
    wire N__38374;
    wire N__38371;
    wire N__38368;
    wire N__38365;
    wire N__38364;
    wire N__38361;
    wire N__38358;
    wire N__38355;
    wire N__38348;
    wire N__38347;
    wire N__38346;
    wire N__38343;
    wire N__38338;
    wire N__38335;
    wire N__38330;
    wire N__38327;
    wire N__38326;
    wire N__38325;
    wire N__38322;
    wire N__38317;
    wire N__38314;
    wire N__38309;
    wire N__38308;
    wire N__38303;
    wire N__38300;
    wire N__38297;
    wire N__38294;
    wire N__38291;
    wire N__38288;
    wire N__38285;
    wire N__38282;
    wire N__38281;
    wire N__38278;
    wire N__38275;
    wire N__38272;
    wire N__38267;
    wire N__38264;
    wire N__38263;
    wire N__38260;
    wire N__38257;
    wire N__38252;
    wire N__38249;
    wire N__38248;
    wire N__38245;
    wire N__38242;
    wire N__38239;
    wire N__38234;
    wire N__38231;
    wire N__38228;
    wire N__38227;
    wire N__38224;
    wire N__38221;
    wire N__38216;
    wire N__38215;
    wire N__38212;
    wire N__38209;
    wire N__38206;
    wire N__38201;
    wire N__38200;
    wire N__38195;
    wire N__38192;
    wire N__38191;
    wire N__38188;
    wire N__38185;
    wire N__38182;
    wire N__38177;
    wire N__38176;
    wire N__38173;
    wire N__38170;
    wire N__38167;
    wire N__38164;
    wire N__38159;
    wire N__38156;
    wire N__38155;
    wire N__38152;
    wire N__38149;
    wire N__38146;
    wire N__38141;
    wire N__38140;
    wire N__38137;
    wire N__38134;
    wire N__38131;
    wire N__38126;
    wire N__38125;
    wire N__38122;
    wire N__38119;
    wire N__38116;
    wire N__38111;
    wire N__38110;
    wire N__38107;
    wire N__38106;
    wire N__38103;
    wire N__38102;
    wire N__38101;
    wire N__38100;
    wire N__38097;
    wire N__38096;
    wire N__38093;
    wire N__38090;
    wire N__38087;
    wire N__38084;
    wire N__38081;
    wire N__38078;
    wire N__38073;
    wire N__38060;
    wire N__38057;
    wire N__38056;
    wire N__38055;
    wire N__38054;
    wire N__38051;
    wire N__38050;
    wire N__38049;
    wire N__38046;
    wire N__38043;
    wire N__38040;
    wire N__38037;
    wire N__38032;
    wire N__38021;
    wire N__38020;
    wire N__38017;
    wire N__38014;
    wire N__38011;
    wire N__38008;
    wire N__38005;
    wire N__38000;
    wire N__37999;
    wire N__37998;
    wire N__37997;
    wire N__37994;
    wire N__37993;
    wire N__37992;
    wire N__37989;
    wire N__37986;
    wire N__37983;
    wire N__37980;
    wire N__37975;
    wire N__37964;
    wire N__37961;
    wire N__37958;
    wire N__37955;
    wire N__37952;
    wire N__37949;
    wire N__37946;
    wire N__37945;
    wire N__37942;
    wire N__37941;
    wire N__37938;
    wire N__37933;
    wire N__37930;
    wire N__37927;
    wire N__37922;
    wire N__37919;
    wire N__37918;
    wire N__37917;
    wire N__37916;
    wire N__37915;
    wire N__37914;
    wire N__37911;
    wire N__37910;
    wire N__37909;
    wire N__37902;
    wire N__37899;
    wire N__37896;
    wire N__37895;
    wire N__37894;
    wire N__37891;
    wire N__37888;
    wire N__37885;
    wire N__37882;
    wire N__37877;
    wire N__37876;
    wire N__37873;
    wire N__37870;
    wire N__37867;
    wire N__37862;
    wire N__37859;
    wire N__37856;
    wire N__37851;
    wire N__37838;
    wire N__37835;
    wire N__37834;
    wire N__37831;
    wire N__37828;
    wire N__37823;
    wire N__37820;
    wire N__37819;
    wire N__37816;
    wire N__37813;
    wire N__37808;
    wire N__37805;
    wire N__37804;
    wire N__37801;
    wire N__37798;
    wire N__37793;
    wire N__37792;
    wire N__37787;
    wire N__37784;
    wire N__37781;
    wire N__37778;
    wire N__37775;
    wire N__37774;
    wire N__37771;
    wire N__37768;
    wire N__37763;
    wire N__37762;
    wire N__37757;
    wire N__37754;
    wire N__37753;
    wire N__37750;
    wire N__37747;
    wire N__37744;
    wire N__37739;
    wire N__37738;
    wire N__37735;
    wire N__37732;
    wire N__37729;
    wire N__37726;
    wire N__37721;
    wire N__37718;
    wire N__37717;
    wire N__37714;
    wire N__37711;
    wire N__37706;
    wire N__37703;
    wire N__37702;
    wire N__37699;
    wire N__37696;
    wire N__37691;
    wire N__37690;
    wire N__37685;
    wire N__37682;
    wire N__37679;
    wire N__37676;
    wire N__37673;
    wire N__37670;
    wire N__37667;
    wire N__37664;
    wire N__37661;
    wire N__37660;
    wire N__37657;
    wire N__37656;
    wire N__37653;
    wire N__37652;
    wire N__37649;
    wire N__37648;
    wire N__37645;
    wire N__37642;
    wire N__37639;
    wire N__37636;
    wire N__37633;
    wire N__37630;
    wire N__37625;
    wire N__37616;
    wire N__37613;
    wire N__37612;
    wire N__37609;
    wire N__37608;
    wire N__37605;
    wire N__37604;
    wire N__37601;
    wire N__37598;
    wire N__37595;
    wire N__37592;
    wire N__37589;
    wire N__37586;
    wire N__37583;
    wire N__37574;
    wire N__37573;
    wire N__37570;
    wire N__37567;
    wire N__37566;
    wire N__37563;
    wire N__37560;
    wire N__37557;
    wire N__37554;
    wire N__37553;
    wire N__37552;
    wire N__37547;
    wire N__37544;
    wire N__37541;
    wire N__37538;
    wire N__37533;
    wire N__37530;
    wire N__37523;
    wire N__37520;
    wire N__37519;
    wire N__37518;
    wire N__37515;
    wire N__37512;
    wire N__37509;
    wire N__37508;
    wire N__37507;
    wire N__37504;
    wire N__37501;
    wire N__37498;
    wire N__37495;
    wire N__37492;
    wire N__37489;
    wire N__37486;
    wire N__37481;
    wire N__37472;
    wire N__37469;
    wire N__37466;
    wire N__37463;
    wire N__37460;
    wire N__37457;
    wire N__37454;
    wire N__37453;
    wire N__37450;
    wire N__37447;
    wire N__37442;
    wire N__37441;
    wire N__37440;
    wire N__37437;
    wire N__37434;
    wire N__37431;
    wire N__37428;
    wire N__37425;
    wire N__37418;
    wire N__37417;
    wire N__37414;
    wire N__37411;
    wire N__37408;
    wire N__37403;
    wire N__37402;
    wire N__37399;
    wire N__37398;
    wire N__37397;
    wire N__37396;
    wire N__37395;
    wire N__37390;
    wire N__37385;
    wire N__37382;
    wire N__37379;
    wire N__37376;
    wire N__37373;
    wire N__37364;
    wire N__37363;
    wire N__37362;
    wire N__37359;
    wire N__37354;
    wire N__37351;
    wire N__37346;
    wire N__37343;
    wire N__37340;
    wire N__37337;
    wire N__37334;
    wire N__37331;
    wire N__37328;
    wire N__37325;
    wire N__37322;
    wire N__37321;
    wire N__37320;
    wire N__37319;
    wire N__37316;
    wire N__37315;
    wire N__37312;
    wire N__37309;
    wire N__37306;
    wire N__37303;
    wire N__37300;
    wire N__37295;
    wire N__37286;
    wire N__37283;
    wire N__37280;
    wire N__37277;
    wire N__37274;
    wire N__37273;
    wire N__37268;
    wire N__37265;
    wire N__37262;
    wire N__37261;
    wire N__37258;
    wire N__37255;
    wire N__37254;
    wire N__37253;
    wire N__37252;
    wire N__37249;
    wire N__37246;
    wire N__37241;
    wire N__37238;
    wire N__37229;
    wire N__37226;
    wire N__37223;
    wire N__37222;
    wire N__37219;
    wire N__37216;
    wire N__37215;
    wire N__37210;
    wire N__37209;
    wire N__37206;
    wire N__37203;
    wire N__37200;
    wire N__37199;
    wire N__37192;
    wire N__37189;
    wire N__37186;
    wire N__37181;
    wire N__37178;
    wire N__37175;
    wire N__37172;
    wire N__37169;
    wire N__37166;
    wire N__37163;
    wire N__37162;
    wire N__37159;
    wire N__37156;
    wire N__37151;
    wire N__37148;
    wire N__37145;
    wire N__37144;
    wire N__37141;
    wire N__37138;
    wire N__37133;
    wire N__37132;
    wire N__37129;
    wire N__37126;
    wire N__37121;
    wire N__37118;
    wire N__37117;
    wire N__37114;
    wire N__37111;
    wire N__37106;
    wire N__37103;
    wire N__37102;
    wire N__37099;
    wire N__37096;
    wire N__37091;
    wire N__37088;
    wire N__37087;
    wire N__37084;
    wire N__37081;
    wire N__37076;
    wire N__37075;
    wire N__37070;
    wire N__37067;
    wire N__37066;
    wire N__37063;
    wire N__37060;
    wire N__37055;
    wire N__37052;
    wire N__37049;
    wire N__37046;
    wire N__37043;
    wire N__37042;
    wire N__37039;
    wire N__37036;
    wire N__37033;
    wire N__37032;
    wire N__37029;
    wire N__37026;
    wire N__37023;
    wire N__37016;
    wire N__37015;
    wire N__37012;
    wire N__37009;
    wire N__37008;
    wire N__37005;
    wire N__37002;
    wire N__36999;
    wire N__36996;
    wire N__36989;
    wire N__36986;
    wire N__36983;
    wire N__36982;
    wire N__36979;
    wire N__36978;
    wire N__36975;
    wire N__36972;
    wire N__36969;
    wire N__36962;
    wire N__36961;
    wire N__36958;
    wire N__36955;
    wire N__36952;
    wire N__36949;
    wire N__36948;
    wire N__36947;
    wire N__36944;
    wire N__36941;
    wire N__36938;
    wire N__36935;
    wire N__36930;
    wire N__36923;
    wire N__36920;
    wire N__36917;
    wire N__36916;
    wire N__36913;
    wire N__36912;
    wire N__36909;
    wire N__36906;
    wire N__36903;
    wire N__36902;
    wire N__36899;
    wire N__36896;
    wire N__36893;
    wire N__36890;
    wire N__36887;
    wire N__36884;
    wire N__36881;
    wire N__36872;
    wire N__36871;
    wire N__36868;
    wire N__36865;
    wire N__36862;
    wire N__36859;
    wire N__36858;
    wire N__36857;
    wire N__36852;
    wire N__36849;
    wire N__36846;
    wire N__36843;
    wire N__36836;
    wire N__36833;
    wire N__36832;
    wire N__36831;
    wire N__36828;
    wire N__36825;
    wire N__36822;
    wire N__36819;
    wire N__36814;
    wire N__36811;
    wire N__36806;
    wire N__36803;
    wire N__36800;
    wire N__36797;
    wire N__36794;
    wire N__36791;
    wire N__36788;
    wire N__36785;
    wire N__36782;
    wire N__36779;
    wire N__36778;
    wire N__36775;
    wire N__36772;
    wire N__36767;
    wire N__36764;
    wire N__36761;
    wire N__36758;
    wire N__36755;
    wire N__36754;
    wire N__36751;
    wire N__36748;
    wire N__36743;
    wire N__36742;
    wire N__36741;
    wire N__36736;
    wire N__36733;
    wire N__36730;
    wire N__36729;
    wire N__36726;
    wire N__36723;
    wire N__36720;
    wire N__36717;
    wire N__36714;
    wire N__36711;
    wire N__36708;
    wire N__36705;
    wire N__36702;
    wire N__36699;
    wire N__36692;
    wire N__36691;
    wire N__36690;
    wire N__36687;
    wire N__36686;
    wire N__36685;
    wire N__36682;
    wire N__36679;
    wire N__36676;
    wire N__36673;
    wire N__36670;
    wire N__36667;
    wire N__36664;
    wire N__36659;
    wire N__36656;
    wire N__36653;
    wire N__36650;
    wire N__36645;
    wire N__36642;
    wire N__36637;
    wire N__36632;
    wire N__36631;
    wire N__36626;
    wire N__36625;
    wire N__36624;
    wire N__36621;
    wire N__36618;
    wire N__36615;
    wire N__36612;
    wire N__36609;
    wire N__36606;
    wire N__36601;
    wire N__36598;
    wire N__36597;
    wire N__36594;
    wire N__36591;
    wire N__36588;
    wire N__36581;
    wire N__36580;
    wire N__36579;
    wire N__36576;
    wire N__36573;
    wire N__36568;
    wire N__36565;
    wire N__36562;
    wire N__36557;
    wire N__36556;
    wire N__36553;
    wire N__36548;
    wire N__36547;
    wire N__36544;
    wire N__36541;
    wire N__36538;
    wire N__36535;
    wire N__36532;
    wire N__36529;
    wire N__36524;
    wire N__36523;
    wire N__36520;
    wire N__36517;
    wire N__36516;
    wire N__36513;
    wire N__36510;
    wire N__36507;
    wire N__36504;
    wire N__36497;
    wire N__36494;
    wire N__36493;
    wire N__36492;
    wire N__36489;
    wire N__36486;
    wire N__36483;
    wire N__36480;
    wire N__36477;
    wire N__36470;
    wire N__36467;
    wire N__36464;
    wire N__36463;
    wire N__36460;
    wire N__36459;
    wire N__36458;
    wire N__36455;
    wire N__36452;
    wire N__36449;
    wire N__36446;
    wire N__36443;
    wire N__36438;
    wire N__36437;
    wire N__36434;
    wire N__36431;
    wire N__36428;
    wire N__36425;
    wire N__36422;
    wire N__36413;
    wire N__36410;
    wire N__36409;
    wire N__36408;
    wire N__36403;
    wire N__36400;
    wire N__36399;
    wire N__36396;
    wire N__36393;
    wire N__36390;
    wire N__36387;
    wire N__36384;
    wire N__36383;
    wire N__36380;
    wire N__36377;
    wire N__36374;
    wire N__36371;
    wire N__36368;
    wire N__36359;
    wire N__36356;
    wire N__36355;
    wire N__36354;
    wire N__36353;
    wire N__36348;
    wire N__36345;
    wire N__36342;
    wire N__36339;
    wire N__36336;
    wire N__36335;
    wire N__36332;
    wire N__36329;
    wire N__36326;
    wire N__36323;
    wire N__36320;
    wire N__36311;
    wire N__36308;
    wire N__36307;
    wire N__36306;
    wire N__36301;
    wire N__36298;
    wire N__36297;
    wire N__36294;
    wire N__36291;
    wire N__36288;
    wire N__36287;
    wire N__36284;
    wire N__36281;
    wire N__36278;
    wire N__36275;
    wire N__36268;
    wire N__36263;
    wire N__36260;
    wire N__36259;
    wire N__36256;
    wire N__36253;
    wire N__36250;
    wire N__36247;
    wire N__36244;
    wire N__36243;
    wire N__36242;
    wire N__36239;
    wire N__36236;
    wire N__36231;
    wire N__36224;
    wire N__36223;
    wire N__36220;
    wire N__36217;
    wire N__36214;
    wire N__36211;
    wire N__36210;
    wire N__36207;
    wire N__36204;
    wire N__36201;
    wire N__36196;
    wire N__36191;
    wire N__36190;
    wire N__36187;
    wire N__36184;
    wire N__36181;
    wire N__36178;
    wire N__36177;
    wire N__36174;
    wire N__36171;
    wire N__36168;
    wire N__36165;
    wire N__36162;
    wire N__36155;
    wire N__36152;
    wire N__36151;
    wire N__36148;
    wire N__36145;
    wire N__36144;
    wire N__36143;
    wire N__36138;
    wire N__36135;
    wire N__36132;
    wire N__36131;
    wire N__36128;
    wire N__36125;
    wire N__36122;
    wire N__36119;
    wire N__36114;
    wire N__36107;
    wire N__36104;
    wire N__36101;
    wire N__36100;
    wire N__36099;
    wire N__36098;
    wire N__36095;
    wire N__36092;
    wire N__36089;
    wire N__36086;
    wire N__36083;
    wire N__36080;
    wire N__36077;
    wire N__36076;
    wire N__36073;
    wire N__36070;
    wire N__36067;
    wire N__36064;
    wire N__36061;
    wire N__36058;
    wire N__36047;
    wire N__36044;
    wire N__36043;
    wire N__36042;
    wire N__36035;
    wire N__36034;
    wire N__36031;
    wire N__36028;
    wire N__36027;
    wire N__36024;
    wire N__36021;
    wire N__36018;
    wire N__36013;
    wire N__36008;
    wire N__36005;
    wire N__36004;
    wire N__36003;
    wire N__36000;
    wire N__35995;
    wire N__35992;
    wire N__35991;
    wire N__35988;
    wire N__35985;
    wire N__35982;
    wire N__35979;
    wire N__35978;
    wire N__35975;
    wire N__35972;
    wire N__35969;
    wire N__35966;
    wire N__35961;
    wire N__35954;
    wire N__35951;
    wire N__35950;
    wire N__35949;
    wire N__35946;
    wire N__35943;
    wire N__35940;
    wire N__35939;
    wire N__35936;
    wire N__35933;
    wire N__35930;
    wire N__35927;
    wire N__35924;
    wire N__35921;
    wire N__35920;
    wire N__35917;
    wire N__35914;
    wire N__35911;
    wire N__35908;
    wire N__35905;
    wire N__35900;
    wire N__35891;
    wire N__35888;
    wire N__35887;
    wire N__35886;
    wire N__35883;
    wire N__35880;
    wire N__35877;
    wire N__35874;
    wire N__35871;
    wire N__35868;
    wire N__35867;
    wire N__35864;
    wire N__35861;
    wire N__35860;
    wire N__35857;
    wire N__35854;
    wire N__35851;
    wire N__35848;
    wire N__35845;
    wire N__35840;
    wire N__35831;
    wire N__35828;
    wire N__35825;
    wire N__35822;
    wire N__35821;
    wire N__35818;
    wire N__35815;
    wire N__35810;
    wire N__35809;
    wire N__35806;
    wire N__35803;
    wire N__35802;
    wire N__35797;
    wire N__35796;
    wire N__35793;
    wire N__35790;
    wire N__35787;
    wire N__35784;
    wire N__35777;
    wire N__35774;
    wire N__35771;
    wire N__35770;
    wire N__35769;
    wire N__35766;
    wire N__35763;
    wire N__35760;
    wire N__35759;
    wire N__35756;
    wire N__35753;
    wire N__35750;
    wire N__35749;
    wire N__35746;
    wire N__35743;
    wire N__35740;
    wire N__35737;
    wire N__35734;
    wire N__35731;
    wire N__35720;
    wire N__35717;
    wire N__35716;
    wire N__35715;
    wire N__35710;
    wire N__35707;
    wire N__35706;
    wire N__35701;
    wire N__35698;
    wire N__35693;
    wire N__35690;
    wire N__35689;
    wire N__35686;
    wire N__35685;
    wire N__35682;
    wire N__35679;
    wire N__35676;
    wire N__35673;
    wire N__35666;
    wire N__35663;
    wire N__35662;
    wire N__35659;
    wire N__35658;
    wire N__35657;
    wire N__35654;
    wire N__35651;
    wire N__35648;
    wire N__35647;
    wire N__35644;
    wire N__35641;
    wire N__35636;
    wire N__35633;
    wire N__35632;
    wire N__35629;
    wire N__35626;
    wire N__35621;
    wire N__35618;
    wire N__35615;
    wire N__35606;
    wire N__35603;
    wire N__35602;
    wire N__35601;
    wire N__35596;
    wire N__35595;
    wire N__35592;
    wire N__35589;
    wire N__35586;
    wire N__35585;
    wire N__35582;
    wire N__35579;
    wire N__35576;
    wire N__35573;
    wire N__35570;
    wire N__35567;
    wire N__35564;
    wire N__35563;
    wire N__35560;
    wire N__35557;
    wire N__35552;
    wire N__35549;
    wire N__35546;
    wire N__35537;
    wire N__35534;
    wire N__35533;
    wire N__35532;
    wire N__35529;
    wire N__35524;
    wire N__35523;
    wire N__35522;
    wire N__35519;
    wire N__35516;
    wire N__35513;
    wire N__35510;
    wire N__35507;
    wire N__35504;
    wire N__35503;
    wire N__35500;
    wire N__35497;
    wire N__35492;
    wire N__35489;
    wire N__35484;
    wire N__35477;
    wire N__35474;
    wire N__35471;
    wire N__35468;
    wire N__35467;
    wire N__35464;
    wire N__35461;
    wire N__35460;
    wire N__35459;
    wire N__35458;
    wire N__35455;
    wire N__35452;
    wire N__35449;
    wire N__35446;
    wire N__35443;
    wire N__35438;
    wire N__35437;
    wire N__35432;
    wire N__35429;
    wire N__35426;
    wire N__35423;
    wire N__35418;
    wire N__35411;
    wire N__35408;
    wire N__35407;
    wire N__35406;
    wire N__35403;
    wire N__35400;
    wire N__35397;
    wire N__35396;
    wire N__35393;
    wire N__35390;
    wire N__35387;
    wire N__35386;
    wire N__35383;
    wire N__35380;
    wire N__35375;
    wire N__35372;
    wire N__35369;
    wire N__35360;
    wire N__35357;
    wire N__35356;
    wire N__35355;
    wire N__35352;
    wire N__35349;
    wire N__35346;
    wire N__35345;
    wire N__35342;
    wire N__35339;
    wire N__35336;
    wire N__35335;
    wire N__35332;
    wire N__35329;
    wire N__35324;
    wire N__35321;
    wire N__35318;
    wire N__35309;
    wire N__35306;
    wire N__35305;
    wire N__35302;
    wire N__35299;
    wire N__35298;
    wire N__35293;
    wire N__35290;
    wire N__35289;
    wire N__35284;
    wire N__35283;
    wire N__35280;
    wire N__35277;
    wire N__35274;
    wire N__35271;
    wire N__35264;
    wire N__35261;
    wire N__35260;
    wire N__35257;
    wire N__35254;
    wire N__35251;
    wire N__35250;
    wire N__35249;
    wire N__35246;
    wire N__35243;
    wire N__35240;
    wire N__35239;
    wire N__35236;
    wire N__35233;
    wire N__35228;
    wire N__35225;
    wire N__35222;
    wire N__35213;
    wire N__35210;
    wire N__35209;
    wire N__35206;
    wire N__35205;
    wire N__35204;
    wire N__35201;
    wire N__35198;
    wire N__35195;
    wire N__35194;
    wire N__35191;
    wire N__35190;
    wire N__35187;
    wire N__35184;
    wire N__35181;
    wire N__35178;
    wire N__35175;
    wire N__35172;
    wire N__35165;
    wire N__35156;
    wire N__35153;
    wire N__35150;
    wire N__35149;
    wire N__35146;
    wire N__35143;
    wire N__35140;
    wire N__35139;
    wire N__35138;
    wire N__35137;
    wire N__35134;
    wire N__35133;
    wire N__35130;
    wire N__35127;
    wire N__35122;
    wire N__35119;
    wire N__35116;
    wire N__35111;
    wire N__35102;
    wire N__35099;
    wire N__35098;
    wire N__35097;
    wire N__35094;
    wire N__35093;
    wire N__35088;
    wire N__35087;
    wire N__35084;
    wire N__35081;
    wire N__35078;
    wire N__35075;
    wire N__35072;
    wire N__35071;
    wire N__35066;
    wire N__35063;
    wire N__35060;
    wire N__35057;
    wire N__35052;
    wire N__35045;
    wire N__35042;
    wire N__35041;
    wire N__35040;
    wire N__35039;
    wire N__35036;
    wire N__35033;
    wire N__35030;
    wire N__35029;
    wire N__35026;
    wire N__35023;
    wire N__35020;
    wire N__35017;
    wire N__35014;
    wire N__35013;
    wire N__35010;
    wire N__35007;
    wire N__35002;
    wire N__34999;
    wire N__34996;
    wire N__34993;
    wire N__34982;
    wire N__34979;
    wire N__34978;
    wire N__34975;
    wire N__34972;
    wire N__34967;
    wire N__34964;
    wire N__34963;
    wire N__34960;
    wire N__34957;
    wire N__34956;
    wire N__34955;
    wire N__34952;
    wire N__34951;
    wire N__34948;
    wire N__34945;
    wire N__34942;
    wire N__34939;
    wire N__34938;
    wire N__34935;
    wire N__34932;
    wire N__34927;
    wire N__34924;
    wire N__34921;
    wire N__34918;
    wire N__34907;
    wire N__34906;
    wire N__34903;
    wire N__34900;
    wire N__34897;
    wire N__34894;
    wire N__34889;
    wire N__34886;
    wire N__34885;
    wire N__34884;
    wire N__34881;
    wire N__34880;
    wire N__34877;
    wire N__34874;
    wire N__34871;
    wire N__34868;
    wire N__34867;
    wire N__34862;
    wire N__34857;
    wire N__34856;
    wire N__34853;
    wire N__34850;
    wire N__34847;
    wire N__34844;
    wire N__34841;
    wire N__34832;
    wire N__34829;
    wire N__34826;
    wire N__34825;
    wire N__34824;
    wire N__34821;
    wire N__34818;
    wire N__34817;
    wire N__34814;
    wire N__34813;
    wire N__34808;
    wire N__34805;
    wire N__34802;
    wire N__34801;
    wire N__34798;
    wire N__34795;
    wire N__34792;
    wire N__34789;
    wire N__34786;
    wire N__34783;
    wire N__34772;
    wire N__34769;
    wire N__34766;
    wire N__34765;
    wire N__34764;
    wire N__34761;
    wire N__34758;
    wire N__34757;
    wire N__34754;
    wire N__34749;
    wire N__34746;
    wire N__34745;
    wire N__34742;
    wire N__34737;
    wire N__34736;
    wire N__34733;
    wire N__34730;
    wire N__34727;
    wire N__34724;
    wire N__34721;
    wire N__34712;
    wire N__34709;
    wire N__34706;
    wire N__34705;
    wire N__34702;
    wire N__34699;
    wire N__34694;
    wire N__34693;
    wire N__34688;
    wire N__34685;
    wire N__34684;
    wire N__34683;
    wire N__34680;
    wire N__34679;
    wire N__34676;
    wire N__34675;
    wire N__34674;
    wire N__34673;
    wire N__34672;
    wire N__34669;
    wire N__34666;
    wire N__34663;
    wire N__34662;
    wire N__34661;
    wire N__34660;
    wire N__34659;
    wire N__34656;
    wire N__34653;
    wire N__34648;
    wire N__34645;
    wire N__34644;
    wire N__34643;
    wire N__34642;
    wire N__34641;
    wire N__34640;
    wire N__34637;
    wire N__34632;
    wire N__34629;
    wire N__34628;
    wire N__34627;
    wire N__34626;
    wire N__34623;
    wire N__34622;
    wire N__34619;
    wire N__34616;
    wire N__34607;
    wire N__34606;
    wire N__34605;
    wire N__34602;
    wire N__34601;
    wire N__34598;
    wire N__34595;
    wire N__34594;
    wire N__34589;
    wire N__34582;
    wire N__34577;
    wire N__34576;
    wire N__34575;
    wire N__34574;
    wire N__34573;
    wire N__34572;
    wire N__34571;
    wire N__34570;
    wire N__34569;
    wire N__34562;
    wire N__34555;
    wire N__34554;
    wire N__34553;
    wire N__34552;
    wire N__34551;
    wire N__34550;
    wire N__34549;
    wire N__34548;
    wire N__34545;
    wire N__34542;
    wire N__34537;
    wire N__34534;
    wire N__34529;
    wire N__34522;
    wire N__34515;
    wire N__34510;
    wire N__34503;
    wire N__34498;
    wire N__34491;
    wire N__34482;
    wire N__34457;
    wire N__34456;
    wire N__34455;
    wire N__34454;
    wire N__34453;
    wire N__34452;
    wire N__34449;
    wire N__34448;
    wire N__34447;
    wire N__34446;
    wire N__34445;
    wire N__34444;
    wire N__34437;
    wire N__34436;
    wire N__34435;
    wire N__34434;
    wire N__34433;
    wire N__34430;
    wire N__34427;
    wire N__34426;
    wire N__34423;
    wire N__34420;
    wire N__34417;
    wire N__34414;
    wire N__34409;
    wire N__34408;
    wire N__34405;
    wire N__34400;
    wire N__34395;
    wire N__34394;
    wire N__34393;
    wire N__34390;
    wire N__34387;
    wire N__34384;
    wire N__34379;
    wire N__34376;
    wire N__34371;
    wire N__34368;
    wire N__34367;
    wire N__34362;
    wire N__34359;
    wire N__34354;
    wire N__34341;
    wire N__34336;
    wire N__34325;
    wire N__34322;
    wire N__34319;
    wire N__34318;
    wire N__34315;
    wire N__34312;
    wire N__34309;
    wire N__34308;
    wire N__34307;
    wire N__34304;
    wire N__34301;
    wire N__34296;
    wire N__34289;
    wire N__34288;
    wire N__34285;
    wire N__34282;
    wire N__34279;
    wire N__34276;
    wire N__34273;
    wire N__34268;
    wire N__34265;
    wire N__34264;
    wire N__34261;
    wire N__34258;
    wire N__34253;
    wire N__34250;
    wire N__34247;
    wire N__34246;
    wire N__34245;
    wire N__34242;
    wire N__34237;
    wire N__34232;
    wire N__34229;
    wire N__34226;
    wire N__34223;
    wire N__34220;
    wire N__34219;
    wire N__34214;
    wire N__34213;
    wire N__34212;
    wire N__34211;
    wire N__34208;
    wire N__34205;
    wire N__34202;
    wire N__34201;
    wire N__34198;
    wire N__34195;
    wire N__34192;
    wire N__34189;
    wire N__34186;
    wire N__34183;
    wire N__34180;
    wire N__34171;
    wire N__34166;
    wire N__34165;
    wire N__34164;
    wire N__34161;
    wire N__34160;
    wire N__34155;
    wire N__34152;
    wire N__34149;
    wire N__34148;
    wire N__34145;
    wire N__34140;
    wire N__34139;
    wire N__34136;
    wire N__34133;
    wire N__34130;
    wire N__34127;
    wire N__34124;
    wire N__34115;
    wire N__34112;
    wire N__34109;
    wire N__34108;
    wire N__34105;
    wire N__34102;
    wire N__34101;
    wire N__34100;
    wire N__34095;
    wire N__34092;
    wire N__34089;
    wire N__34088;
    wire N__34085;
    wire N__34082;
    wire N__34079;
    wire N__34078;
    wire N__34075;
    wire N__34070;
    wire N__34067;
    wire N__34064;
    wire N__34061;
    wire N__34052;
    wire N__34049;
    wire N__34046;
    wire N__34045;
    wire N__34042;
    wire N__34039;
    wire N__34034;
    wire N__34033;
    wire N__34030;
    wire N__34027;
    wire N__34024;
    wire N__34021;
    wire N__34018;
    wire N__34015;
    wire N__34012;
    wire N__34009;
    wire N__34006;
    wire N__34003;
    wire N__33998;
    wire N__33997;
    wire N__33994;
    wire N__33991;
    wire N__33988;
    wire N__33985;
    wire N__33980;
    wire N__33977;
    wire N__33976;
    wire N__33973;
    wire N__33970;
    wire N__33965;
    wire N__33962;
    wire N__33959;
    wire N__33956;
    wire N__33953;
    wire N__33952;
    wire N__33949;
    wire N__33946;
    wire N__33941;
    wire N__33938;
    wire N__33935;
    wire N__33932;
    wire N__33931;
    wire N__33928;
    wire N__33925;
    wire N__33924;
    wire N__33919;
    wire N__33916;
    wire N__33911;
    wire N__33910;
    wire N__33907;
    wire N__33904;
    wire N__33903;
    wire N__33902;
    wire N__33895;
    wire N__33892;
    wire N__33887;
    wire N__33884;
    wire N__33881;
    wire N__33878;
    wire N__33877;
    wire N__33874;
    wire N__33871;
    wire N__33866;
    wire N__33863;
    wire N__33860;
    wire N__33859;
    wire N__33856;
    wire N__33853;
    wire N__33852;
    wire N__33849;
    wire N__33846;
    wire N__33843;
    wire N__33840;
    wire N__33833;
    wire N__33832;
    wire N__33831;
    wire N__33828;
    wire N__33825;
    wire N__33822;
    wire N__33819;
    wire N__33814;
    wire N__33811;
    wire N__33808;
    wire N__33803;
    wire N__33800;
    wire N__33797;
    wire N__33794;
    wire N__33793;
    wire N__33790;
    wire N__33789;
    wire N__33786;
    wire N__33783;
    wire N__33780;
    wire N__33773;
    wire N__33770;
    wire N__33767;
    wire N__33764;
    wire N__33763;
    wire N__33760;
    wire N__33757;
    wire N__33754;
    wire N__33751;
    wire N__33750;
    wire N__33747;
    wire N__33744;
    wire N__33741;
    wire N__33738;
    wire N__33731;
    wire N__33728;
    wire N__33725;
    wire N__33724;
    wire N__33721;
    wire N__33718;
    wire N__33713;
    wire N__33710;
    wire N__33709;
    wire N__33706;
    wire N__33703;
    wire N__33698;
    wire N__33697;
    wire N__33694;
    wire N__33693;
    wire N__33692;
    wire N__33689;
    wire N__33686;
    wire N__33683;
    wire N__33682;
    wire N__33679;
    wire N__33678;
    wire N__33677;
    wire N__33674;
    wire N__33671;
    wire N__33668;
    wire N__33667;
    wire N__33666;
    wire N__33663;
    wire N__33660;
    wire N__33657;
    wire N__33654;
    wire N__33651;
    wire N__33646;
    wire N__33645;
    wire N__33640;
    wire N__33637;
    wire N__33634;
    wire N__33633;
    wire N__33630;
    wire N__33627;
    wire N__33622;
    wire N__33619;
    wire N__33614;
    wire N__33611;
    wire N__33608;
    wire N__33605;
    wire N__33600;
    wire N__33595;
    wire N__33592;
    wire N__33589;
    wire N__33586;
    wire N__33583;
    wire N__33580;
    wire N__33577;
    wire N__33572;
    wire N__33569;
    wire N__33560;
    wire N__33557;
    wire N__33554;
    wire N__33551;
    wire N__33548;
    wire N__33547;
    wire N__33544;
    wire N__33541;
    wire N__33538;
    wire N__33535;
    wire N__33530;
    wire N__33529;
    wire N__33526;
    wire N__33523;
    wire N__33522;
    wire N__33519;
    wire N__33518;
    wire N__33517;
    wire N__33516;
    wire N__33515;
    wire N__33514;
    wire N__33509;
    wire N__33508;
    wire N__33505;
    wire N__33498;
    wire N__33495;
    wire N__33492;
    wire N__33491;
    wire N__33488;
    wire N__33485;
    wire N__33480;
    wire N__33477;
    wire N__33474;
    wire N__33471;
    wire N__33468;
    wire N__33465;
    wire N__33462;
    wire N__33461;
    wire N__33460;
    wire N__33459;
    wire N__33456;
    wire N__33453;
    wire N__33448;
    wire N__33445;
    wire N__33442;
    wire N__33435;
    wire N__33428;
    wire N__33425;
    wire N__33422;
    wire N__33413;
    wire N__33410;
    wire N__33407;
    wire N__33404;
    wire N__33401;
    wire N__33398;
    wire N__33395;
    wire N__33392;
    wire N__33389;
    wire N__33388;
    wire N__33387;
    wire N__33384;
    wire N__33381;
    wire N__33380;
    wire N__33379;
    wire N__33378;
    wire N__33375;
    wire N__33368;
    wire N__33367;
    wire N__33364;
    wire N__33363;
    wire N__33360;
    wire N__33357;
    wire N__33354;
    wire N__33351;
    wire N__33346;
    wire N__33345;
    wire N__33342;
    wire N__33339;
    wire N__33336;
    wire N__33333;
    wire N__33330;
    wire N__33327;
    wire N__33326;
    wire N__33323;
    wire N__33322;
    wire N__33321;
    wire N__33320;
    wire N__33317;
    wire N__33312;
    wire N__33307;
    wire N__33304;
    wire N__33301;
    wire N__33296;
    wire N__33293;
    wire N__33288;
    wire N__33285;
    wire N__33272;
    wire N__33269;
    wire N__33268;
    wire N__33267;
    wire N__33266;
    wire N__33265;
    wire N__33262;
    wire N__33255;
    wire N__33252;
    wire N__33251;
    wire N__33250;
    wire N__33249;
    wire N__33246;
    wire N__33243;
    wire N__33242;
    wire N__33241;
    wire N__33238;
    wire N__33231;
    wire N__33230;
    wire N__33229;
    wire N__33226;
    wire N__33223;
    wire N__33218;
    wire N__33217;
    wire N__33214;
    wire N__33211;
    wire N__33208;
    wire N__33205;
    wire N__33200;
    wire N__33197;
    wire N__33194;
    wire N__33187;
    wire N__33182;
    wire N__33175;
    wire N__33170;
    wire N__33167;
    wire N__33166;
    wire N__33163;
    wire N__33160;
    wire N__33159;
    wire N__33158;
    wire N__33153;
    wire N__33150;
    wire N__33149;
    wire N__33148;
    wire N__33145;
    wire N__33140;
    wire N__33137;
    wire N__33134;
    wire N__33131;
    wire N__33126;
    wire N__33123;
    wire N__33120;
    wire N__33117;
    wire N__33114;
    wire N__33111;
    wire N__33108;
    wire N__33105;
    wire N__33098;
    wire N__33095;
    wire N__33092;
    wire N__33089;
    wire N__33086;
    wire N__33083;
    wire N__33080;
    wire N__33077;
    wire N__33074;
    wire N__33071;
    wire N__33068;
    wire N__33065;
    wire N__33062;
    wire N__33061;
    wire N__33060;
    wire N__33057;
    wire N__33054;
    wire N__33051;
    wire N__33048;
    wire N__33045;
    wire N__33038;
    wire N__33037;
    wire N__33034;
    wire N__33031;
    wire N__33028;
    wire N__33027;
    wire N__33024;
    wire N__33021;
    wire N__33018;
    wire N__33015;
    wire N__33014;
    wire N__33011;
    wire N__33008;
    wire N__33005;
    wire N__33002;
    wire N__32999;
    wire N__32994;
    wire N__32987;
    wire N__32986;
    wire N__32985;
    wire N__32984;
    wire N__32983;
    wire N__32980;
    wire N__32977;
    wire N__32974;
    wire N__32971;
    wire N__32968;
    wire N__32965;
    wire N__32962;
    wire N__32957;
    wire N__32952;
    wire N__32949;
    wire N__32946;
    wire N__32941;
    wire N__32936;
    wire N__32935;
    wire N__32932;
    wire N__32929;
    wire N__32924;
    wire N__32921;
    wire N__32920;
    wire N__32919;
    wire N__32912;
    wire N__32909;
    wire N__32908;
    wire N__32905;
    wire N__32902;
    wire N__32899;
    wire N__32896;
    wire N__32893;
    wire N__32892;
    wire N__32889;
    wire N__32886;
    wire N__32883;
    wire N__32880;
    wire N__32873;
    wire N__32870;
    wire N__32869;
    wire N__32866;
    wire N__32863;
    wire N__32858;
    wire N__32857;
    wire N__32852;
    wire N__32849;
    wire N__32846;
    wire N__32843;
    wire N__32842;
    wire N__32841;
    wire N__32838;
    wire N__32835;
    wire N__32834;
    wire N__32833;
    wire N__32832;
    wire N__32829;
    wire N__32828;
    wire N__32827;
    wire N__32826;
    wire N__32825;
    wire N__32824;
    wire N__32823;
    wire N__32822;
    wire N__32821;
    wire N__32820;
    wire N__32819;
    wire N__32818;
    wire N__32817;
    wire N__32816;
    wire N__32815;
    wire N__32814;
    wire N__32813;
    wire N__32812;
    wire N__32811;
    wire N__32810;
    wire N__32809;
    wire N__32806;
    wire N__32801;
    wire N__32800;
    wire N__32799;
    wire N__32798;
    wire N__32797;
    wire N__32796;
    wire N__32793;
    wire N__32792;
    wire N__32791;
    wire N__32790;
    wire N__32789;
    wire N__32788;
    wire N__32787;
    wire N__32784;
    wire N__32781;
    wire N__32778;
    wire N__32775;
    wire N__32772;
    wire N__32771;
    wire N__32768;
    wire N__32765;
    wire N__32764;
    wire N__32763;
    wire N__32762;
    wire N__32761;
    wire N__32760;
    wire N__32759;
    wire N__32758;
    wire N__32757;
    wire N__32756;
    wire N__32755;
    wire N__32754;
    wire N__32753;
    wire N__32752;
    wire N__32751;
    wire N__32750;
    wire N__32749;
    wire N__32748;
    wire N__32747;
    wire N__32746;
    wire N__32745;
    wire N__32744;
    wire N__32743;
    wire N__32738;
    wire N__32729;
    wire N__32724;
    wire N__32723;
    wire N__32722;
    wire N__32721;
    wire N__32720;
    wire N__32719;
    wire N__32718;
    wire N__32717;
    wire N__32716;
    wire N__32715;
    wire N__32712;
    wire N__32709;
    wire N__32706;
    wire N__32699;
    wire N__32696;
    wire N__32691;
    wire N__32682;
    wire N__32679;
    wire N__32678;
    wire N__32675;
    wire N__32672;
    wire N__32661;
    wire N__32656;
    wire N__32653;
    wire N__32652;
    wire N__32651;
    wire N__32650;
    wire N__32649;
    wire N__32648;
    wire N__32647;
    wire N__32644;
    wire N__32643;
    wire N__32640;
    wire N__32639;
    wire N__32638;
    wire N__32637;
    wire N__32636;
    wire N__32635;
    wire N__32634;
    wire N__32633;
    wire N__32632;
    wire N__32631;
    wire N__32630;
    wire N__32629;
    wire N__32628;
    wire N__32627;
    wire N__32626;
    wire N__32625;
    wire N__32624;
    wire N__32623;
    wire N__32622;
    wire N__32621;
    wire N__32620;
    wire N__32619;
    wire N__32618;
    wire N__32617;
    wire N__32616;
    wire N__32615;
    wire N__32614;
    wire N__32613;
    wire N__32612;
    wire N__32611;
    wire N__32610;
    wire N__32609;
    wire N__32608;
    wire N__32607;
    wire N__32606;
    wire N__32605;
    wire N__32604;
    wire N__32603;
    wire N__32602;
    wire N__32601;
    wire N__32600;
    wire N__32599;
    wire N__32598;
    wire N__32595;
    wire N__32588;
    wire N__32581;
    wire N__32566;
    wire N__32549;
    wire N__32542;
    wire N__32539;
    wire N__32536;
    wire N__32533;
    wire N__32526;
    wire N__32513;
    wire N__32508;
    wire N__32497;
    wire N__32494;
    wire N__32491;
    wire N__32488;
    wire N__32485;
    wire N__32478;
    wire N__32475;
    wire N__32464;
    wire N__32461;
    wire N__32458;
    wire N__32455;
    wire N__32438;
    wire N__32421;
    wire N__32404;
    wire N__32387;
    wire N__32372;
    wire N__32365;
    wire N__32360;
    wire N__32345;
    wire N__32334;
    wire N__32329;
    wire N__32324;
    wire N__32317;
    wire N__32312;
    wire N__32285;
    wire N__32282;
    wire N__32279;
    wire N__32278;
    wire N__32275;
    wire N__32272;
    wire N__32269;
    wire N__32264;
    wire N__32263;
    wire N__32260;
    wire N__32257;
    wire N__32256;
    wire N__32253;
    wire N__32250;
    wire N__32247;
    wire N__32246;
    wire N__32241;
    wire N__32238;
    wire N__32235;
    wire N__32232;
    wire N__32229;
    wire N__32226;
    wire N__32223;
    wire N__32216;
    wire N__32215;
    wire N__32214;
    wire N__32213;
    wire N__32208;
    wire N__32205;
    wire N__32202;
    wire N__32199;
    wire N__32196;
    wire N__32193;
    wire N__32190;
    wire N__32187;
    wire N__32184;
    wire N__32181;
    wire N__32178;
    wire N__32175;
    wire N__32172;
    wire N__32165;
    wire N__32162;
    wire N__32161;
    wire N__32158;
    wire N__32155;
    wire N__32152;
    wire N__32149;
    wire N__32144;
    wire N__32141;
    wire N__32140;
    wire N__32137;
    wire N__32134;
    wire N__32131;
    wire N__32126;
    wire N__32123;
    wire N__32120;
    wire N__32117;
    wire N__32114;
    wire N__32111;
    wire N__32110;
    wire N__32107;
    wire N__32106;
    wire N__32103;
    wire N__32100;
    wire N__32097;
    wire N__32094;
    wire N__32089;
    wire N__32084;
    wire N__32081;
    wire N__32078;
    wire N__32075;
    wire N__32072;
    wire N__32069;
    wire N__32066;
    wire N__32065;
    wire N__32064;
    wire N__32061;
    wire N__32058;
    wire N__32057;
    wire N__32054;
    wire N__32049;
    wire N__32046;
    wire N__32045;
    wire N__32042;
    wire N__32039;
    wire N__32036;
    wire N__32033;
    wire N__32026;
    wire N__32023;
    wire N__32020;
    wire N__32017;
    wire N__32014;
    wire N__32009;
    wire N__32006;
    wire N__32003;
    wire N__32000;
    wire N__31997;
    wire N__31996;
    wire N__31995;
    wire N__31994;
    wire N__31993;
    wire N__31992;
    wire N__31989;
    wire N__31988;
    wire N__31985;
    wire N__31982;
    wire N__31981;
    wire N__31980;
    wire N__31979;
    wire N__31978;
    wire N__31977;
    wire N__31976;
    wire N__31975;
    wire N__31974;
    wire N__31973;
    wire N__31972;
    wire N__31971;
    wire N__31970;
    wire N__31969;
    wire N__31968;
    wire N__31959;
    wire N__31952;
    wire N__31951;
    wire N__31950;
    wire N__31947;
    wire N__31944;
    wire N__31943;
    wire N__31942;
    wire N__31941;
    wire N__31938;
    wire N__31937;
    wire N__31934;
    wire N__31929;
    wire N__31928;
    wire N__31927;
    wire N__31926;
    wire N__31925;
    wire N__31924;
    wire N__31923;
    wire N__31922;
    wire N__31921;
    wire N__31920;
    wire N__31919;
    wire N__31918;
    wire N__31917;
    wire N__31914;
    wire N__31911;
    wire N__31908;
    wire N__31907;
    wire N__31906;
    wire N__31903;
    wire N__31894;
    wire N__31893;
    wire N__31892;
    wire N__31887;
    wire N__31878;
    wire N__31877;
    wire N__31876;
    wire N__31875;
    wire N__31872;
    wire N__31871;
    wire N__31870;
    wire N__31867;
    wire N__31864;
    wire N__31861;
    wire N__31856;
    wire N__31853;
    wire N__31852;
    wire N__31851;
    wire N__31850;
    wire N__31849;
    wire N__31848;
    wire N__31847;
    wire N__31844;
    wire N__31841;
    wire N__31840;
    wire N__31839;
    wire N__31838;
    wire N__31835;
    wire N__31832;
    wire N__31831;
    wire N__31830;
    wire N__31829;
    wire N__31828;
    wire N__31825;
    wire N__31824;
    wire N__31823;
    wire N__31822;
    wire N__31821;
    wire N__31820;
    wire N__31819;
    wire N__31818;
    wire N__31817;
    wire N__31816;
    wire N__31813;
    wire N__31810;
    wire N__31809;
    wire N__31808;
    wire N__31807;
    wire N__31806;
    wire N__31805;
    wire N__31804;
    wire N__31803;
    wire N__31800;
    wire N__31799;
    wire N__31798;
    wire N__31797;
    wire N__31796;
    wire N__31795;
    wire N__31792;
    wire N__31791;
    wire N__31790;
    wire N__31789;
    wire N__31786;
    wire N__31783;
    wire N__31780;
    wire N__31777;
    wire N__31774;
    wire N__31771;
    wire N__31768;
    wire N__31765;
    wire N__31760;
    wire N__31755;
    wire N__31750;
    wire N__31747;
    wire N__31740;
    wire N__31731;
    wire N__31724;
    wire N__31723;
    wire N__31720;
    wire N__31717;
    wire N__31714;
    wire N__31713;
    wire N__31712;
    wire N__31701;
    wire N__31686;
    wire N__31675;
    wire N__31664;
    wire N__31655;
    wire N__31642;
    wire N__31631;
    wire N__31618;
    wire N__31615;
    wire N__31604;
    wire N__31597;
    wire N__31592;
    wire N__31583;
    wire N__31570;
    wire N__31541;
    wire N__31538;
    wire N__31537;
    wire N__31534;
    wire N__31531;
    wire N__31528;
    wire N__31525;
    wire N__31520;
    wire N__31517;
    wire N__31516;
    wire N__31513;
    wire N__31512;
    wire N__31509;
    wire N__31506;
    wire N__31505;
    wire N__31502;
    wire N__31499;
    wire N__31496;
    wire N__31493;
    wire N__31486;
    wire N__31483;
    wire N__31478;
    wire N__31475;
    wire N__31472;
    wire N__31469;
    wire N__31466;
    wire N__31463;
    wire N__31462;
    wire N__31459;
    wire N__31456;
    wire N__31451;
    wire N__31450;
    wire N__31447;
    wire N__31444;
    wire N__31439;
    wire N__31436;
    wire N__31433;
    wire N__31430;
    wire N__31429;
    wire N__31426;
    wire N__31423;
    wire N__31418;
    wire N__31415;
    wire N__31414;
    wire N__31411;
    wire N__31410;
    wire N__31409;
    wire N__31406;
    wire N__31403;
    wire N__31400;
    wire N__31397;
    wire N__31392;
    wire N__31389;
    wire N__31382;
    wire N__31379;
    wire N__31378;
    wire N__31377;
    wire N__31376;
    wire N__31373;
    wire N__31370;
    wire N__31367;
    wire N__31364;
    wire N__31363;
    wire N__31358;
    wire N__31355;
    wire N__31352;
    wire N__31349;
    wire N__31346;
    wire N__31341;
    wire N__31334;
    wire N__31333;
    wire N__31328;
    wire N__31325;
    wire N__31324;
    wire N__31319;
    wire N__31316;
    wire N__31313;
    wire N__31310;
    wire N__31309;
    wire N__31306;
    wire N__31303;
    wire N__31298;
    wire N__31295;
    wire N__31292;
    wire N__31291;
    wire N__31288;
    wire N__31287;
    wire N__31284;
    wire N__31281;
    wire N__31276;
    wire N__31271;
    wire N__31270;
    wire N__31267;
    wire N__31264;
    wire N__31263;
    wire N__31260;
    wire N__31257;
    wire N__31254;
    wire N__31251;
    wire N__31248;
    wire N__31247;
    wire N__31244;
    wire N__31239;
    wire N__31236;
    wire N__31233;
    wire N__31226;
    wire N__31223;
    wire N__31220;
    wire N__31219;
    wire N__31216;
    wire N__31213;
    wire N__31210;
    wire N__31205;
    wire N__31204;
    wire N__31201;
    wire N__31198;
    wire N__31195;
    wire N__31190;
    wire N__31187;
    wire N__31184;
    wire N__31181;
    wire N__31178;
    wire N__31175;
    wire N__31172;
    wire N__31171;
    wire N__31168;
    wire N__31165;
    wire N__31162;
    wire N__31157;
    wire N__31156;
    wire N__31155;
    wire N__31154;
    wire N__31147;
    wire N__31144;
    wire N__31143;
    wire N__31142;
    wire N__31141;
    wire N__31140;
    wire N__31135;
    wire N__31134;
    wire N__31133;
    wire N__31132;
    wire N__31131;
    wire N__31130;
    wire N__31129;
    wire N__31128;
    wire N__31125;
    wire N__31124;
    wire N__31123;
    wire N__31122;
    wire N__31119;
    wire N__31118;
    wire N__31113;
    wire N__31110;
    wire N__31101;
    wire N__31100;
    wire N__31097;
    wire N__31096;
    wire N__31095;
    wire N__31094;
    wire N__31091;
    wire N__31088;
    wire N__31085;
    wire N__31084;
    wire N__31081;
    wire N__31078;
    wire N__31077;
    wire N__31076;
    wire N__31075;
    wire N__31074;
    wire N__31073;
    wire N__31066;
    wire N__31059;
    wire N__31054;
    wire N__31053;
    wire N__31052;
    wire N__31049;
    wire N__31044;
    wire N__31043;
    wire N__31036;
    wire N__31035;
    wire N__31034;
    wire N__31033;
    wire N__31032;
    wire N__31031;
    wire N__31030;
    wire N__31027;
    wire N__31024;
    wire N__31021;
    wire N__31016;
    wire N__31009;
    wire N__31002;
    wire N__30995;
    wire N__30992;
    wire N__30991;
    wire N__30990;
    wire N__30989;
    wire N__30988;
    wire N__30987;
    wire N__30986;
    wire N__30985;
    wire N__30984;
    wire N__30983;
    wire N__30982;
    wire N__30981;
    wire N__30980;
    wire N__30979;
    wire N__30978;
    wire N__30975;
    wire N__30972;
    wire N__30969;
    wire N__30968;
    wire N__30967;
    wire N__30966;
    wire N__30965;
    wire N__30964;
    wire N__30963;
    wire N__30962;
    wire N__30957;
    wire N__30954;
    wire N__30951;
    wire N__30948;
    wire N__30945;
    wire N__30942;
    wire N__30931;
    wire N__30930;
    wire N__30927;
    wire N__30924;
    wire N__30921;
    wire N__30916;
    wire N__30911;
    wire N__30908;
    wire N__30899;
    wire N__30892;
    wire N__30885;
    wire N__30876;
    wire N__30875;
    wire N__30874;
    wire N__30871;
    wire N__30866;
    wire N__30861;
    wire N__30854;
    wire N__30849;
    wire N__30846;
    wire N__30841;
    wire N__30824;
    wire N__30817;
    wire N__30808;
    wire N__30797;
    wire N__30796;
    wire N__30795;
    wire N__30794;
    wire N__30793;
    wire N__30792;
    wire N__30791;
    wire N__30790;
    wire N__30789;
    wire N__30782;
    wire N__30777;
    wire N__30774;
    wire N__30773;
    wire N__30772;
    wire N__30771;
    wire N__30770;
    wire N__30769;
    wire N__30768;
    wire N__30767;
    wire N__30766;
    wire N__30765;
    wire N__30764;
    wire N__30763;
    wire N__30762;
    wire N__30761;
    wire N__30760;
    wire N__30759;
    wire N__30758;
    wire N__30755;
    wire N__30754;
    wire N__30753;
    wire N__30750;
    wire N__30747;
    wire N__30740;
    wire N__30739;
    wire N__30738;
    wire N__30737;
    wire N__30736;
    wire N__30735;
    wire N__30734;
    wire N__30733;
    wire N__30726;
    wire N__30723;
    wire N__30722;
    wire N__30719;
    wire N__30714;
    wire N__30699;
    wire N__30696;
    wire N__30695;
    wire N__30694;
    wire N__30691;
    wire N__30688;
    wire N__30685;
    wire N__30682;
    wire N__30675;
    wire N__30674;
    wire N__30673;
    wire N__30672;
    wire N__30671;
    wire N__30670;
    wire N__30669;
    wire N__30664;
    wire N__30655;
    wire N__30652;
    wire N__30649;
    wire N__30646;
    wire N__30645;
    wire N__30644;
    wire N__30643;
    wire N__30640;
    wire N__30631;
    wire N__30626;
    wire N__30625;
    wire N__30622;
    wire N__30617;
    wire N__30612;
    wire N__30609;
    wire N__30604;
    wire N__30601;
    wire N__30598;
    wire N__30595;
    wire N__30590;
    wire N__30585;
    wire N__30582;
    wire N__30575;
    wire N__30568;
    wire N__30565;
    wire N__30564;
    wire N__30563;
    wire N__30562;
    wire N__30561;
    wire N__30560;
    wire N__30555;
    wire N__30550;
    wire N__30537;
    wire N__30532;
    wire N__30529;
    wire N__30526;
    wire N__30523;
    wire N__30514;
    wire N__30509;
    wire N__30504;
    wire N__30501;
    wire N__30488;
    wire N__30485;
    wire N__30482;
    wire N__30479;
    wire N__30476;
    wire N__30473;
    wire N__30472;
    wire N__30469;
    wire N__30466;
    wire N__30463;
    wire N__30462;
    wire N__30457;
    wire N__30454;
    wire N__30451;
    wire N__30446;
    wire N__30445;
    wire N__30440;
    wire N__30437;
    wire N__30436;
    wire N__30431;
    wire N__30428;
    wire N__30427;
    wire N__30422;
    wire N__30419;
    wire N__30418;
    wire N__30413;
    wire N__30410;
    wire N__30407;
    wire N__30406;
    wire N__30403;
    wire N__30400;
    wire N__30395;
    wire N__30394;
    wire N__30389;
    wire N__30386;
    wire N__30383;
    wire N__30380;
    wire N__30377;
    wire N__30376;
    wire N__30375;
    wire N__30374;
    wire N__30373;
    wire N__30372;
    wire N__30367;
    wire N__30364;
    wire N__30359;
    wire N__30356;
    wire N__30347;
    wire N__30344;
    wire N__30341;
    wire N__30338;
    wire N__30335;
    wire N__30334;
    wire N__30333;
    wire N__30330;
    wire N__30327;
    wire N__30324;
    wire N__30317;
    wire N__30316;
    wire N__30315;
    wire N__30314;
    wire N__30311;
    wire N__30310;
    wire N__30309;
    wire N__30306;
    wire N__30295;
    wire N__30294;
    wire N__30293;
    wire N__30288;
    wire N__30283;
    wire N__30278;
    wire N__30275;
    wire N__30272;
    wire N__30269;
    wire N__30266;
    wire N__30263;
    wire N__30260;
    wire N__30257;
    wire N__30254;
    wire N__30251;
    wire N__30250;
    wire N__30247;
    wire N__30244;
    wire N__30239;
    wire N__30236;
    wire N__30235;
    wire N__30232;
    wire N__30229;
    wire N__30226;
    wire N__30221;
    wire N__30218;
    wire N__30215;
    wire N__30214;
    wire N__30211;
    wire N__30208;
    wire N__30205;
    wire N__30200;
    wire N__30197;
    wire N__30194;
    wire N__30191;
    wire N__30188;
    wire N__30185;
    wire N__30182;
    wire N__30179;
    wire N__30176;
    wire N__30173;
    wire N__30170;
    wire N__30167;
    wire N__30164;
    wire N__30161;
    wire N__30158;
    wire N__30157;
    wire N__30152;
    wire N__30149;
    wire N__30148;
    wire N__30143;
    wire N__30140;
    wire N__30139;
    wire N__30138;
    wire N__30133;
    wire N__30130;
    wire N__30125;
    wire N__30122;
    wire N__30119;
    wire N__30118;
    wire N__30113;
    wire N__30110;
    wire N__30109;
    wire N__30108;
    wire N__30107;
    wire N__30104;
    wire N__30101;
    wire N__30096;
    wire N__30089;
    wire N__30086;
    wire N__30085;
    wire N__30084;
    wire N__30077;
    wire N__30074;
    wire N__30071;
    wire N__30070;
    wire N__30069;
    wire N__30068;
    wire N__30065;
    wire N__30062;
    wire N__30059;
    wire N__30056;
    wire N__30047;
    wire N__30044;
    wire N__30041;
    wire N__30040;
    wire N__30037;
    wire N__30034;
    wire N__30031;
    wire N__30026;
    wire N__30025;
    wire N__30020;
    wire N__30017;
    wire N__30014;
    wire N__30013;
    wire N__30010;
    wire N__30007;
    wire N__30002;
    wire N__29999;
    wire N__29996;
    wire N__29993;
    wire N__29992;
    wire N__29989;
    wire N__29988;
    wire N__29985;
    wire N__29982;
    wire N__29979;
    wire N__29976;
    wire N__29969;
    wire N__29966;
    wire N__29965;
    wire N__29962;
    wire N__29959;
    wire N__29958;
    wire N__29955;
    wire N__29952;
    wire N__29949;
    wire N__29942;
    wire N__29939;
    wire N__29938;
    wire N__29935;
    wire N__29932;
    wire N__29927;
    wire N__29926;
    wire N__29923;
    wire N__29920;
    wire N__29919;
    wire N__29916;
    wire N__29913;
    wire N__29910;
    wire N__29907;
    wire N__29904;
    wire N__29897;
    wire N__29896;
    wire N__29893;
    wire N__29890;
    wire N__29887;
    wire N__29882;
    wire N__29881;
    wire N__29878;
    wire N__29875;
    wire N__29870;
    wire N__29869;
    wire N__29866;
    wire N__29863;
    wire N__29858;
    wire N__29855;
    wire N__29852;
    wire N__29851;
    wire N__29848;
    wire N__29845;
    wire N__29844;
    wire N__29841;
    wire N__29838;
    wire N__29835;
    wire N__29828;
    wire N__29827;
    wire N__29826;
    wire N__29823;
    wire N__29820;
    wire N__29817;
    wire N__29814;
    wire N__29807;
    wire N__29804;
    wire N__29801;
    wire N__29800;
    wire N__29797;
    wire N__29794;
    wire N__29791;
    wire N__29788;
    wire N__29785;
    wire N__29784;
    wire N__29781;
    wire N__29778;
    wire N__29775;
    wire N__29772;
    wire N__29769;
    wire N__29762;
    wire N__29759;
    wire N__29756;
    wire N__29753;
    wire N__29750;
    wire N__29747;
    wire N__29744;
    wire N__29741;
    wire N__29738;
    wire N__29735;
    wire N__29734;
    wire N__29733;
    wire N__29730;
    wire N__29727;
    wire N__29724;
    wire N__29717;
    wire N__29714;
    wire N__29713;
    wire N__29712;
    wire N__29705;
    wire N__29702;
    wire N__29701;
    wire N__29700;
    wire N__29699;
    wire N__29696;
    wire N__29689;
    wire N__29684;
    wire N__29681;
    wire N__29678;
    wire N__29677;
    wire N__29676;
    wire N__29673;
    wire N__29668;
    wire N__29665;
    wire N__29660;
    wire N__29659;
    wire N__29658;
    wire N__29655;
    wire N__29652;
    wire N__29649;
    wire N__29642;
    wire N__29641;
    wire N__29640;
    wire N__29637;
    wire N__29634;
    wire N__29631;
    wire N__29628;
    wire N__29621;
    wire N__29620;
    wire N__29619;
    wire N__29616;
    wire N__29613;
    wire N__29610;
    wire N__29603;
    wire N__29602;
    wire N__29601;
    wire N__29598;
    wire N__29595;
    wire N__29592;
    wire N__29585;
    wire N__29582;
    wire N__29579;
    wire N__29578;
    wire N__29577;
    wire N__29574;
    wire N__29569;
    wire N__29564;
    wire N__29563;
    wire N__29558;
    wire N__29557;
    wire N__29554;
    wire N__29553;
    wire N__29550;
    wire N__29547;
    wire N__29544;
    wire N__29541;
    wire N__29538;
    wire N__29531;
    wire N__29530;
    wire N__29527;
    wire N__29524;
    wire N__29523;
    wire N__29518;
    wire N__29515;
    wire N__29512;
    wire N__29507;
    wire N__29506;
    wire N__29503;
    wire N__29500;
    wire N__29497;
    wire N__29494;
    wire N__29491;
    wire N__29488;
    wire N__29485;
    wire N__29480;
    wire N__29479;
    wire N__29476;
    wire N__29473;
    wire N__29470;
    wire N__29467;
    wire N__29464;
    wire N__29461;
    wire N__29458;
    wire N__29453;
    wire N__29450;
    wire N__29447;
    wire N__29446;
    wire N__29443;
    wire N__29440;
    wire N__29437;
    wire N__29434;
    wire N__29429;
    wire N__29426;
    wire N__29423;
    wire N__29420;
    wire N__29419;
    wire N__29416;
    wire N__29413;
    wire N__29412;
    wire N__29409;
    wire N__29406;
    wire N__29403;
    wire N__29400;
    wire N__29393;
    wire N__29392;
    wire N__29391;
    wire N__29390;
    wire N__29389;
    wire N__29388;
    wire N__29385;
    wire N__29382;
    wire N__29375;
    wire N__29372;
    wire N__29365;
    wire N__29362;
    wire N__29357;
    wire N__29354;
    wire N__29351;
    wire N__29348;
    wire N__29345;
    wire N__29344;
    wire N__29341;
    wire N__29338;
    wire N__29333;
    wire N__29330;
    wire N__29327;
    wire N__29324;
    wire N__29323;
    wire N__29320;
    wire N__29317;
    wire N__29312;
    wire N__29309;
    wire N__29306;
    wire N__29303;
    wire N__29300;
    wire N__29297;
    wire N__29294;
    wire N__29291;
    wire N__29288;
    wire N__29285;
    wire N__29282;
    wire N__29279;
    wire N__29276;
    wire N__29273;
    wire N__29270;
    wire N__29269;
    wire N__29266;
    wire N__29263;
    wire N__29258;
    wire N__29257;
    wire N__29254;
    wire N__29251;
    wire N__29248;
    wire N__29247;
    wire N__29246;
    wire N__29245;
    wire N__29240;
    wire N__29235;
    wire N__29232;
    wire N__29229;
    wire N__29226;
    wire N__29223;
    wire N__29220;
    wire N__29215;
    wire N__29210;
    wire N__29207;
    wire N__29204;
    wire N__29201;
    wire N__29198;
    wire N__29197;
    wire N__29194;
    wire N__29191;
    wire N__29188;
    wire N__29185;
    wire N__29180;
    wire N__29177;
    wire N__29174;
    wire N__29173;
    wire N__29170;
    wire N__29167;
    wire N__29162;
    wire N__29159;
    wire N__29156;
    wire N__29153;
    wire N__29150;
    wire N__29147;
    wire N__29144;
    wire N__29141;
    wire N__29138;
    wire N__29135;
    wire N__29134;
    wire N__29133;
    wire N__29130;
    wire N__29127;
    wire N__29126;
    wire N__29123;
    wire N__29122;
    wire N__29119;
    wire N__29116;
    wire N__29113;
    wire N__29110;
    wire N__29107;
    wire N__29102;
    wire N__29093;
    wire N__29090;
    wire N__29089;
    wire N__29088;
    wire N__29085;
    wire N__29084;
    wire N__29081;
    wire N__29078;
    wire N__29075;
    wire N__29072;
    wire N__29069;
    wire N__29060;
    wire N__29057;
    wire N__29056;
    wire N__29053;
    wire N__29050;
    wire N__29047;
    wire N__29044;
    wire N__29041;
    wire N__29040;
    wire N__29035;
    wire N__29032;
    wire N__29031;
    wire N__29030;
    wire N__29027;
    wire N__29022;
    wire N__29019;
    wire N__29012;
    wire N__29011;
    wire N__29010;
    wire N__29007;
    wire N__29002;
    wire N__29001;
    wire N__28998;
    wire N__28995;
    wire N__28992;
    wire N__28989;
    wire N__28986;
    wire N__28979;
    wire N__28978;
    wire N__28975;
    wire N__28974;
    wire N__28971;
    wire N__28968;
    wire N__28965;
    wire N__28962;
    wire N__28959;
    wire N__28956;
    wire N__28953;
    wire N__28950;
    wire N__28947;
    wire N__28942;
    wire N__28937;
    wire N__28934;
    wire N__28933;
    wire N__28930;
    wire N__28927;
    wire N__28924;
    wire N__28921;
    wire N__28920;
    wire N__28917;
    wire N__28914;
    wire N__28911;
    wire N__28908;
    wire N__28905;
    wire N__28902;
    wire N__28895;
    wire N__28894;
    wire N__28891;
    wire N__28888;
    wire N__28885;
    wire N__28880;
    wire N__28877;
    wire N__28874;
    wire N__28873;
    wire N__28870;
    wire N__28867;
    wire N__28864;
    wire N__28861;
    wire N__28856;
    wire N__28853;
    wire N__28850;
    wire N__28849;
    wire N__28846;
    wire N__28843;
    wire N__28840;
    wire N__28837;
    wire N__28832;
    wire N__28829;
    wire N__28826;
    wire N__28823;
    wire N__28820;
    wire N__28819;
    wire N__28816;
    wire N__28813;
    wire N__28808;
    wire N__28807;
    wire N__28804;
    wire N__28801;
    wire N__28798;
    wire N__28795;
    wire N__28790;
    wire N__28787;
    wire N__28784;
    wire N__28781;
    wire N__28778;
    wire N__28775;
    wire N__28774;
    wire N__28773;
    wire N__28768;
    wire N__28767;
    wire N__28764;
    wire N__28761;
    wire N__28760;
    wire N__28759;
    wire N__28756;
    wire N__28753;
    wire N__28750;
    wire N__28745;
    wire N__28740;
    wire N__28733;
    wire N__28732;
    wire N__28727;
    wire N__28724;
    wire N__28723;
    wire N__28720;
    wire N__28717;
    wire N__28716;
    wire N__28715;
    wire N__28714;
    wire N__28711;
    wire N__28706;
    wire N__28701;
    wire N__28694;
    wire N__28693;
    wire N__28692;
    wire N__28689;
    wire N__28686;
    wire N__28683;
    wire N__28680;
    wire N__28679;
    wire N__28672;
    wire N__28669;
    wire N__28664;
    wire N__28661;
    wire N__28658;
    wire N__28655;
    wire N__28652;
    wire N__28649;
    wire N__28646;
    wire N__28645;
    wire N__28642;
    wire N__28641;
    wire N__28638;
    wire N__28635;
    wire N__28632;
    wire N__28631;
    wire N__28628;
    wire N__28625;
    wire N__28622;
    wire N__28621;
    wire N__28618;
    wire N__28615;
    wire N__28610;
    wire N__28607;
    wire N__28604;
    wire N__28595;
    wire N__28592;
    wire N__28591;
    wire N__28588;
    wire N__28585;
    wire N__28582;
    wire N__28579;
    wire N__28576;
    wire N__28573;
    wire N__28568;
    wire N__28565;
    wire N__28564;
    wire N__28563;
    wire N__28560;
    wire N__28557;
    wire N__28554;
    wire N__28551;
    wire N__28546;
    wire N__28541;
    wire N__28538;
    wire N__28535;
    wire N__28534;
    wire N__28531;
    wire N__28530;
    wire N__28527;
    wire N__28524;
    wire N__28521;
    wire N__28518;
    wire N__28513;
    wire N__28510;
    wire N__28507;
    wire N__28502;
    wire N__28499;
    wire N__28496;
    wire N__28493;
    wire N__28492;
    wire N__28491;
    wire N__28488;
    wire N__28485;
    wire N__28482;
    wire N__28481;
    wire N__28478;
    wire N__28477;
    wire N__28476;
    wire N__28473;
    wire N__28470;
    wire N__28467;
    wire N__28464;
    wire N__28459;
    wire N__28454;
    wire N__28451;
    wire N__28446;
    wire N__28439;
    wire N__28438;
    wire N__28435;
    wire N__28434;
    wire N__28433;
    wire N__28432;
    wire N__28429;
    wire N__28426;
    wire N__28423;
    wire N__28420;
    wire N__28417;
    wire N__28412;
    wire N__28409;
    wire N__28404;
    wire N__28397;
    wire N__28394;
    wire N__28391;
    wire N__28388;
    wire N__28385;
    wire N__28384;
    wire N__28381;
    wire N__28378;
    wire N__28375;
    wire N__28372;
    wire N__28369;
    wire N__28366;
    wire N__28365;
    wire N__28362;
    wire N__28359;
    wire N__28356;
    wire N__28353;
    wire N__28350;
    wire N__28343;
    wire N__28342;
    wire N__28341;
    wire N__28340;
    wire N__28339;
    wire N__28336;
    wire N__28335;
    wire N__28332;
    wire N__28329;
    wire N__28326;
    wire N__28323;
    wire N__28320;
    wire N__28317;
    wire N__28316;
    wire N__28315;
    wire N__28312;
    wire N__28305;
    wire N__28300;
    wire N__28297;
    wire N__28294;
    wire N__28291;
    wire N__28286;
    wire N__28283;
    wire N__28274;
    wire N__28271;
    wire N__28268;
    wire N__28265;
    wire N__28262;
    wire N__28261;
    wire N__28258;
    wire N__28255;
    wire N__28254;
    wire N__28251;
    wire N__28248;
    wire N__28245;
    wire N__28242;
    wire N__28239;
    wire N__28236;
    wire N__28233;
    wire N__28230;
    wire N__28227;
    wire N__28220;
    wire N__28217;
    wire N__28216;
    wire N__28213;
    wire N__28210;
    wire N__28207;
    wire N__28204;
    wire N__28199;
    wire N__28196;
    wire N__28193;
    wire N__28190;
    wire N__28187;
    wire N__28184;
    wire N__28183;
    wire N__28182;
    wire N__28181;
    wire N__28178;
    wire N__28175;
    wire N__28174;
    wire N__28171;
    wire N__28168;
    wire N__28165;
    wire N__28162;
    wire N__28159;
    wire N__28148;
    wire N__28145;
    wire N__28144;
    wire N__28143;
    wire N__28142;
    wire N__28141;
    wire N__28138;
    wire N__28131;
    wire N__28128;
    wire N__28125;
    wire N__28118;
    wire N__28117;
    wire N__28114;
    wire N__28111;
    wire N__28108;
    wire N__28105;
    wire N__28100;
    wire N__28099;
    wire N__28098;
    wire N__28095;
    wire N__28094;
    wire N__28089;
    wire N__28086;
    wire N__28083;
    wire N__28080;
    wire N__28077;
    wire N__28072;
    wire N__28067;
    wire N__28066;
    wire N__28063;
    wire N__28062;
    wire N__28059;
    wire N__28058;
    wire N__28053;
    wire N__28052;
    wire N__28049;
    wire N__28046;
    wire N__28045;
    wire N__28044;
    wire N__28043;
    wire N__28042;
    wire N__28039;
    wire N__28036;
    wire N__28035;
    wire N__28034;
    wire N__28033;
    wire N__28028;
    wire N__28025;
    wire N__28024;
    wire N__28023;
    wire N__28016;
    wire N__28013;
    wire N__28010;
    wire N__28009;
    wire N__28008;
    wire N__28007;
    wire N__28006;
    wire N__28005;
    wire N__28004;
    wire N__28001;
    wire N__27998;
    wire N__27995;
    wire N__27990;
    wire N__27985;
    wire N__27978;
    wire N__27971;
    wire N__27964;
    wire N__27947;
    wire N__27946;
    wire N__27943;
    wire N__27942;
    wire N__27939;
    wire N__27936;
    wire N__27933;
    wire N__27930;
    wire N__27925;
    wire N__27922;
    wire N__27917;
    wire N__27914;
    wire N__27911;
    wire N__27908;
    wire N__27905;
    wire N__27904;
    wire N__27901;
    wire N__27898;
    wire N__27897;
    wire N__27896;
    wire N__27895;
    wire N__27890;
    wire N__27885;
    wire N__27882;
    wire N__27877;
    wire N__27872;
    wire N__27869;
    wire N__27866;
    wire N__27865;
    wire N__27862;
    wire N__27859;
    wire N__27856;
    wire N__27851;
    wire N__27850;
    wire N__27847;
    wire N__27844;
    wire N__27839;
    wire N__27836;
    wire N__27835;
    wire N__27832;
    wire N__27831;
    wire N__27828;
    wire N__27825;
    wire N__27824;
    wire N__27823;
    wire N__27820;
    wire N__27817;
    wire N__27814;
    wire N__27811;
    wire N__27808;
    wire N__27797;
    wire N__27796;
    wire N__27793;
    wire N__27790;
    wire N__27789;
    wire N__27786;
    wire N__27783;
    wire N__27782;
    wire N__27779;
    wire N__27778;
    wire N__27773;
    wire N__27770;
    wire N__27767;
    wire N__27764;
    wire N__27761;
    wire N__27756;
    wire N__27749;
    wire N__27746;
    wire N__27743;
    wire N__27742;
    wire N__27741;
    wire N__27740;
    wire N__27737;
    wire N__27734;
    wire N__27731;
    wire N__27728;
    wire N__27719;
    wire N__27718;
    wire N__27715;
    wire N__27714;
    wire N__27711;
    wire N__27708;
    wire N__27707;
    wire N__27704;
    wire N__27699;
    wire N__27696;
    wire N__27689;
    wire N__27686;
    wire N__27683;
    wire N__27682;
    wire N__27681;
    wire N__27680;
    wire N__27677;
    wire N__27672;
    wire N__27669;
    wire N__27662;
    wire N__27659;
    wire N__27658;
    wire N__27657;
    wire N__27654;
    wire N__27649;
    wire N__27644;
    wire N__27643;
    wire N__27640;
    wire N__27637;
    wire N__27634;
    wire N__27631;
    wire N__27630;
    wire N__27629;
    wire N__27626;
    wire N__27623;
    wire N__27618;
    wire N__27611;
    wire N__27608;
    wire N__27605;
    wire N__27604;
    wire N__27601;
    wire N__27598;
    wire N__27597;
    wire N__27596;
    wire N__27593;
    wire N__27590;
    wire N__27585;
    wire N__27578;
    wire N__27575;
    wire N__27572;
    wire N__27571;
    wire N__27568;
    wire N__27565;
    wire N__27564;
    wire N__27561;
    wire N__27558;
    wire N__27555;
    wire N__27548;
    wire N__27545;
    wire N__27542;
    wire N__27539;
    wire N__27538;
    wire N__27537;
    wire N__27536;
    wire N__27533;
    wire N__27528;
    wire N__27525;
    wire N__27518;
    wire N__27517;
    wire N__27516;
    wire N__27513;
    wire N__27510;
    wire N__27509;
    wire N__27506;
    wire N__27503;
    wire N__27500;
    wire N__27497;
    wire N__27494;
    wire N__27491;
    wire N__27486;
    wire N__27481;
    wire N__27478;
    wire N__27473;
    wire N__27470;
    wire N__27467;
    wire N__27466;
    wire N__27463;
    wire N__27460;
    wire N__27455;
    wire N__27454;
    wire N__27453;
    wire N__27450;
    wire N__27447;
    wire N__27442;
    wire N__27437;
    wire N__27434;
    wire N__27431;
    wire N__27428;
    wire N__27427;
    wire N__27426;
    wire N__27423;
    wire N__27420;
    wire N__27417;
    wire N__27414;
    wire N__27407;
    wire N__27404;
    wire N__27403;
    wire N__27400;
    wire N__27397;
    wire N__27394;
    wire N__27391;
    wire N__27390;
    wire N__27389;
    wire N__27384;
    wire N__27379;
    wire N__27376;
    wire N__27371;
    wire N__27368;
    wire N__27365;
    wire N__27364;
    wire N__27361;
    wire N__27358;
    wire N__27357;
    wire N__27354;
    wire N__27351;
    wire N__27348;
    wire N__27341;
    wire N__27338;
    wire N__27335;
    wire N__27332;
    wire N__27329;
    wire N__27326;
    wire N__27325;
    wire N__27322;
    wire N__27319;
    wire N__27316;
    wire N__27315;
    wire N__27314;
    wire N__27311;
    wire N__27308;
    wire N__27305;
    wire N__27302;
    wire N__27299;
    wire N__27296;
    wire N__27293;
    wire N__27284;
    wire N__27281;
    wire N__27280;
    wire N__27277;
    wire N__27276;
    wire N__27275;
    wire N__27272;
    wire N__27271;
    wire N__27268;
    wire N__27265;
    wire N__27262;
    wire N__27259;
    wire N__27256;
    wire N__27245;
    wire N__27242;
    wire N__27239;
    wire N__27236;
    wire N__27233;
    wire N__27232;
    wire N__27231;
    wire N__27228;
    wire N__27225;
    wire N__27222;
    wire N__27215;
    wire N__27212;
    wire N__27209;
    wire N__27206;
    wire N__27203;
    wire N__27200;
    wire N__27199;
    wire N__27198;
    wire N__27195;
    wire N__27192;
    wire N__27189;
    wire N__27182;
    wire N__27179;
    wire N__27176;
    wire N__27175;
    wire N__27174;
    wire N__27173;
    wire N__27172;
    wire N__27169;
    wire N__27166;
    wire N__27161;
    wire N__27158;
    wire N__27149;
    wire N__27146;
    wire N__27143;
    wire N__27140;
    wire N__27137;
    wire N__27134;
    wire N__27133;
    wire N__27130;
    wire N__27127;
    wire N__27122;
    wire N__27119;
    wire N__27116;
    wire N__27115;
    wire N__27112;
    wire N__27111;
    wire N__27108;
    wire N__27105;
    wire N__27104;
    wire N__27103;
    wire N__27100;
    wire N__27097;
    wire N__27094;
    wire N__27091;
    wire N__27088;
    wire N__27077;
    wire N__27074;
    wire N__27073;
    wire N__27070;
    wire N__27067;
    wire N__27064;
    wire N__27063;
    wire N__27062;
    wire N__27059;
    wire N__27056;
    wire N__27053;
    wire N__27050;
    wire N__27041;
    wire N__27038;
    wire N__27037;
    wire N__27034;
    wire N__27033;
    wire N__27032;
    wire N__27029;
    wire N__27026;
    wire N__27023;
    wire N__27022;
    wire N__27019;
    wire N__27016;
    wire N__27013;
    wire N__27010;
    wire N__27007;
    wire N__26996;
    wire N__26993;
    wire N__26990;
    wire N__26989;
    wire N__26986;
    wire N__26985;
    wire N__26982;
    wire N__26979;
    wire N__26978;
    wire N__26977;
    wire N__26974;
    wire N__26971;
    wire N__26968;
    wire N__26965;
    wire N__26962;
    wire N__26951;
    wire N__26948;
    wire N__26945;
    wire N__26942;
    wire N__26941;
    wire N__26938;
    wire N__26935;
    wire N__26934;
    wire N__26933;
    wire N__26930;
    wire N__26929;
    wire N__26926;
    wire N__26925;
    wire N__26922;
    wire N__26919;
    wire N__26916;
    wire N__26913;
    wire N__26910;
    wire N__26907;
    wire N__26906;
    wire N__26905;
    wire N__26902;
    wire N__26895;
    wire N__26890;
    wire N__26887;
    wire N__26884;
    wire N__26879;
    wire N__26870;
    wire N__26867;
    wire N__26864;
    wire N__26863;
    wire N__26860;
    wire N__26857;
    wire N__26854;
    wire N__26849;
    wire N__26846;
    wire N__26845;
    wire N__26844;
    wire N__26843;
    wire N__26842;
    wire N__26841;
    wire N__26840;
    wire N__26835;
    wire N__26834;
    wire N__26833;
    wire N__26828;
    wire N__26827;
    wire N__26826;
    wire N__26823;
    wire N__26818;
    wire N__26815;
    wire N__26812;
    wire N__26809;
    wire N__26806;
    wire N__26801;
    wire N__26800;
    wire N__26799;
    wire N__26798;
    wire N__26795;
    wire N__26786;
    wire N__26785;
    wire N__26784;
    wire N__26783;
    wire N__26782;
    wire N__26781;
    wire N__26780;
    wire N__26775;
    wire N__26768;
    wire N__26765;
    wire N__26762;
    wire N__26759;
    wire N__26758;
    wire N__26755;
    wire N__26750;
    wire N__26745;
    wire N__26742;
    wire N__26733;
    wire N__26730;
    wire N__26719;
    wire N__26714;
    wire N__26711;
    wire N__26710;
    wire N__26707;
    wire N__26704;
    wire N__26701;
    wire N__26696;
    wire N__26693;
    wire N__26690;
    wire N__26687;
    wire N__26684;
    wire N__26681;
    wire N__26678;
    wire N__26677;
    wire N__26676;
    wire N__26675;
    wire N__26674;
    wire N__26673;
    wire N__26672;
    wire N__26669;
    wire N__26668;
    wire N__26667;
    wire N__26666;
    wire N__26665;
    wire N__26664;
    wire N__26663;
    wire N__26662;
    wire N__26661;
    wire N__26654;
    wire N__26647;
    wire N__26644;
    wire N__26641;
    wire N__26638;
    wire N__26635;
    wire N__26628;
    wire N__26627;
    wire N__26626;
    wire N__26625;
    wire N__26624;
    wire N__26621;
    wire N__26620;
    wire N__26619;
    wire N__26618;
    wire N__26617;
    wire N__26616;
    wire N__26613;
    wire N__26608;
    wire N__26603;
    wire N__26602;
    wire N__26599;
    wire N__26594;
    wire N__26589;
    wire N__26584;
    wire N__26581;
    wire N__26576;
    wire N__26569;
    wire N__26564;
    wire N__26561;
    wire N__26558;
    wire N__26555;
    wire N__26552;
    wire N__26537;
    wire N__26528;
    wire N__26525;
    wire N__26522;
    wire N__26521;
    wire N__26520;
    wire N__26519;
    wire N__26518;
    wire N__26515;
    wire N__26512;
    wire N__26509;
    wire N__26508;
    wire N__26505;
    wire N__26502;
    wire N__26501;
    wire N__26500;
    wire N__26495;
    wire N__26492;
    wire N__26489;
    wire N__26486;
    wire N__26483;
    wire N__26480;
    wire N__26477;
    wire N__26476;
    wire N__26473;
    wire N__26466;
    wire N__26459;
    wire N__26456;
    wire N__26455;
    wire N__26450;
    wire N__26445;
    wire N__26442;
    wire N__26439;
    wire N__26432;
    wire N__26429;
    wire N__26426;
    wire N__26423;
    wire N__26420;
    wire N__26417;
    wire N__26416;
    wire N__26413;
    wire N__26410;
    wire N__26409;
    wire N__26406;
    wire N__26405;
    wire N__26404;
    wire N__26401;
    wire N__26400;
    wire N__26397;
    wire N__26394;
    wire N__26391;
    wire N__26388;
    wire N__26385;
    wire N__26382;
    wire N__26379;
    wire N__26378;
    wire N__26377;
    wire N__26374;
    wire N__26371;
    wire N__26368;
    wire N__26365;
    wire N__26362;
    wire N__26359;
    wire N__26356;
    wire N__26353;
    wire N__26350;
    wire N__26347;
    wire N__26344;
    wire N__26341;
    wire N__26338;
    wire N__26335;
    wire N__26318;
    wire N__26315;
    wire N__26312;
    wire N__26309;
    wire N__26306;
    wire N__26303;
    wire N__26300;
    wire N__26297;
    wire N__26294;
    wire N__26291;
    wire N__26288;
    wire N__26285;
    wire N__26282;
    wire N__26279;
    wire N__26276;
    wire N__26273;
    wire N__26270;
    wire N__26267;
    wire N__26264;
    wire N__26261;
    wire N__26260;
    wire N__26257;
    wire N__26254;
    wire N__26251;
    wire N__26246;
    wire N__26243;
    wire N__26240;
    wire N__26237;
    wire N__26234;
    wire N__26231;
    wire N__26228;
    wire N__26225;
    wire N__26222;
    wire N__26221;
    wire N__26218;
    wire N__26215;
    wire N__26212;
    wire N__26207;
    wire N__26204;
    wire N__26201;
    wire N__26200;
    wire N__26197;
    wire N__26194;
    wire N__26191;
    wire N__26186;
    wire N__26185;
    wire N__26182;
    wire N__26181;
    wire N__26180;
    wire N__26177;
    wire N__26174;
    wire N__26171;
    wire N__26170;
    wire N__26169;
    wire N__26168;
    wire N__26167;
    wire N__26164;
    wire N__26161;
    wire N__26156;
    wire N__26153;
    wire N__26144;
    wire N__26135;
    wire N__26132;
    wire N__26131;
    wire N__26130;
    wire N__26129;
    wire N__26126;
    wire N__26121;
    wire N__26120;
    wire N__26119;
    wire N__26118;
    wire N__26115;
    wire N__26110;
    wire N__26103;
    wire N__26100;
    wire N__26093;
    wire N__26090;
    wire N__26087;
    wire N__26084;
    wire N__26081;
    wire N__26078;
    wire N__26075;
    wire N__26072;
    wire N__26069;
    wire N__26066;
    wire N__26063;
    wire N__26060;
    wire N__26057;
    wire N__26054;
    wire N__26051;
    wire N__26048;
    wire N__26045;
    wire N__26042;
    wire N__26039;
    wire N__26036;
    wire N__26035;
    wire N__26032;
    wire N__26029;
    wire N__26026;
    wire N__26021;
    wire N__26018;
    wire N__26015;
    wire N__26012;
    wire N__26009;
    wire N__26006;
    wire N__26003;
    wire N__26000;
    wire N__25999;
    wire N__25996;
    wire N__25993;
    wire N__25990;
    wire N__25985;
    wire N__25982;
    wire N__25979;
    wire N__25978;
    wire N__25975;
    wire N__25972;
    wire N__25969;
    wire N__25964;
    wire N__25961;
    wire N__25958;
    wire N__25955;
    wire N__25952;
    wire N__25949;
    wire N__25946;
    wire N__25943;
    wire N__25942;
    wire N__25939;
    wire N__25936;
    wire N__25935;
    wire N__25932;
    wire N__25927;
    wire N__25926;
    wire N__25923;
    wire N__25920;
    wire N__25917;
    wire N__25910;
    wire N__25907;
    wire N__25906;
    wire N__25905;
    wire N__25902;
    wire N__25897;
    wire N__25892;
    wire N__25889;
    wire N__25888;
    wire N__25885;
    wire N__25884;
    wire N__25881;
    wire N__25878;
    wire N__25875;
    wire N__25872;
    wire N__25871;
    wire N__25866;
    wire N__25863;
    wire N__25860;
    wire N__25857;
    wire N__25854;
    wire N__25847;
    wire N__25844;
    wire N__25841;
    wire N__25838;
    wire N__25835;
    wire N__25832;
    wire N__25831;
    wire N__25828;
    wire N__25825;
    wire N__25822;
    wire N__25819;
    wire N__25816;
    wire N__25811;
    wire N__25810;
    wire N__25807;
    wire N__25804;
    wire N__25801;
    wire N__25796;
    wire N__25793;
    wire N__25790;
    wire N__25789;
    wire N__25786;
    wire N__25783;
    wire N__25778;
    wire N__25777;
    wire N__25774;
    wire N__25771;
    wire N__25766;
    wire N__25765;
    wire N__25760;
    wire N__25757;
    wire N__25754;
    wire N__25751;
    wire N__25748;
    wire N__25745;
    wire N__25742;
    wire N__25739;
    wire N__25736;
    wire N__25733;
    wire N__25730;
    wire N__25727;
    wire N__25724;
    wire N__25723;
    wire N__25720;
    wire N__25717;
    wire N__25714;
    wire N__25711;
    wire N__25710;
    wire N__25705;
    wire N__25702;
    wire N__25699;
    wire N__25694;
    wire N__25691;
    wire N__25688;
    wire N__25687;
    wire N__25684;
    wire N__25681;
    wire N__25678;
    wire N__25673;
    wire N__25670;
    wire N__25669;
    wire N__25666;
    wire N__25663;
    wire N__25658;
    wire N__25655;
    wire N__25652;
    wire N__25651;
    wire N__25648;
    wire N__25645;
    wire N__25642;
    wire N__25637;
    wire N__25636;
    wire N__25635;
    wire N__25632;
    wire N__25631;
    wire N__25628;
    wire N__25625;
    wire N__25622;
    wire N__25619;
    wire N__25614;
    wire N__25611;
    wire N__25608;
    wire N__25605;
    wire N__25600;
    wire N__25597;
    wire N__25594;
    wire N__25589;
    wire N__25588;
    wire N__25587;
    wire N__25584;
    wire N__25583;
    wire N__25582;
    wire N__25579;
    wire N__25576;
    wire N__25573;
    wire N__25570;
    wire N__25567;
    wire N__25564;
    wire N__25561;
    wire N__25556;
    wire N__25555;
    wire N__25550;
    wire N__25545;
    wire N__25542;
    wire N__25539;
    wire N__25536;
    wire N__25529;
    wire N__25526;
    wire N__25525;
    wire N__25522;
    wire N__25519;
    wire N__25516;
    wire N__25513;
    wire N__25510;
    wire N__25507;
    wire N__25502;
    wire N__25501;
    wire N__25498;
    wire N__25495;
    wire N__25492;
    wire N__25489;
    wire N__25486;
    wire N__25483;
    wire N__25480;
    wire N__25475;
    wire N__25472;
    wire N__25471;
    wire N__25468;
    wire N__25465;
    wire N__25462;
    wire N__25461;
    wire N__25458;
    wire N__25455;
    wire N__25452;
    wire N__25445;
    wire N__25444;
    wire N__25443;
    wire N__25440;
    wire N__25437;
    wire N__25434;
    wire N__25433;
    wire N__25432;
    wire N__25429;
    wire N__25424;
    wire N__25421;
    wire N__25418;
    wire N__25413;
    wire N__25410;
    wire N__25403;
    wire N__25400;
    wire N__25399;
    wire N__25396;
    wire N__25393;
    wire N__25390;
    wire N__25389;
    wire N__25386;
    wire N__25385;
    wire N__25382;
    wire N__25379;
    wire N__25376;
    wire N__25373;
    wire N__25366;
    wire N__25361;
    wire N__25358;
    wire N__25355;
    wire N__25352;
    wire N__25349;
    wire N__25346;
    wire N__25345;
    wire N__25342;
    wire N__25339;
    wire N__25336;
    wire N__25333;
    wire N__25332;
    wire N__25331;
    wire N__25326;
    wire N__25321;
    wire N__25316;
    wire N__25313;
    wire N__25310;
    wire N__25309;
    wire N__25306;
    wire N__25303;
    wire N__25300;
    wire N__25295;
    wire N__25292;
    wire N__25289;
    wire N__25286;
    wire N__25283;
    wire N__25280;
    wire N__25277;
    wire N__25274;
    wire N__25273;
    wire N__25272;
    wire N__25271;
    wire N__25270;
    wire N__25267;
    wire N__25264;
    wire N__25263;
    wire N__25260;
    wire N__25257;
    wire N__25254;
    wire N__25251;
    wire N__25248;
    wire N__25241;
    wire N__25232;
    wire N__25229;
    wire N__25226;
    wire N__25223;
    wire N__25220;
    wire N__25217;
    wire N__25214;
    wire N__25211;
    wire N__25208;
    wire N__25207;
    wire N__25204;
    wire N__25201;
    wire N__25198;
    wire N__25193;
    wire N__25190;
    wire N__25189;
    wire N__25186;
    wire N__25183;
    wire N__25178;
    wire N__25175;
    wire N__25174;
    wire N__25171;
    wire N__25168;
    wire N__25165;
    wire N__25162;
    wire N__25159;
    wire N__25156;
    wire N__25153;
    wire N__25150;
    wire N__25145;
    wire N__25142;
    wire N__25139;
    wire N__25136;
    wire N__25133;
    wire N__25132;
    wire N__25129;
    wire N__25126;
    wire N__25123;
    wire N__25120;
    wire N__25117;
    wire N__25112;
    wire N__25109;
    wire N__25108;
    wire N__25107;
    wire N__25106;
    wire N__25103;
    wire N__25100;
    wire N__25097;
    wire N__25094;
    wire N__25089;
    wire N__25086;
    wire N__25083;
    wire N__25080;
    wire N__25073;
    wire N__25070;
    wire N__25067;
    wire N__25064;
    wire N__25063;
    wire N__25062;
    wire N__25059;
    wire N__25056;
    wire N__25053;
    wire N__25052;
    wire N__25049;
    wire N__25046;
    wire N__25043;
    wire N__25040;
    wire N__25037;
    wire N__25032;
    wire N__25025;
    wire N__25022;
    wire N__25021;
    wire N__25018;
    wire N__25015;
    wire N__25012;
    wire N__25009;
    wire N__25006;
    wire N__25003;
    wire N__25000;
    wire N__24995;
    wire N__24994;
    wire N__24991;
    wire N__24988;
    wire N__24985;
    wire N__24982;
    wire N__24979;
    wire N__24976;
    wire N__24971;
    wire N__24970;
    wire N__24967;
    wire N__24964;
    wire N__24963;
    wire N__24960;
    wire N__24957;
    wire N__24956;
    wire N__24955;
    wire N__24952;
    wire N__24947;
    wire N__24942;
    wire N__24935;
    wire N__24932;
    wire N__24931;
    wire N__24928;
    wire N__24925;
    wire N__24922;
    wire N__24919;
    wire N__24916;
    wire N__24911;
    wire N__24908;
    wire N__24905;
    wire N__24902;
    wire N__24901;
    wire N__24900;
    wire N__24897;
    wire N__24894;
    wire N__24891;
    wire N__24884;
    wire N__24883;
    wire N__24880;
    wire N__24879;
    wire N__24876;
    wire N__24873;
    wire N__24870;
    wire N__24867;
    wire N__24864;
    wire N__24861;
    wire N__24856;
    wire N__24853;
    wire N__24848;
    wire N__24845;
    wire N__24842;
    wire N__24839;
    wire N__24838;
    wire N__24835;
    wire N__24832;
    wire N__24829;
    wire N__24826;
    wire N__24821;
    wire N__24818;
    wire N__24815;
    wire N__24812;
    wire N__24809;
    wire N__24806;
    wire N__24803;
    wire N__24800;
    wire N__24797;
    wire N__24794;
    wire N__24791;
    wire N__24790;
    wire N__24785;
    wire N__24782;
    wire N__24781;
    wire N__24778;
    wire N__24775;
    wire N__24772;
    wire N__24769;
    wire N__24764;
    wire N__24763;
    wire N__24760;
    wire N__24759;
    wire N__24758;
    wire N__24755;
    wire N__24754;
    wire N__24753;
    wire N__24750;
    wire N__24747;
    wire N__24744;
    wire N__24741;
    wire N__24736;
    wire N__24733;
    wire N__24730;
    wire N__24725;
    wire N__24722;
    wire N__24721;
    wire N__24720;
    wire N__24715;
    wire N__24710;
    wire N__24705;
    wire N__24698;
    wire N__24695;
    wire N__24694;
    wire N__24693;
    wire N__24692;
    wire N__24691;
    wire N__24688;
    wire N__24683;
    wire N__24682;
    wire N__24679;
    wire N__24678;
    wire N__24677;
    wire N__24674;
    wire N__24673;
    wire N__24670;
    wire N__24667;
    wire N__24660;
    wire N__24657;
    wire N__24654;
    wire N__24651;
    wire N__24648;
    wire N__24643;
    wire N__24640;
    wire N__24637;
    wire N__24634;
    wire N__24631;
    wire N__24628;
    wire N__24621;
    wire N__24614;
    wire N__24611;
    wire N__24608;
    wire N__24605;
    wire N__24602;
    wire N__24599;
    wire N__24598;
    wire N__24595;
    wire N__24594;
    wire N__24591;
    wire N__24588;
    wire N__24585;
    wire N__24578;
    wire N__24575;
    wire N__24572;
    wire N__24569;
    wire N__24566;
    wire N__24563;
    wire N__24560;
    wire N__24557;
    wire N__24556;
    wire N__24555;
    wire N__24552;
    wire N__24549;
    wire N__24546;
    wire N__24543;
    wire N__24540;
    wire N__24537;
    wire N__24532;
    wire N__24529;
    wire N__24524;
    wire N__24523;
    wire N__24520;
    wire N__24517;
    wire N__24514;
    wire N__24509;
    wire N__24506;
    wire N__24503;
    wire N__24500;
    wire N__24499;
    wire N__24496;
    wire N__24493;
    wire N__24490;
    wire N__24487;
    wire N__24482;
    wire N__24479;
    wire N__24476;
    wire N__24473;
    wire N__24470;
    wire N__24467;
    wire N__24464;
    wire N__24461;
    wire N__24458;
    wire N__24455;
    wire N__24452;
    wire N__24449;
    wire N__24446;
    wire N__24443;
    wire N__24440;
    wire N__24439;
    wire N__24438;
    wire N__24435;
    wire N__24430;
    wire N__24427;
    wire N__24424;
    wire N__24419;
    wire N__24416;
    wire N__24415;
    wire N__24412;
    wire N__24409;
    wire N__24406;
    wire N__24403;
    wire N__24400;
    wire N__24395;
    wire N__24392;
    wire N__24389;
    wire N__24386;
    wire N__24383;
    wire N__24380;
    wire N__24379;
    wire N__24378;
    wire N__24377;
    wire N__24374;
    wire N__24371;
    wire N__24370;
    wire N__24367;
    wire N__24364;
    wire N__24361;
    wire N__24358;
    wire N__24355;
    wire N__24344;
    wire N__24343;
    wire N__24340;
    wire N__24337;
    wire N__24332;
    wire N__24329;
    wire N__24326;
    wire N__24323;
    wire N__24320;
    wire N__24319;
    wire N__24318;
    wire N__24317;
    wire N__24316;
    wire N__24315;
    wire N__24310;
    wire N__24307;
    wire N__24304;
    wire N__24299;
    wire N__24294;
    wire N__24291;
    wire N__24284;
    wire N__24281;
    wire N__24278;
    wire N__24277;
    wire N__24276;
    wire N__24275;
    wire N__24274;
    wire N__24273;
    wire N__24272;
    wire N__24271;
    wire N__24270;
    wire N__24269;
    wire N__24268;
    wire N__24267;
    wire N__24266;
    wire N__24265;
    wire N__24264;
    wire N__24263;
    wire N__24262;
    wire N__24261;
    wire N__24260;
    wire N__24259;
    wire N__24258;
    wire N__24257;
    wire N__24256;
    wire N__24255;
    wire N__24254;
    wire N__24253;
    wire N__24252;
    wire N__24251;
    wire N__24250;
    wire N__24247;
    wire N__24246;
    wire N__24245;
    wire N__24244;
    wire N__24243;
    wire N__24242;
    wire N__24241;
    wire N__24240;
    wire N__24239;
    wire N__24238;
    wire N__24237;
    wire N__24230;
    wire N__24227;
    wire N__24222;
    wire N__24219;
    wire N__24218;
    wire N__24217;
    wire N__24216;
    wire N__24215;
    wire N__24214;
    wire N__24213;
    wire N__24212;
    wire N__24205;
    wire N__24202;
    wire N__24193;
    wire N__24184;
    wire N__24181;
    wire N__24176;
    wire N__24171;
    wire N__24162;
    wire N__24159;
    wire N__24152;
    wire N__24143;
    wire N__24136;
    wire N__24131;
    wire N__24126;
    wire N__24125;
    wire N__24122;
    wire N__24119;
    wire N__24118;
    wire N__24115;
    wire N__24106;
    wire N__24103;
    wire N__24096;
    wire N__24091;
    wire N__24086;
    wire N__24073;
    wire N__24072;
    wire N__24071;
    wire N__24070;
    wire N__24069;
    wire N__24066;
    wire N__24061;
    wire N__24058;
    wire N__24049;
    wire N__24044;
    wire N__24041;
    wire N__24032;
    wire N__24025;
    wire N__24014;
    wire N__24011;
    wire N__24008;
    wire N__24007;
    wire N__24004;
    wire N__24003;
    wire N__24002;
    wire N__23999;
    wire N__23996;
    wire N__23991;
    wire N__23984;
    wire N__23981;
    wire N__23978;
    wire N__23977;
    wire N__23974;
    wire N__23973;
    wire N__23970;
    wire N__23969;
    wire N__23966;
    wire N__23959;
    wire N__23954;
    wire N__23951;
    wire N__23948;
    wire N__23947;
    wire N__23946;
    wire N__23945;
    wire N__23944;
    wire N__23941;
    wire N__23938;
    wire N__23931;
    wire N__23924;
    wire N__23921;
    wire N__23918;
    wire N__23915;
    wire N__23912;
    wire N__23909;
    wire N__23906;
    wire N__23905;
    wire N__23902;
    wire N__23899;
    wire N__23894;
    wire N__23893;
    wire N__23890;
    wire N__23887;
    wire N__23882;
    wire N__23881;
    wire N__23878;
    wire N__23877;
    wire N__23874;
    wire N__23873;
    wire N__23870;
    wire N__23867;
    wire N__23866;
    wire N__23863;
    wire N__23860;
    wire N__23859;
    wire N__23856;
    wire N__23853;
    wire N__23850;
    wire N__23845;
    wire N__23842;
    wire N__23831;
    wire N__23830;
    wire N__23827;
    wire N__23824;
    wire N__23823;
    wire N__23820;
    wire N__23817;
    wire N__23814;
    wire N__23811;
    wire N__23804;
    wire N__23801;
    wire N__23798;
    wire N__23795;
    wire N__23794;
    wire N__23793;
    wire N__23790;
    wire N__23787;
    wire N__23784;
    wire N__23777;
    wire N__23774;
    wire N__23773;
    wire N__23770;
    wire N__23767;
    wire N__23764;
    wire N__23761;
    wire N__23756;
    wire N__23753;
    wire N__23750;
    wire N__23747;
    wire N__23744;
    wire N__23741;
    wire N__23738;
    wire N__23737;
    wire N__23736;
    wire N__23733;
    wire N__23730;
    wire N__23727;
    wire N__23720;
    wire N__23717;
    wire N__23714;
    wire N__23711;
    wire N__23708;
    wire N__23705;
    wire N__23702;
    wire N__23699;
    wire N__23698;
    wire N__23695;
    wire N__23692;
    wire N__23689;
    wire N__23686;
    wire N__23683;
    wire N__23680;
    wire N__23679;
    wire N__23678;
    wire N__23675;
    wire N__23672;
    wire N__23669;
    wire N__23666;
    wire N__23663;
    wire N__23654;
    wire N__23651;
    wire N__23648;
    wire N__23645;
    wire N__23642;
    wire N__23641;
    wire N__23638;
    wire N__23635;
    wire N__23632;
    wire N__23627;
    wire N__23624;
    wire N__23621;
    wire N__23618;
    wire N__23615;
    wire N__23612;
    wire N__23609;
    wire N__23606;
    wire N__23603;
    wire N__23600;
    wire N__23597;
    wire N__23594;
    wire N__23591;
    wire N__23588;
    wire N__23585;
    wire N__23582;
    wire N__23579;
    wire N__23576;
    wire N__23573;
    wire N__23570;
    wire N__23567;
    wire N__23564;
    wire N__23561;
    wire N__23558;
    wire N__23555;
    wire N__23552;
    wire N__23549;
    wire N__23546;
    wire N__23543;
    wire N__23540;
    wire N__23537;
    wire N__23534;
    wire N__23531;
    wire N__23528;
    wire N__23527;
    wire N__23524;
    wire N__23521;
    wire N__23516;
    wire N__23513;
    wire N__23510;
    wire N__23509;
    wire N__23506;
    wire N__23503;
    wire N__23500;
    wire N__23497;
    wire N__23492;
    wire N__23491;
    wire N__23488;
    wire N__23485;
    wire N__23480;
    wire N__23477;
    wire N__23474;
    wire N__23471;
    wire N__23468;
    wire N__23465;
    wire N__23464;
    wire N__23461;
    wire N__23458;
    wire N__23455;
    wire N__23450;
    wire N__23447;
    wire N__23444;
    wire N__23441;
    wire N__23438;
    wire N__23435;
    wire N__23432;
    wire N__23431;
    wire N__23428;
    wire N__23425;
    wire N__23420;
    wire N__23419;
    wire N__23416;
    wire N__23413;
    wire N__23410;
    wire N__23405;
    wire N__23402;
    wire N__23399;
    wire N__23396;
    wire N__23393;
    wire N__23390;
    wire N__23387;
    wire N__23384;
    wire N__23381;
    wire N__23378;
    wire N__23377;
    wire N__23374;
    wire N__23371;
    wire N__23368;
    wire N__23363;
    wire N__23362;
    wire N__23359;
    wire N__23356;
    wire N__23351;
    wire N__23350;
    wire N__23347;
    wire N__23344;
    wire N__23341;
    wire N__23336;
    wire N__23333;
    wire N__23330;
    wire N__23329;
    wire N__23326;
    wire N__23323;
    wire N__23320;
    wire N__23315;
    wire N__23312;
    wire N__23311;
    wire N__23308;
    wire N__23305;
    wire N__23300;
    wire N__23299;
    wire N__23296;
    wire N__23293;
    wire N__23288;
    wire N__23285;
    wire N__23282;
    wire N__23279;
    wire N__23276;
    wire N__23273;
    wire N__23270;
    wire N__23267;
    wire N__23264;
    wire N__23263;
    wire N__23260;
    wire N__23257;
    wire N__23252;
    wire N__23249;
    wire N__23246;
    wire N__23243;
    wire N__23242;
    wire N__23239;
    wire N__23236;
    wire N__23233;
    wire N__23228;
    wire N__23225;
    wire N__23222;
    wire N__23219;
    wire N__23216;
    wire N__23213;
    wire N__23210;
    wire N__23207;
    wire N__23206;
    wire N__23203;
    wire N__23200;
    wire N__23199;
    wire N__23198;
    wire N__23195;
    wire N__23192;
    wire N__23187;
    wire N__23184;
    wire N__23181;
    wire N__23174;
    wire N__23171;
    wire N__23168;
    wire N__23165;
    wire N__23162;
    wire N__23159;
    wire N__23156;
    wire N__23153;
    wire N__23150;
    wire N__23147;
    wire N__23144;
    wire N__23141;
    wire N__23138;
    wire N__23135;
    wire N__23132;
    wire N__23129;
    wire N__23126;
    wire N__23125;
    wire N__23122;
    wire N__23119;
    wire N__23116;
    wire N__23113;
    wire N__23108;
    wire N__23105;
    wire N__23102;
    wire N__23099;
    wire N__23098;
    wire N__23095;
    wire N__23092;
    wire N__23087;
    wire N__23084;
    wire N__23083;
    wire N__23080;
    wire N__23077;
    wire N__23072;
    wire N__23069;
    wire N__23066;
    wire N__23065;
    wire N__23062;
    wire N__23059;
    wire N__23056;
    wire N__23051;
    wire N__23050;
    wire N__23047;
    wire N__23044;
    wire N__23043;
    wire N__23040;
    wire N__23037;
    wire N__23034;
    wire N__23029;
    wire N__23024;
    wire N__23023;
    wire N__23022;
    wire N__23019;
    wire N__23016;
    wire N__23013;
    wire N__23010;
    wire N__23007;
    wire N__23004;
    wire N__23001;
    wire N__22998;
    wire N__22991;
    wire N__22988;
    wire N__22985;
    wire N__22982;
    wire N__22979;
    wire N__22976;
    wire N__22973;
    wire N__22970;
    wire N__22967;
    wire N__22964;
    wire N__22961;
    wire N__22960;
    wire N__22957;
    wire N__22954;
    wire N__22953;
    wire N__22952;
    wire N__22949;
    wire N__22946;
    wire N__22943;
    wire N__22940;
    wire N__22935;
    wire N__22928;
    wire N__22927;
    wire N__22926;
    wire N__22925;
    wire N__22922;
    wire N__22917;
    wire N__22914;
    wire N__22909;
    wire N__22904;
    wire N__22903;
    wire N__22902;
    wire N__22897;
    wire N__22894;
    wire N__22893;
    wire N__22890;
    wire N__22887;
    wire N__22884;
    wire N__22881;
    wire N__22876;
    wire N__22871;
    wire N__22870;
    wire N__22865;
    wire N__22862;
    wire N__22859;
    wire N__22856;
    wire N__22853;
    wire N__22850;
    wire N__22847;
    wire N__22846;
    wire N__22843;
    wire N__22840;
    wire N__22839;
    wire N__22836;
    wire N__22833;
    wire N__22832;
    wire N__22831;
    wire N__22828;
    wire N__22823;
    wire N__22820;
    wire N__22817;
    wire N__22814;
    wire N__22805;
    wire N__22802;
    wire N__22801;
    wire N__22798;
    wire N__22795;
    wire N__22792;
    wire N__22789;
    wire N__22784;
    wire N__22783;
    wire N__22780;
    wire N__22777;
    wire N__22774;
    wire N__22769;
    wire N__22768;
    wire N__22767;
    wire N__22762;
    wire N__22759;
    wire N__22756;
    wire N__22755;
    wire N__22752;
    wire N__22749;
    wire N__22746;
    wire N__22739;
    wire N__22736;
    wire N__22733;
    wire N__22730;
    wire N__22729;
    wire N__22726;
    wire N__22723;
    wire N__22718;
    wire N__22715;
    wire N__22712;
    wire N__22709;
    wire N__22706;
    wire N__22705;
    wire N__22702;
    wire N__22699;
    wire N__22696;
    wire N__22695;
    wire N__22692;
    wire N__22689;
    wire N__22686;
    wire N__22683;
    wire N__22680;
    wire N__22677;
    wire N__22670;
    wire N__22669;
    wire N__22668;
    wire N__22665;
    wire N__22662;
    wire N__22659;
    wire N__22654;
    wire N__22653;
    wire N__22650;
    wire N__22647;
    wire N__22644;
    wire N__22637;
    wire N__22636;
    wire N__22635;
    wire N__22632;
    wire N__22629;
    wire N__22628;
    wire N__22627;
    wire N__22624;
    wire N__22621;
    wire N__22618;
    wire N__22615;
    wire N__22612;
    wire N__22609;
    wire N__22604;
    wire N__22595;
    wire N__22592;
    wire N__22591;
    wire N__22590;
    wire N__22587;
    wire N__22584;
    wire N__22581;
    wire N__22580;
    wire N__22577;
    wire N__22574;
    wire N__22571;
    wire N__22568;
    wire N__22563;
    wire N__22560;
    wire N__22553;
    wire N__22552;
    wire N__22549;
    wire N__22548;
    wire N__22545;
    wire N__22544;
    wire N__22543;
    wire N__22542;
    wire N__22539;
    wire N__22536;
    wire N__22533;
    wire N__22530;
    wire N__22525;
    wire N__22518;
    wire N__22511;
    wire N__22508;
    wire N__22505;
    wire N__22502;
    wire N__22499;
    wire N__22496;
    wire N__22493;
    wire N__22492;
    wire N__22489;
    wire N__22486;
    wire N__22485;
    wire N__22484;
    wire N__22481;
    wire N__22480;
    wire N__22477;
    wire N__22474;
    wire N__22471;
    wire N__22468;
    wire N__22465;
    wire N__22460;
    wire N__22451;
    wire N__22450;
    wire N__22447;
    wire N__22444;
    wire N__22441;
    wire N__22438;
    wire N__22433;
    wire N__22430;
    wire N__22427;
    wire N__22424;
    wire N__22421;
    wire N__22420;
    wire N__22417;
    wire N__22414;
    wire N__22411;
    wire N__22406;
    wire N__22405;
    wire N__22402;
    wire N__22399;
    wire N__22396;
    wire N__22393;
    wire N__22390;
    wire N__22387;
    wire N__22382;
    wire N__22379;
    wire N__22376;
    wire N__22375;
    wire N__22372;
    wire N__22369;
    wire N__22366;
    wire N__22361;
    wire N__22358;
    wire N__22355;
    wire N__22352;
    wire N__22349;
    wire N__22346;
    wire N__22345;
    wire N__22342;
    wire N__22339;
    wire N__22334;
    wire N__22333;
    wire N__22330;
    wire N__22327;
    wire N__22324;
    wire N__22321;
    wire N__22316;
    wire N__22313;
    wire N__22310;
    wire N__22307;
    wire N__22304;
    wire N__22301;
    wire N__22298;
    wire N__22297;
    wire N__22296;
    wire N__22293;
    wire N__22288;
    wire N__22285;
    wire N__22280;
    wire N__22277;
    wire N__22274;
    wire N__22273;
    wire N__22270;
    wire N__22267;
    wire N__22262;
    wire N__22261;
    wire N__22258;
    wire N__22255;
    wire N__22250;
    wire N__22247;
    wire N__22244;
    wire N__22241;
    wire N__22238;
    wire N__22235;
    wire N__22232;
    wire N__22229;
    wire N__22226;
    wire N__22225;
    wire N__22224;
    wire N__22221;
    wire N__22218;
    wire N__22215;
    wire N__22212;
    wire N__22209;
    wire N__22202;
    wire N__22201;
    wire N__22196;
    wire N__22193;
    wire N__22190;
    wire N__22187;
    wire N__22184;
    wire N__22183;
    wire N__22180;
    wire N__22177;
    wire N__22172;
    wire N__22169;
    wire N__22168;
    wire N__22165;
    wire N__22162;
    wire N__22161;
    wire N__22156;
    wire N__22155;
    wire N__22152;
    wire N__22149;
    wire N__22146;
    wire N__22139;
    wire N__22138;
    wire N__22135;
    wire N__22134;
    wire N__22133;
    wire N__22130;
    wire N__22127;
    wire N__22124;
    wire N__22121;
    wire N__22114;
    wire N__22111;
    wire N__22108;
    wire N__22103;
    wire N__22102;
    wire N__22099;
    wire N__22098;
    wire N__22095;
    wire N__22092;
    wire N__22087;
    wire N__22086;
    wire N__22083;
    wire N__22080;
    wire N__22077;
    wire N__22074;
    wire N__22071;
    wire N__22064;
    wire N__22063;
    wire N__22060;
    wire N__22059;
    wire N__22056;
    wire N__22049;
    wire N__22046;
    wire N__22043;
    wire N__22042;
    wire N__22041;
    wire N__22038;
    wire N__22035;
    wire N__22034;
    wire N__22033;
    wire N__22030;
    wire N__22027;
    wire N__22022;
    wire N__22017;
    wire N__22010;
    wire N__22009;
    wire N__22006;
    wire N__22003;
    wire N__22002;
    wire N__21999;
    wire N__21996;
    wire N__21993;
    wire N__21990;
    wire N__21985;
    wire N__21982;
    wire N__21977;
    wire N__21976;
    wire N__21973;
    wire N__21970;
    wire N__21967;
    wire N__21964;
    wire N__21961;
    wire N__21958;
    wire N__21953;
    wire N__21950;
    wire N__21947;
    wire N__21946;
    wire N__21943;
    wire N__21940;
    wire N__21937;
    wire N__21934;
    wire N__21929;
    wire N__21928;
    wire N__21925;
    wire N__21922;
    wire N__21919;
    wire N__21916;
    wire N__21913;
    wire N__21908;
    wire N__21907;
    wire N__21906;
    wire N__21905;
    wire N__21902;
    wire N__21899;
    wire N__21896;
    wire N__21895;
    wire N__21892;
    wire N__21885;
    wire N__21882;
    wire N__21877;
    wire N__21874;
    wire N__21869;
    wire N__21868;
    wire N__21865;
    wire N__21862;
    wire N__21859;
    wire N__21858;
    wire N__21857;
    wire N__21854;
    wire N__21851;
    wire N__21846;
    wire N__21839;
    wire N__21838;
    wire N__21837;
    wire N__21834;
    wire N__21833;
    wire N__21830;
    wire N__21829;
    wire N__21826;
    wire N__21823;
    wire N__21820;
    wire N__21817;
    wire N__21814;
    wire N__21811;
    wire N__21808;
    wire N__21805;
    wire N__21802;
    wire N__21795;
    wire N__21790;
    wire N__21785;
    wire N__21782;
    wire N__21779;
    wire N__21776;
    wire N__21773;
    wire N__21772;
    wire N__21769;
    wire N__21768;
    wire N__21765;
    wire N__21764;
    wire N__21761;
    wire N__21758;
    wire N__21755;
    wire N__21754;
    wire N__21751;
    wire N__21748;
    wire N__21745;
    wire N__21742;
    wire N__21737;
    wire N__21728;
    wire N__21727;
    wire N__21724;
    wire N__21723;
    wire N__21722;
    wire N__21719;
    wire N__21718;
    wire N__21715;
    wire N__21712;
    wire N__21709;
    wire N__21706;
    wire N__21703;
    wire N__21700;
    wire N__21689;
    wire N__21686;
    wire N__21685;
    wire N__21684;
    wire N__21683;
    wire N__21680;
    wire N__21677;
    wire N__21674;
    wire N__21671;
    wire N__21668;
    wire N__21665;
    wire N__21662;
    wire N__21653;
    wire N__21650;
    wire N__21647;
    wire N__21646;
    wire N__21645;
    wire N__21642;
    wire N__21637;
    wire N__21632;
    wire N__21629;
    wire N__21628;
    wire N__21625;
    wire N__21624;
    wire N__21621;
    wire N__21618;
    wire N__21615;
    wire N__21608;
    wire N__21607;
    wire N__21606;
    wire N__21605;
    wire N__21602;
    wire N__21599;
    wire N__21596;
    wire N__21593;
    wire N__21592;
    wire N__21589;
    wire N__21584;
    wire N__21583;
    wire N__21582;
    wire N__21579;
    wire N__21576;
    wire N__21573;
    wire N__21570;
    wire N__21565;
    wire N__21554;
    wire N__21553;
    wire N__21552;
    wire N__21549;
    wire N__21546;
    wire N__21543;
    wire N__21540;
    wire N__21533;
    wire N__21530;
    wire N__21527;
    wire N__21524;
    wire N__21523;
    wire N__21520;
    wire N__21517;
    wire N__21512;
    wire N__21509;
    wire N__21506;
    wire N__21505;
    wire N__21502;
    wire N__21501;
    wire N__21500;
    wire N__21497;
    wire N__21494;
    wire N__21491;
    wire N__21488;
    wire N__21479;
    wire N__21476;
    wire N__21473;
    wire N__21470;
    wire N__21469;
    wire N__21468;
    wire N__21467;
    wire N__21466;
    wire N__21465;
    wire N__21462;
    wire N__21455;
    wire N__21452;
    wire N__21449;
    wire N__21444;
    wire N__21437;
    wire N__21434;
    wire N__21433;
    wire N__21432;
    wire N__21431;
    wire N__21430;
    wire N__21427;
    wire N__21426;
    wire N__21425;
    wire N__21422;
    wire N__21421;
    wire N__21418;
    wire N__21417;
    wire N__21416;
    wire N__21415;
    wire N__21414;
    wire N__21413;
    wire N__21412;
    wire N__21411;
    wire N__21410;
    wire N__21409;
    wire N__21406;
    wire N__21401;
    wire N__21398;
    wire N__21391;
    wire N__21382;
    wire N__21379;
    wire N__21368;
    wire N__21365;
    wire N__21360;
    wire N__21347;
    wire N__21344;
    wire N__21343;
    wire N__21342;
    wire N__21341;
    wire N__21340;
    wire N__21337;
    wire N__21330;
    wire N__21327;
    wire N__21326;
    wire N__21325;
    wire N__21324;
    wire N__21323;
    wire N__21320;
    wire N__21315;
    wire N__21312;
    wire N__21305;
    wire N__21296;
    wire N__21295;
    wire N__21294;
    wire N__21293;
    wire N__21292;
    wire N__21289;
    wire N__21288;
    wire N__21285;
    wire N__21284;
    wire N__21283;
    wire N__21280;
    wire N__21279;
    wire N__21276;
    wire N__21267;
    wire N__21266;
    wire N__21261;
    wire N__21258;
    wire N__21255;
    wire N__21250;
    wire N__21247;
    wire N__21236;
    wire N__21233;
    wire N__21232;
    wire N__21229;
    wire N__21226;
    wire N__21221;
    wire N__21218;
    wire N__21215;
    wire N__21212;
    wire N__21209;
    wire N__21206;
    wire N__21205;
    wire N__21202;
    wire N__21199;
    wire N__21196;
    wire N__21191;
    wire N__21188;
    wire N__21185;
    wire N__21182;
    wire N__21179;
    wire N__21176;
    wire N__21173;
    wire N__21170;
    wire N__21167;
    wire N__21164;
    wire N__21161;
    wire N__21158;
    wire N__21155;
    wire N__21152;
    wire N__21149;
    wire N__21148;
    wire N__21145;
    wire N__21142;
    wire N__21139;
    wire N__21136;
    wire N__21135;
    wire N__21130;
    wire N__21127;
    wire N__21122;
    wire N__21119;
    wire N__21116;
    wire N__21113;
    wire N__21110;
    wire N__21107;
    wire N__21104;
    wire N__21101;
    wire N__21098;
    wire N__21095;
    wire N__21092;
    wire N__21089;
    wire N__21086;
    wire N__21083;
    wire N__21080;
    wire N__21077;
    wire N__21074;
    wire N__21073;
    wire N__21068;
    wire N__21065;
    wire N__21064;
    wire N__21061;
    wire N__21058;
    wire N__21053;
    wire N__21050;
    wire N__21047;
    wire N__21044;
    wire N__21041;
    wire N__21038;
    wire N__21035;
    wire N__21032;
    wire N__21029;
    wire N__21026;
    wire N__21023;
    wire N__21020;
    wire N__21017;
    wire N__21014;
    wire N__21011;
    wire N__21008;
    wire N__21005;
    wire N__21002;
    wire N__20999;
    wire N__20996;
    wire N__20995;
    wire N__20992;
    wire N__20989;
    wire N__20986;
    wire N__20981;
    wire N__20980;
    wire N__20977;
    wire N__20974;
    wire N__20971;
    wire N__20966;
    wire N__20963;
    wire N__20960;
    wire N__20959;
    wire N__20956;
    wire N__20953;
    wire N__20950;
    wire N__20945;
    wire N__20942;
    wire N__20939;
    wire N__20938;
    wire N__20935;
    wire N__20932;
    wire N__20929;
    wire N__20924;
    wire N__20923;
    wire N__20920;
    wire N__20917;
    wire N__20912;
    wire N__20909;
    wire N__20906;
    wire N__20905;
    wire N__20902;
    wire N__20899;
    wire N__20894;
    wire N__20891;
    wire N__20888;
    wire N__20885;
    wire N__20882;
    wire N__20879;
    wire N__20876;
    wire N__20873;
    wire N__20870;
    wire N__20867;
    wire N__20864;
    wire N__20861;
    wire N__20858;
    wire N__20855;
    wire N__20852;
    wire N__20849;
    wire N__20846;
    wire N__20843;
    wire N__20840;
    wire N__20837;
    wire N__20834;
    wire N__20831;
    wire N__20830;
    wire N__20827;
    wire N__20824;
    wire N__20821;
    wire N__20816;
    wire N__20813;
    wire N__20812;
    wire N__20809;
    wire N__20806;
    wire N__20803;
    wire N__20798;
    wire N__20795;
    wire N__20792;
    wire N__20791;
    wire N__20788;
    wire N__20785;
    wire N__20782;
    wire N__20777;
    wire N__20774;
    wire N__20773;
    wire N__20770;
    wire N__20767;
    wire N__20764;
    wire N__20759;
    wire N__20756;
    wire N__20753;
    wire N__20752;
    wire N__20749;
    wire N__20746;
    wire N__20743;
    wire N__20738;
    wire N__20735;
    wire N__20732;
    wire N__20729;
    wire N__20728;
    wire N__20725;
    wire N__20722;
    wire N__20719;
    wire N__20716;
    wire N__20713;
    wire N__20712;
    wire N__20709;
    wire N__20706;
    wire N__20703;
    wire N__20696;
    wire N__20693;
    wire N__20690;
    wire N__20689;
    wire N__20686;
    wire N__20683;
    wire N__20680;
    wire N__20677;
    wire N__20674;
    wire N__20669;
    wire N__20668;
    wire N__20665;
    wire N__20662;
    wire N__20659;
    wire N__20656;
    wire N__20653;
    wire N__20648;
    wire N__20645;
    wire N__20642;
    wire N__20639;
    wire N__20636;
    wire N__20633;
    wire N__20630;
    wire N__20627;
    wire N__20624;
    wire N__20621;
    wire N__20618;
    wire N__20615;
    wire N__20612;
    wire N__20611;
    wire N__20608;
    wire N__20605;
    wire N__20600;
    wire N__20599;
    wire N__20596;
    wire N__20593;
    wire N__20590;
    wire N__20587;
    wire N__20584;
    wire N__20579;
    wire N__20576;
    wire N__20573;
    wire N__20570;
    wire N__20567;
    wire N__20566;
    wire N__20563;
    wire N__20560;
    wire N__20557;
    wire N__20556;
    wire N__20553;
    wire N__20550;
    wire N__20547;
    wire N__20544;
    wire N__20537;
    wire N__20534;
    wire N__20531;
    wire N__20528;
    wire N__20527;
    wire N__20524;
    wire N__20523;
    wire N__20520;
    wire N__20517;
    wire N__20514;
    wire N__20513;
    wire N__20510;
    wire N__20507;
    wire N__20502;
    wire N__20499;
    wire N__20492;
    wire N__20491;
    wire N__20486;
    wire N__20483;
    wire N__20482;
    wire N__20481;
    wire N__20478;
    wire N__20475;
    wire N__20472;
    wire N__20467;
    wire N__20462;
    wire N__20461;
    wire N__20458;
    wire N__20455;
    wire N__20452;
    wire N__20449;
    wire N__20446;
    wire N__20441;
    wire N__20438;
    wire N__20437;
    wire N__20434;
    wire N__20431;
    wire N__20428;
    wire N__20427;
    wire N__20426;
    wire N__20425;
    wire N__20424;
    wire N__20419;
    wire N__20414;
    wire N__20409;
    wire N__20402;
    wire N__20401;
    wire N__20398;
    wire N__20395;
    wire N__20392;
    wire N__20389;
    wire N__20386;
    wire N__20381;
    wire N__20380;
    wire N__20377;
    wire N__20376;
    wire N__20375;
    wire N__20372;
    wire N__20369;
    wire N__20366;
    wire N__20363;
    wire N__20360;
    wire N__20355;
    wire N__20350;
    wire N__20345;
    wire N__20342;
    wire N__20341;
    wire N__20338;
    wire N__20335;
    wire N__20332;
    wire N__20327;
    wire N__20324;
    wire N__20321;
    wire N__20318;
    wire N__20315;
    wire N__20312;
    wire N__20309;
    wire N__20306;
    wire N__20305;
    wire N__20302;
    wire N__20299;
    wire N__20296;
    wire N__20291;
    wire N__20290;
    wire N__20289;
    wire N__20286;
    wire N__20281;
    wire N__20276;
    wire N__20275;
    wire N__20274;
    wire N__20273;
    wire N__20270;
    wire N__20267;
    wire N__20266;
    wire N__20265;
    wire N__20262;
    wire N__20261;
    wire N__20254;
    wire N__20247;
    wire N__20244;
    wire N__20237;
    wire N__20234;
    wire N__20231;
    wire N__20228;
    wire N__20225;
    wire N__20222;
    wire N__20219;
    wire N__20216;
    wire N__20213;
    wire N__20210;
    wire N__20207;
    wire N__20204;
    wire N__20201;
    wire N__20198;
    wire N__20195;
    wire N__20192;
    wire N__20189;
    wire N__20186;
    wire N__20183;
    wire N__20182;
    wire N__20179;
    wire N__20178;
    wire N__20175;
    wire N__20172;
    wire N__20169;
    wire N__20166;
    wire N__20159;
    wire N__20156;
    wire N__20153;
    wire N__20150;
    wire N__20147;
    wire N__20144;
    wire N__20143;
    wire N__20140;
    wire N__20137;
    wire N__20136;
    wire N__20135;
    wire N__20132;
    wire N__20129;
    wire N__20126;
    wire N__20123;
    wire N__20122;
    wire N__20115;
    wire N__20112;
    wire N__20109;
    wire N__20104;
    wire N__20099;
    wire N__20098;
    wire N__20095;
    wire N__20094;
    wire N__20093;
    wire N__20090;
    wire N__20087;
    wire N__20082;
    wire N__20075;
    wire N__20074;
    wire N__20073;
    wire N__20072;
    wire N__20071;
    wire N__20068;
    wire N__20065;
    wire N__20062;
    wire N__20057;
    wire N__20054;
    wire N__20051;
    wire N__20048;
    wire N__20045;
    wire N__20036;
    wire N__20033;
    wire N__20030;
    wire N__20027;
    wire N__20024;
    wire N__20021;
    wire N__20018;
    wire N__20015;
    wire N__20012;
    wire N__20009;
    wire N__20006;
    wire N__20003;
    wire N__20000;
    wire N__19997;
    wire N__19996;
    wire N__19993;
    wire N__19990;
    wire N__19987;
    wire N__19984;
    wire N__19981;
    wire N__19978;
    wire N__19975;
    wire N__19972;
    wire N__19967;
    wire N__19964;
    wire N__19963;
    wire N__19960;
    wire N__19959;
    wire N__19958;
    wire N__19955;
    wire N__19952;
    wire N__19947;
    wire N__19940;
    wire N__19937;
    wire N__19936;
    wire N__19933;
    wire N__19930;
    wire N__19925;
    wire N__19922;
    wire N__19919;
    wire N__19918;
    wire N__19915;
    wire N__19912;
    wire N__19909;
    wire N__19904;
    wire N__19903;
    wire N__19902;
    wire N__19899;
    wire N__19898;
    wire N__19893;
    wire N__19888;
    wire N__19885;
    wire N__19880;
    wire N__19877;
    wire N__19874;
    wire N__19871;
    wire N__19868;
    wire N__19865;
    wire N__19862;
    wire N__19859;
    wire N__19858;
    wire N__19855;
    wire N__19852;
    wire N__19851;
    wire N__19848;
    wire N__19845;
    wire N__19842;
    wire N__19839;
    wire N__19832;
    wire N__19829;
    wire N__19826;
    wire N__19823;
    wire N__19822;
    wire N__19817;
    wire N__19814;
    wire N__19811;
    wire N__19808;
    wire N__19807;
    wire N__19804;
    wire N__19801;
    wire N__19796;
    wire N__19793;
    wire N__19790;
    wire N__19787;
    wire N__19784;
    wire N__19781;
    wire N__19778;
    wire N__19775;
    wire N__19772;
    wire N__19769;
    wire N__19766;
    wire N__19763;
    wire N__19760;
    wire N__19757;
    wire N__19754;
    wire N__19753;
    wire N__19750;
    wire N__19749;
    wire N__19748;
    wire N__19745;
    wire N__19742;
    wire N__19737;
    wire N__19730;
    wire N__19729;
    wire N__19726;
    wire N__19721;
    wire N__19718;
    wire N__19717;
    wire N__19714;
    wire N__19711;
    wire N__19708;
    wire N__19703;
    wire N__19700;
    wire N__19697;
    wire N__19694;
    wire N__19691;
    wire N__19688;
    wire N__19687;
    wire N__19684;
    wire N__19681;
    wire N__19678;
    wire N__19673;
    wire N__19670;
    wire N__19667;
    wire N__19664;
    wire N__19663;
    wire N__19660;
    wire N__19657;
    wire N__19654;
    wire N__19649;
    wire N__19646;
    wire N__19643;
    wire N__19640;
    wire N__19637;
    wire N__19636;
    wire N__19633;
    wire N__19630;
    wire N__19627;
    wire N__19622;
    wire N__19619;
    wire N__19616;
    wire N__19613;
    wire N__19610;
    wire N__19607;
    wire N__19604;
    wire N__19601;
    wire N__19598;
    wire N__19595;
    wire N__19592;
    wire N__19589;
    wire N__19586;
    wire N__19583;
    wire N__19580;
    wire N__19577;
    wire N__19574;
    wire N__19571;
    wire N__19568;
    wire N__19565;
    wire N__19562;
    wire N__19559;
    wire N__19556;
    wire N__19555;
    wire N__19552;
    wire N__19549;
    wire N__19544;
    wire N__19541;
    wire N__19540;
    wire N__19537;
    wire N__19534;
    wire N__19531;
    wire N__19526;
    wire N__19523;
    wire N__19520;
    wire N__19517;
    wire N__19514;
    wire N__19511;
    wire N__19508;
    wire N__19505;
    wire N__19502;
    wire N__19499;
    wire N__19496;
    wire N__19493;
    wire N__19490;
    wire N__19487;
    wire N__19484;
    wire N__19481;
    wire N__19478;
    wire N__19475;
    wire N__19474;
    wire N__19471;
    wire N__19468;
    wire N__19465;
    wire N__19460;
    wire N__19457;
    wire N__19454;
    wire N__19451;
    wire N__19448;
    wire N__19445;
    wire N__19444;
    wire N__19441;
    wire N__19438;
    wire N__19435;
    wire N__19430;
    wire N__19429;
    wire N__19426;
    wire N__19423;
    wire N__19420;
    wire N__19415;
    wire N__19414;
    wire N__19409;
    wire N__19406;
    wire N__19403;
    wire N__19402;
    wire N__19399;
    wire N__19396;
    wire N__19393;
    wire N__19388;
    wire N__19387;
    wire N__19384;
    wire N__19381;
    wire N__19376;
    wire N__19373;
    wire N__19372;
    wire N__19369;
    wire N__19366;
    wire N__19363;
    wire N__19358;
    wire N__19355;
    wire N__19352;
    wire N__19349;
    wire N__19346;
    wire N__19343;
    wire N__19340;
    wire N__19337;
    wire N__19334;
    wire N__19331;
    wire N__19328;
    wire N__19325;
    wire N__19324;
    wire N__19321;
    wire N__19318;
    wire N__19315;
    wire N__19310;
    wire N__19309;
    wire N__19306;
    wire N__19303;
    wire N__19300;
    wire N__19295;
    wire N__19292;
    wire N__19291;
    wire N__19288;
    wire N__19285;
    wire N__19282;
    wire N__19277;
    wire N__19276;
    wire N__19271;
    wire N__19268;
    wire N__19267;
    wire N__19264;
    wire N__19261;
    wire N__19258;
    wire N__19253;
    wire N__19252;
    wire N__19249;
    wire N__19244;
    wire N__19241;
    wire N__19238;
    wire N__19235;
    wire N__19232;
    wire N__19229;
    wire N__19228;
    wire N__19225;
    wire N__19222;
    wire N__19219;
    wire N__19216;
    wire N__19213;
    wire N__19208;
    wire N__19207;
    wire N__19204;
    wire N__19201;
    wire N__19198;
    wire N__19193;
    wire N__19192;
    wire N__19189;
    wire N__19186;
    wire N__19181;
    wire N__19178;
    wire N__19175;
    wire N__19174;
    wire N__19171;
    wire N__19168;
    wire N__19165;
    wire N__19160;
    wire N__19157;
    wire N__19154;
    wire N__19153;
    wire N__19150;
    wire N__19147;
    wire N__19144;
    wire N__19139;
    wire N__19136;
    wire N__19135;
    wire N__19132;
    wire N__19129;
    wire N__19126;
    wire N__19121;
    wire N__19118;
    wire N__19117;
    wire N__19114;
    wire N__19111;
    wire N__19108;
    wire N__19103;
    wire N__19100;
    wire N__19097;
    wire N__19096;
    wire N__19093;
    wire N__19090;
    wire N__19087;
    wire N__19082;
    wire N__19079;
    wire N__19078;
    wire N__19075;
    wire N__19072;
    wire N__19069;
    wire N__19064;
    wire N__19061;
    wire N__19058;
    wire N__19057;
    wire N__19054;
    wire N__19053;
    wire N__19050;
    wire N__19047;
    wire N__19044;
    wire N__19041;
    wire N__19038;
    wire N__19031;
    wire N__19028;
    wire N__19025;
    wire N__19022;
    wire N__19019;
    wire N__19016;
    wire N__19013;
    wire N__19012;
    wire N__19009;
    wire N__19006;
    wire N__19003;
    wire N__18998;
    wire N__18995;
    wire N__18994;
    wire N__18991;
    wire N__18988;
    wire N__18985;
    wire N__18980;
    wire N__18977;
    wire N__18974;
    wire N__18971;
    wire N__18968;
    wire N__18965;
    wire N__18962;
    wire N__18959;
    wire N__18956;
    wire N__18953;
    wire N__18950;
    wire N__18947;
    wire N__18944;
    wire N__18941;
    wire N__18938;
    wire N__18937;
    wire N__18936;
    wire N__18933;
    wire N__18930;
    wire N__18927;
    wire N__18924;
    wire N__18919;
    wire N__18916;
    wire N__18911;
    wire N__18908;
    wire N__18907;
    wire N__18904;
    wire N__18903;
    wire N__18900;
    wire N__18897;
    wire N__18894;
    wire N__18891;
    wire N__18884;
    wire N__18883;
    wire N__18880;
    wire N__18877;
    wire N__18876;
    wire N__18873;
    wire N__18868;
    wire N__18863;
    wire N__18862;
    wire N__18859;
    wire N__18856;
    wire N__18855;
    wire N__18850;
    wire N__18847;
    wire N__18842;
    wire N__18839;
    wire N__18836;
    wire N__18833;
    wire N__18830;
    wire N__18827;
    wire N__18824;
    wire N__18821;
    wire N__18818;
    wire N__18815;
    wire N__18812;
    wire N__18809;
    wire N__18806;
    wire N__18803;
    wire N__18800;
    wire N__18797;
    wire N__18794;
    wire N__18793;
    wire N__18790;
    wire N__18789;
    wire N__18786;
    wire N__18783;
    wire N__18780;
    wire N__18773;
    wire N__18770;
    wire N__18769;
    wire N__18768;
    wire N__18767;
    wire N__18764;
    wire N__18761;
    wire N__18758;
    wire N__18755;
    wire N__18750;
    wire N__18743;
    wire N__18740;
    wire N__18739;
    wire N__18736;
    wire N__18735;
    wire N__18732;
    wire N__18731;
    wire N__18728;
    wire N__18725;
    wire N__18722;
    wire N__18719;
    wire N__18714;
    wire N__18707;
    wire N__18706;
    wire N__18705;
    wire N__18700;
    wire N__18697;
    wire N__18694;
    wire N__18689;
    wire N__18686;
    wire N__18683;
    wire N__18680;
    wire N__18679;
    wire N__18678;
    wire N__18675;
    wire N__18672;
    wire N__18669;
    wire N__18662;
    wire N__18659;
    wire N__18658;
    wire N__18657;
    wire N__18654;
    wire N__18649;
    wire N__18644;
    wire N__18641;
    wire N__18640;
    wire N__18639;
    wire N__18638;
    wire N__18635;
    wire N__18632;
    wire N__18629;
    wire N__18626;
    wire N__18617;
    wire N__18614;
    wire N__18611;
    wire N__18608;
    wire N__18605;
    wire N__18604;
    wire N__18603;
    wire N__18600;
    wire N__18595;
    wire N__18590;
    wire N__18589;
    wire N__18588;
    wire N__18585;
    wire N__18582;
    wire N__18579;
    wire N__18572;
    wire N__18571;
    wire N__18570;
    wire N__18567;
    wire N__18564;
    wire N__18559;
    wire N__18554;
    wire N__18553;
    wire N__18552;
    wire N__18549;
    wire N__18544;
    wire N__18539;
    wire N__18538;
    wire N__18537;
    wire N__18534;
    wire N__18531;
    wire N__18528;
    wire N__18521;
    wire N__18518;
    wire N__18517;
    wire N__18516;
    wire N__18513;
    wire N__18510;
    wire N__18507;
    wire N__18500;
    wire N__18499;
    wire N__18498;
    wire N__18495;
    wire N__18492;
    wire N__18489;
    wire N__18482;
    wire N__18479;
    wire N__18478;
    wire N__18477;
    wire N__18474;
    wire N__18469;
    wire N__18466;
    wire N__18461;
    wire N__18458;
    wire N__18455;
    wire N__18452;
    wire N__18449;
    wire N__18446;
    wire N__18445;
    wire N__18444;
    wire N__18443;
    wire N__18442;
    wire N__18441;
    wire N__18440;
    wire N__18439;
    wire N__18438;
    wire N__18435;
    wire N__18432;
    wire N__18423;
    wire N__18420;
    wire N__18417;
    wire N__18414;
    wire N__18401;
    wire N__18398;
    wire N__18397;
    wire N__18396;
    wire N__18393;
    wire N__18390;
    wire N__18387;
    wire N__18380;
    wire N__18377;
    wire N__18376;
    wire N__18373;
    wire N__18370;
    wire N__18365;
    wire N__18362;
    wire N__18359;
    wire N__18356;
    wire N__18353;
    wire N__18350;
    wire N__18347;
    wire N__18344;
    wire N__18341;
    wire N__18338;
    wire N__18335;
    wire N__18332;
    wire N__18329;
    wire N__18326;
    wire N__18323;
    wire N__18320;
    wire N__18317;
    wire N__18314;
    wire N__18311;
    wire N__18310;
    wire N__18307;
    wire N__18304;
    wire N__18301;
    wire N__18296;
    wire N__18293;
    wire N__18290;
    wire N__18287;
    wire N__18284;
    wire N__18283;
    wire N__18280;
    wire N__18277;
    wire N__18274;
    wire N__18269;
    wire N__18266;
    wire N__18263;
    wire N__18262;
    wire N__18259;
    wire N__18256;
    wire N__18251;
    wire N__18250;
    wire N__18247;
    wire N__18244;
    wire N__18241;
    wire N__18236;
    wire N__18233;
    wire N__18230;
    wire N__18227;
    wire N__18226;
    wire N__18223;
    wire N__18220;
    wire N__18217;
    wire N__18212;
    wire N__18211;
    wire N__18208;
    wire N__18205;
    wire N__18200;
    wire N__18197;
    wire N__18194;
    wire N__18191;
    wire N__18188;
    wire N__18185;
    wire N__18182;
    wire N__18179;
    wire N__18176;
    wire N__18173;
    wire N__18170;
    wire N__18167;
    wire N__18164;
    wire N__18161;
    wire N__18158;
    wire N__18155;
    wire N__18152;
    wire N__18149;
    wire N__18148;
    wire N__18145;
    wire N__18142;
    wire N__18139;
    wire N__18134;
    wire N__18131;
    wire N__18128;
    wire N__18125;
    wire N__18122;
    wire N__18121;
    wire N__18118;
    wire N__18115;
    wire N__18112;
    wire N__18107;
    wire N__18104;
    wire N__18101;
    wire N__18098;
    wire N__18095;
    wire N__18092;
    wire N__18089;
    wire N__18086;
    wire N__18083;
    wire N__18080;
    wire N__18079;
    wire N__18076;
    wire N__18073;
    wire N__18068;
    wire N__18065;
    wire N__18064;
    wire N__18061;
    wire N__18058;
    wire N__18055;
    wire N__18050;
    wire N__18047;
    wire N__18046;
    wire N__18043;
    wire N__18040;
    wire N__18037;
    wire N__18032;
    wire N__18029;
    wire N__18026;
    wire N__18025;
    wire N__18022;
    wire N__18017;
    wire N__18014;
    wire N__18011;
    wire N__18008;
    wire N__18005;
    wire N__18002;
    wire N__17999;
    wire N__17998;
    wire N__17995;
    wire N__17992;
    wire N__17989;
    wire N__17984;
    wire N__17981;
    wire N__17978;
    wire N__17977;
    wire N__17974;
    wire N__17971;
    wire N__17968;
    wire N__17963;
    wire N__17962;
    wire N__17959;
    wire N__17956;
    wire N__17951;
    wire N__17950;
    wire N__17947;
    wire N__17944;
    wire N__17939;
    wire N__17938;
    wire N__17935;
    wire N__17932;
    wire N__17927;
    wire N__17924;
    wire N__17921;
    wire N__17920;
    wire N__17917;
    wire N__17914;
    wire N__17911;
    wire N__17906;
    wire N__17905;
    wire N__17902;
    wire N__17899;
    wire N__17894;
    wire N__17893;
    wire N__17890;
    wire N__17887;
    wire N__17884;
    wire N__17879;
    wire N__17876;
    wire N__17875;
    wire N__17872;
    wire N__17869;
    wire N__17866;
    wire N__17861;
    wire N__17860;
    wire N__17857;
    wire N__17854;
    wire N__17851;
    wire N__17846;
    wire N__17843;
    wire N__17842;
    wire N__17839;
    wire N__17836;
    wire N__17833;
    wire N__17828;
    wire N__17825;
    wire N__17824;
    wire N__17821;
    wire N__17818;
    wire N__17815;
    wire N__17810;
    wire N__17807;
    wire N__17806;
    wire N__17803;
    wire N__17800;
    wire N__17797;
    wire N__17792;
    wire N__17789;
    wire N__17788;
    wire N__17783;
    wire N__17780;
    wire N__17777;
    wire N__17774;
    wire N__17771;
    wire N__17768;
    wire N__17765;
    wire N__17762;
    wire N__17759;
    wire N__17758;
    wire N__17753;
    wire N__17750;
    wire N__17747;
    wire N__17744;
    wire N__17743;
    wire N__17740;
    wire N__17737;
    wire N__17734;
    wire N__17729;
    wire N__17726;
    wire N__17725;
    wire N__17722;
    wire N__17719;
    wire N__17716;
    wire N__17711;
    wire N__17708;
    wire N__17705;
    wire N__17704;
    wire N__17701;
    wire N__17698;
    wire N__17695;
    wire N__17690;
    wire N__17687;
    wire N__17684;
    wire N__17681;
    wire N__17680;
    wire N__17677;
    wire N__17674;
    wire N__17671;
    wire N__17666;
    wire N__17663;
    wire N__17660;
    wire N__17657;
    wire N__17654;
    wire N__17651;
    wire N__17648;
    wire N__17645;
    wire N__17642;
    wire N__17639;
    wire N__17636;
    wire N__17633;
    wire N__17630;
    wire N__17627;
    wire N__17624;
    wire N__17621;
    wire N__17618;
    wire N__17615;
    wire N__17614;
    wire N__17611;
    wire N__17608;
    wire N__17603;
    wire N__17600;
    wire N__17597;
    wire N__17594;
    wire N__17591;
    wire N__17588;
    wire N__17585;
    wire N__17582;
    wire N__17579;
    wire N__17578;
    wire N__17577;
    wire N__17576;
    wire N__17569;
    wire N__17566;
    wire N__17563;
    wire N__17558;
    wire N__17555;
    wire N__17552;
    wire N__17549;
    wire N__17548;
    wire N__17545;
    wire N__17542;
    wire N__17537;
    wire N__17536;
    wire N__17533;
    wire N__17530;
    wire N__17527;
    wire N__17524;
    wire N__17519;
    wire N__17516;
    wire N__17513;
    wire N__17510;
    wire N__17507;
    wire N__17504;
    wire N__17501;
    wire N__17500;
    wire N__17499;
    wire N__17498;
    wire N__17495;
    wire N__17494;
    wire N__17489;
    wire N__17486;
    wire N__17483;
    wire N__17480;
    wire N__17471;
    wire N__17470;
    wire N__17467;
    wire N__17464;
    wire N__17459;
    wire N__17456;
    wire N__17453;
    wire N__17452;
    wire N__17451;
    wire N__17448;
    wire N__17443;
    wire N__17438;
    wire N__17435;
    wire N__17432;
    wire N__17429;
    wire N__17426;
    wire N__17423;
    wire N__17420;
    wire N__17417;
    wire N__17414;
    wire N__17411;
    wire N__17408;
    wire N__17405;
    wire N__17402;
    wire N__17399;
    wire N__17396;
    wire N__17393;
    wire N__17392;
    wire N__17391;
    wire N__17390;
    wire N__17385;
    wire N__17382;
    wire N__17379;
    wire N__17372;
    wire N__17369;
    wire N__17366;
    wire N__17363;
    wire N__17360;
    wire N__17357;
    wire N__17354;
    wire N__17351;
    wire N__17348;
    wire N__17345;
    wire N__17342;
    wire N__17339;
    wire N__17336;
    wire N__17333;
    wire N__17330;
    wire N__17327;
    wire N__17324;
    wire N__17321;
    wire N__17318;
    wire N__17315;
    wire N__17312;
    wire N__17309;
    wire N__17306;
    wire N__17303;
    wire N__17300;
    wire N__17297;
    wire N__17294;
    wire N__17291;
    wire N__17288;
    wire N__17285;
    wire N__17282;
    wire N__17281;
    wire N__17276;
    wire N__17273;
    wire N__17270;
    wire N__17267;
    wire N__17264;
    wire N__17261;
    wire N__17258;
    wire N__17255;
    wire N__17252;
    wire N__17249;
    wire N__17246;
    wire N__17245;
    wire N__17242;
    wire N__17239;
    wire N__17236;
    wire N__17231;
    wire N__17228;
    wire N__17225;
    wire N__17222;
    wire N__17219;
    wire N__17216;
    wire N__17213;
    wire N__17210;
    wire N__17207;
    wire N__17204;
    wire N__17201;
    wire N__17198;
    wire N__17197;
    wire N__17194;
    wire N__17191;
    wire N__17188;
    wire N__17183;
    wire N__17180;
    wire N__17177;
    wire N__17174;
    wire N__17171;
    wire N__17170;
    wire N__17167;
    wire N__17164;
    wire N__17159;
    wire N__17158;
    wire N__17155;
    wire N__17152;
    wire N__17149;
    wire N__17144;
    wire N__17141;
    wire N__17140;
    wire N__17137;
    wire N__17134;
    wire N__17131;
    wire N__17126;
    wire N__17123;
    wire N__17120;
    wire N__17117;
    wire N__17116;
    wire N__17113;
    wire N__17110;
    wire N__17105;
    wire N__17102;
    wire N__17099;
    wire N__17096;
    wire N__17093;
    wire N__17090;
    wire N__17087;
    wire N__17084;
    wire N__17081;
    wire N__17078;
    wire N__17077;
    wire N__17072;
    wire N__17069;
    wire N__17068;
    wire N__17063;
    wire N__17060;
    wire N__17059;
    wire N__17056;
    wire N__17053;
    wire N__17050;
    wire N__17045;
    wire N__17042;
    wire N__17041;
    wire N__17038;
    wire N__17033;
    wire N__17030;
    wire N__17027;
    wire N__17024;
    wire N__17021;
    wire N__17018;
    wire N__17015;
    wire N__17012;
    wire N__17009;
    wire N__17006;
    wire N__17003;
    wire N__17002;
    wire N__16999;
    wire N__16996;
    wire N__16991;
    wire N__16988;
    wire N__16985;
    wire N__16982;
    wire N__16979;
    wire N__16976;
    wire N__16973;
    wire N__16970;
    wire N__16967;
    wire N__16964;
    wire N__16961;
    wire N__16958;
    wire N__16955;
    wire N__16952;
    wire N__16949;
    wire N__16946;
    wire N__16945;
    wire N__16942;
    wire N__16941;
    wire N__16938;
    wire N__16937;
    wire N__16928;
    wire N__16925;
    wire N__16922;
    wire N__16919;
    wire N__16916;
    wire N__16913;
    wire N__16910;
    wire CLK_pad_gb_input;
    wire VCCG0;
    wire GNDG0;
    wire \c0.data_in_frame_0_3 ;
    wire \c0.n9186_cascade_ ;
    wire \c0.n8857_cascade_ ;
    wire \c0.n8725_cascade_ ;
    wire \c0.n8063_cascade_ ;
    wire \c0.n20_adj_2547_cascade_ ;
    wire \c0.n9317 ;
    wire \c0.n8063 ;
    wire \c0.n17650 ;
    wire \c0.n8645_cascade_ ;
    wire \c0.n9186 ;
    wire \c0.n30_adj_2489_cascade_ ;
    wire \c0.n18_adj_2545 ;
    wire bfn_1_22_0_;
    wire \c0.n16405 ;
    wire \c0.n16406 ;
    wire \c0.n16407 ;
    wire \c0.n16408 ;
    wire \c0.n16409 ;
    wire \c0.n16410 ;
    wire \c0.n16411 ;
    wire \c0.data_out_frame2_0_0 ;
    wire data_out_frame2_7_2;
    wire \c0.data_out_frame2_0_6 ;
    wire \c0.n18546_cascade_ ;
    wire data_out_frame2_11_5;
    wire \c0.n18474 ;
    wire \c0.n18534_cascade_ ;
    wire data_out_frame2_17_5;
    wire \c0.n18537_cascade_ ;
    wire \c0.n17803 ;
    wire \c0.n18080 ;
    wire \c0.n18384_cascade_ ;
    wire \c0.n22_adj_2523 ;
    wire \c0.n18387_cascade_ ;
    wire \c0.n5_adj_2463 ;
    wire data_out_frame2_16_5;
    wire data_out_frame2_9_5;
    wire data_out_frame2_6_2;
    wire data_out_frame2_16_2;
    wire \c0.n18486_cascade_ ;
    wire \c0.n18489_cascade_ ;
    wire \c0.n18084 ;
    wire \c0.n18366_cascade_ ;
    wire \c0.n6_adj_2466 ;
    wire \c0.n22_adj_2529 ;
    wire \c0.n18369_cascade_ ;
    wire data_out_frame2_7_5;
    wire \c0.n5_adj_2503_cascade_ ;
    wire data_out_frame2_14_2;
    wire \c0.n18606_cascade_ ;
    wire \c0.n18570_cascade_ ;
    wire \c0.n17779 ;
    wire \c0.n17773_cascade_ ;
    wire \c0.n18074 ;
    wire \c0.n18432_cascade_ ;
    wire \c0.n18435_cascade_ ;
    wire \c0.n17836 ;
    wire \c0.n18360_cascade_ ;
    wire \c0.n6_adj_2504 ;
    wire \c0.n18471_cascade_ ;
    wire \c0.n18363 ;
    wire \c0.n22_adj_2530_cascade_ ;
    wire bfn_1_31_0_;
    wire \c0.tx2.n16372 ;
    wire \c0.tx2.n16373 ;
    wire \c0.tx2.n16374 ;
    wire \c0.tx2.n16375 ;
    wire \c0.tx2.n16376 ;
    wire \c0.tx2.n16377 ;
    wire \c0.tx2.n16378 ;
    wire \c0.tx2.n16379 ;
    wire bfn_1_32_0_;
    wire \c0.tx2.n17953 ;
    wire \c0.tx2.n18013 ;
    wire \c0.tx2.n17939 ;
    wire n316;
    wire \c0.n17507_cascade_ ;
    wire \c0.data_in_frame_0_4 ;
    wire \c0.n17507 ;
    wire \c0.n17476_cascade_ ;
    wire \c0.n17476 ;
    wire \c0.n17478_cascade_ ;
    wire \c0.n17629_cascade_ ;
    wire \c0.n16_adj_2546 ;
    wire \c0.n9254 ;
    wire \c0.n9254_cascade_ ;
    wire \c0.data_in_frame_2_5 ;
    wire \c0.n8976 ;
    wire \c0.data_in_frame_1_3 ;
    wire \c0.n5_adj_2515 ;
    wire \c0.data_out_frame2_0_5 ;
    wire \c0.data_in_frame_3_3 ;
    wire \c0.n2607 ;
    wire \c0.n17513 ;
    wire \c0.n2602 ;
    wire \c0.data_in_frame_3_2 ;
    wire \c0.n9_adj_2500 ;
    wire \c0.n9_adj_2507 ;
    wire \c0.n17325_cascade_ ;
    wire \c0.n8_adj_2459_cascade_ ;
    wire \c0.n2604 ;
    wire \c0.n11_adj_2460 ;
    wire \c0.n9605 ;
    wire \c0.n9900 ;
    wire \c0.n17806 ;
    wire data_out_frame2_18_5;
    wire data_out_frame2_13_2;
    wire \c0.n18492 ;
    wire \c0.n17827 ;
    wire data_out_frame2_12_5;
    wire \c0.n9043_cascade_ ;
    wire data_out_frame2_14_6;
    wire data_out_frame2_10_6;
    wire data_out_frame2_11_0;
    wire data_out_frame2_6_6;
    wire data_out_frame2_7_6;
    wire data_out_frame2_8_5;
    wire data_out_frame2_15_1;
    wire data_out_frame2_11_6;
    wire data_out_frame2_15_6;
    wire data_out_frame2_5_2;
    wire data_out_frame2_15_2;
    wire data_out_frame2_15_0;
    wire data_out_frame2_8_6;
    wire \c0.n18564 ;
    wire data_out_frame2_16_1;
    wire data_out_frame2_17_1;
    wire data_out_frame2_18_0;
    wire data_out_frame2_10_3;
    wire data_out_frame2_14_4;
    wire \c0.n5_adj_2495 ;
    wire data_out_frame2_5_5;
    wire \c0.n6_adj_2496 ;
    wire data_out_frame2_11_3;
    wire \c0.n17629 ;
    wire \c0.n8725 ;
    wire data_out_frame2_10_0;
    wire data_out_frame2_17_0;
    wire data_out_frame2_16_0;
    wire \c0.n18600 ;
    wire data_out_frame2_5_0;
    wire \c0.n5_adj_2477_cascade_ ;
    wire \c0.n6_adj_2436 ;
    wire data_out_frame2_18_1;
    wire \c0.n18468 ;
    wire data_out_frame2_5_1;
    wire data_out_frame2_10_2;
    wire data_out_frame2_11_2;
    wire data_out_frame2_12_0;
    wire \c0.n17794 ;
    wire \c0.n18078 ;
    wire \c0.n18408_cascade_ ;
    wire \c0.n6_adj_2506 ;
    wire \c0.n18411_cascade_ ;
    wire data_out_frame2_18_6;
    wire \c0.n18552_cascade_ ;
    wire \c0.n18555_cascade_ ;
    wire \c0.n22_adj_2521 ;
    wire n317;
    wire n318;
    wire n319;
    wire n321;
    wire r_Clock_Count_0_adj_2634;
    wire r_Clock_Count_2_adj_2632;
    wire r_Clock_Count_4_adj_2630;
    wire r_Clock_Count_3_adj_2631;
    wire r_Clock_Count_5_adj_2629;
    wire \c0.tx2.n10_cascade_ ;
    wire \c0.tx2.r_Clock_Count_7 ;
    wire \c0.tx2.r_Clock_Count_6 ;
    wire \c0.tx2.r_Clock_Count_8 ;
    wire \c0.tx2.n16452 ;
    wire \c0.tx2.r_SM_Main_2_N_2323_1_cascade_ ;
    wire n320;
    wire n10244;
    wire r_Clock_Count_1_adj_2633;
    wire \c0.tx2.o_Tx_Serial_N_2354 ;
    wire \c0.tx2.n12306_cascade_ ;
    wire \c0.n12_adj_2492 ;
    wire \c0.data_in_frame_0_7 ;
    wire \c0.data_in_frame_2_0 ;
    wire \c0.n17553_cascade_ ;
    wire \c0.data_in_frame_3_7 ;
    wire \c0.n17406_cascade_ ;
    wire data_in_frame_5_5;
    wire \c0.data_in_frame_2_4 ;
    wire \c0.data_in_frame_1_5 ;
    wire n9419_cascade_;
    wire \c0.n25_adj_2491 ;
    wire n1396_cascade_;
    wire n2589_cascade_;
    wire n2589;
    wire \c0.n18558 ;
    wire \c0.n17797 ;
    wire \c0.n17424 ;
    wire \c0.n17569 ;
    wire \c0.n10_adj_2505 ;
    wire \c0.n9028 ;
    wire \c0.n8061_cascade_ ;
    wire \c0.data_in_frame_6_4 ;
    wire n2595;
    wire \c0.data_in_frame_0_0 ;
    wire \c0.n2839 ;
    wire \c0.n9151_cascade_ ;
    wire \c0.n17588_cascade_ ;
    wire data_in_frame_8_5;
    wire \c0.n6_adj_2429 ;
    wire \c0.data_out_frame2_20_5 ;
    wire data_out_frame2_12_2;
    wire data_out_frame2_13_1;
    wire data_out_frame2_12_1;
    wire data_out_frame2_7_0;
    wire n9606_cascade_;
    wire data_out_frame2_10_5;
    wire data_out_frame2_13_5;
    wire data_out_frame2_9_0;
    wire data_out_frame2_6_1;
    wire data_out_frame2_17_2;
    wire data_out_frame2_5_7;
    wire data_out_frame2_6_5;
    wire data_out_frame2_6_0;
    wire data_out_frame2_7_1;
    wire data_out_frame2_16_6;
    wire data_out_frame2_11_7;
    wire data_out_frame2_9_1;
    wire data_out_frame2_8_1;
    wire \c0.n17833 ;
    wire data_out_frame2_19_0;
    wire \c0.n18603 ;
    wire \c0.n22_adj_2510 ;
    wire data_out_frame2_14_7;
    wire data_out_frame2_15_7;
    wire data_out_frame2_12_7;
    wire \c0.n18582_cascade_ ;
    wire data_out_frame2_13_7;
    wire data_out_frame2_9_2;
    wire data_out_frame2_8_2;
    wire \c0.n18504 ;
    wire \c0.n17824 ;
    wire \c0.tx2.r_Tx_Data_2 ;
    wire \c0.tx2.r_Tx_Data_0 ;
    wire \c0.tx2.r_Tx_Data_1 ;
    wire \c0.tx2.n18612_cascade_ ;
    wire \c0.tx2.n18615 ;
    wire \c0.tx2.r_Tx_Data_6 ;
    wire data_out_frame2_17_6;
    wire data_out_frame2_13_4;
    wire \c0.n12 ;
    wire \c0.n11_cascade_ ;
    wire \c0.tx2.r_Tx_Data_5 ;
    wire \c0.tx2.n18450 ;
    wire \c0.tx2.n18453 ;
    wire data_out_frame2_5_3;
    wire data_out_frame2_7_3;
    wire \c0.n5_adj_2509 ;
    wire \c0.byte_transmit_counter2_5 ;
    wire \c0.byte_transmit_counter2_6 ;
    wire \c0.n18_adj_2544_cascade_ ;
    wire \c0.byte_transmit_counter2_7 ;
    wire \c0.n19_adj_2540_cascade_ ;
    wire \c0.tx2_transmit_N_2287 ;
    wire \c0.tx2_transmit_N_2287_cascade_ ;
    wire \c0.n19_adj_2540 ;
    wire \c0.n67_cascade_ ;
    wire \c0.n13530 ;
    wire \c0.n17656 ;
    wire \c0.n20_adj_2427 ;
    wire \c0.n10_adj_2428_cascade_ ;
    wire \c0.n17442 ;
    wire \c0.n17553 ;
    wire \c0.n17442_cascade_ ;
    wire \c0.n17550 ;
    wire \c0.data_in_frame_4_0 ;
    wire \c0.n8874 ;
    wire \c0.data_in_frame_1_4 ;
    wire \c0.n8874_cascade_ ;
    wire \c0.n9349 ;
    wire \c0.n9368_cascade_ ;
    wire \c0.n23_adj_2426 ;
    wire \c0.data_in_frame_1_6 ;
    wire \c0.n17632 ;
    wire \c0.n17485 ;
    wire \c0.data_in_frame_3_1 ;
    wire \c0.n17406 ;
    wire \c0.n12_adj_2449_cascade_ ;
    wire n2598;
    wire \c0.n23_adj_2462 ;
    wire \c0.n24_adj_2454_cascade_ ;
    wire data_in_frame_5_3;
    wire \c0.data_in_frame_2_7 ;
    wire \c0.data_in_frame_7_7 ;
    wire n2584;
    wire \c0.n9151 ;
    wire n2584_cascade_;
    wire \c0.n21_adj_2465 ;
    wire n9419;
    wire \c0.n8061 ;
    wire \c0.n8857 ;
    wire \c0.n18_adj_2468 ;
    wire \c0.n26_adj_2469_cascade_ ;
    wire \c0.n30 ;
    wire data_out_frame2_6_7;
    wire \c0.n5_adj_2501 ;
    wire \c0.n17534 ;
    wire \c0.n8674 ;
    wire \c0.n9163 ;
    wire \c0.n17470 ;
    wire n9148;
    wire n9148_cascade_;
    wire \c0.n22_adj_2508 ;
    wire \c0.n12_adj_2542 ;
    wire \c0.data_in_frame_2_2 ;
    wire \c0.n9058 ;
    wire \c0.n17467 ;
    wire \c0.data_in_frame_4_3 ;
    wire \c0.n17562 ;
    wire data_in_frame_8_7;
    wire \c0.n17647_cascade_ ;
    wire \c0.n12_adj_2549 ;
    wire data_in_8_5;
    wire \c0.n17602 ;
    wire \c0.n30_adj_2489 ;
    wire \c0.n9345 ;
    wire \c0.n9345_cascade_ ;
    wire \c0.n10_cascade_ ;
    wire \c0.data_out_frame2_20_6 ;
    wire \c0.n17647 ;
    wire \c0.n8995 ;
    wire \c0.n6_adj_2550 ;
    wire \c0.data_out_frame2_20_0 ;
    wire \c0.n6_adj_2502_cascade_ ;
    wire \c0.data_out_frame2_20_2 ;
    wire \c0.data_out_frame2_19_5 ;
    wire data_out_frame2_14_0;
    wire data_out_frame2_18_2;
    wire data_out_frame2_5_6;
    wire data_out_frame2_6_3;
    wire data_out_frame2_12_6;
    wire data_out_frame2_13_6;
    wire data_out_frame2_8_0;
    wire data_out_frame2_10_7;
    wire data_out_frame2_15_4;
    wire data_out_frame2_12_4;
    wire \c0.n17535_cascade_ ;
    wire \c0.data_out_frame2_19_6 ;
    wire \c0.n9240 ;
    wire \c0.n9240_cascade_ ;
    wire \c0.n9131 ;
    wire \c0.n17409_cascade_ ;
    wire \c0.n10_adj_2470 ;
    wire \c0.data_out_frame2_20_1 ;
    wire \c0.data_out_frame2_19_1 ;
    wire \c0.n6_adj_2464 ;
    wire \c0.n18423_cascade_ ;
    wire \c0.tx2.r_Tx_Data_7 ;
    wire data_out_frame2_18_7;
    wire \c0.data_out_frame2_19_7 ;
    wire \c0.n18576_cascade_ ;
    wire data_out_frame2_17_7;
    wire \c0.n18579_cascade_ ;
    wire \c0.n22_adj_2520 ;
    wire \c0.n17788 ;
    wire \c0.n18420 ;
    wire \c0.n4_adj_2480 ;
    wire tx_enable;
    wire tx2_o;
    wire tx2_enable;
    wire \c0.tx2.n4 ;
    wire \c0.tx2.n9568_cascade_ ;
    wire \c0.tx2.tx2_active ;
    wire \c0.tx2.n23 ;
    wire \c0.r_SM_Main_2_N_2326_0 ;
    wire \c0.tx2.n17990 ;
    wire \c0.tx2.r_SM_Main_2_N_2323_1 ;
    wire \c0.tx2.n12_cascade_ ;
    wire r_SM_Main_2_adj_2628;
    wire \c0.tx2.r_SM_Main_0 ;
    wire \c0.tx2.r_SM_Main_1 ;
    wire \c0.tx2.n6812_cascade_ ;
    wire data_in_0_7;
    wire \c0.n17697_cascade_ ;
    wire data_in_0_4;
    wire data_in_frame_5_0;
    wire \c0.n9306 ;
    wire \c0.data_in_frame_1_2 ;
    wire \c0.data_in_frame_6_1 ;
    wire \c0.n9328 ;
    wire \c0.n8645 ;
    wire n9100;
    wire \c0.data_in_frame_4_5 ;
    wire \c0.data_in_frame_0_5 ;
    wire \c0.data_in_frame_4_4 ;
    wire \c0.n9176 ;
    wire \c0.data_in_frame_4_2 ;
    wire \c0.data_in_frame_2_3 ;
    wire \c0.n10_adj_2430_cascade_ ;
    wire \c0.data_in_frame_4_1 ;
    wire \c0.n8695_cascade_ ;
    wire \c0.n8867 ;
    wire \c0.data_in_frame_0_6 ;
    wire \c0.data_in_frame_3_4 ;
    wire data_in_5_0;
    wire data_in_7_6;
    wire n2593;
    wire n2593_cascade_;
    wire \c0.n22_adj_2461 ;
    wire n2586;
    wire \c0.n9279 ;
    wire n2590_cascade_;
    wire \c0.n10_adj_2450 ;
    wire data_in_6_3;
    wire n2596;
    wire \c0.n17529 ;
    wire n2596_cascade_;
    wire \c0.n10_adj_2498 ;
    wire \c0.data_in_frame_7_3 ;
    wire n2588;
    wire \c0.n8687 ;
    wire n2585;
    wire \c0.n17 ;
    wire n2590;
    wire \c0.data_in_frame_7_1 ;
    wire \c0.data_in_frame_1_0 ;
    wire \c0.data_in_frame_4_6 ;
    wire \c0.data_in_frame_3_0 ;
    wire \c0.data_in_frame_4_7 ;
    wire \c0.n17403 ;
    wire \c0.n17403_cascade_ ;
    wire \c0.data_in_frame_2_6 ;
    wire n9283;
    wire n9283_cascade_;
    wire data_out_frame2_16_7;
    wire \c0.n9219 ;
    wire \c0.n8695 ;
    wire \c0.data_in_frame_6_6 ;
    wire \c0.n9208 ;
    wire \c0.n22_cascade_ ;
    wire n16_adj_2656;
    wire \c0.n17519 ;
    wire \c0.n24_cascade_ ;
    wire \c0.n11_adj_2453 ;
    wire data_in_frame_8_2;
    wire data_in_frame_8_1;
    wire \c0.data_in_frame_6_3 ;
    wire \c0.n17605 ;
    wire \c0.n20 ;
    wire \c0.data_in_frame_7_6 ;
    wire \c0.n9144 ;
    wire \c0.n8064 ;
    wire \c0.n17582_cascade_ ;
    wire \c0.data_out_frame2_20_7 ;
    wire n2560;
    wire \c0.n17588 ;
    wire \c0.n17582 ;
    wire n2560_cascade_;
    wire n17585;
    wire \c0.n17648 ;
    wire \c0.n18_cascade_ ;
    wire \c0.n17418 ;
    wire n2572;
    wire bfn_5_25_0_;
    wire \c0.tx.n16357 ;
    wire \c0.tx.n16358 ;
    wire \c0.tx.n16359 ;
    wire \c0.tx.n16360 ;
    wire \c0.tx.n16361 ;
    wire \c0.tx.n16362 ;
    wire \c0.tx.n16363 ;
    wire \c0.tx.n16364 ;
    wire bfn_5_26_0_;
    wire \c0.n31 ;
    wire data_out_frame2_9_6;
    wire data_out_frame2_15_3;
    wire data_out_frame2_14_3;
    wire \c0.n18516_cascade_ ;
    wire data_out_frame2_13_3;
    wire data_out_frame2_11_1;
    wire data_out_frame2_10_1;
    wire \c0.n18480 ;
    wire \c0.n136 ;
    wire \c0.n1_adj_2443 ;
    wire \c0.n14631_cascade_ ;
    wire \c0.data_out_frame2_0_2 ;
    wire \c0.n17482 ;
    wire data_out_frame2_9_3;
    wire data_out_frame2_8_3;
    wire \c0.n18522 ;
    wire \c0.data_out_frame2_0_7 ;
    wire \c0.n18076 ;
    wire data_out_frame2_9_7;
    wire data_out_frame2_8_7;
    wire \c0.n18588 ;
    wire \c0.n17785 ;
    wire bfn_5_29_0_;
    wire n16319;
    wire n16320;
    wire n16321;
    wire n16322;
    wire n16323;
    wire n16324;
    wire n16325;
    wire n16326;
    wire bfn_5_30_0_;
    wire n16327;
    wire n16328;
    wire n16329;
    wire n16330;
    wire n16331;
    wire n16332;
    wire n16333;
    wire n16334;
    wire bfn_5_31_0_;
    wire n16335;
    wire n16336;
    wire n16337;
    wire n16338;
    wire n16339;
    wire n16340;
    wire n16341;
    wire n16342;
    wire bfn_5_32_0_;
    wire n16343;
    wire n16344;
    wire n16345;
    wire n16346;
    wire n16347;
    wire n16348;
    wire n16349;
    wire data_in_5_3;
    wire \c0.n17715_cascade_ ;
    wire data_out_frame2_15_5;
    wire \c0.n18540 ;
    wire \c0.data_in_1_0 ;
    wire \c0.data_in_0_0 ;
    wire data_in_3_7;
    wire \c0.n6_adj_2473 ;
    wire data_in_8_0;
    wire \c0.n81 ;
    wire data_in_6_0;
    wire \c0.data_in_frame_6_0 ;
    wire n2599;
    wire n2599_cascade_;
    wire \c0.n20_adj_2452 ;
    wire data_in_0_2;
    wire \c0.n12_adj_2472_cascade_ ;
    wire \c0.n17765 ;
    wire \c0.n8556_cascade_ ;
    wire \c0.n7_cascade_ ;
    wire \c0.n6_adj_2478 ;
    wire data_in_2_2;
    wire \c0.n8460 ;
    wire \c0.n17745 ;
    wire \c0.n16_adj_2485_cascade_ ;
    wire data_in_frame_10_6;
    wire n63_adj_2642_cascade_;
    wire n16468;
    wire data_in_7_0;
    wire \c0.n4_adj_2512_cascade_ ;
    wire n2591;
    wire \c0.n8751 ;
    wire \c0.n17532 ;
    wire n2591_cascade_;
    wire \c0.n9324 ;
    wire \c0.n17533 ;
    wire \c0.n2605 ;
    wire n2570;
    wire n2570_cascade_;
    wire \c0.n8556 ;
    wire \c0.n17_adj_2514_cascade_ ;
    wire \c0.data_in_frame_6_2 ;
    wire FRAME_MATCHER_next_state_31_N_2026_1_cascade_;
    wire n2567;
    wire \c0.n8658 ;
    wire data_in_frame_5_1;
    wire \c0.n17516 ;
    wire \c0.n2601_cascade_ ;
    wire n2597;
    wire \c0.n9039 ;
    wire \c0.n17522 ;
    wire \c0.n2606 ;
    wire \c0.n17428_cascade_ ;
    wire \c0.n11_adj_2494 ;
    wire \c0.n14 ;
    wire \c0.n17575 ;
    wire \c0.n9103 ;
    wire data_in_frame_5_2;
    wire data_in_frame_5_6;
    wire \c0.n17430 ;
    wire data_in_frame_5_4;
    wire \c0.n2603 ;
    wire n2568;
    wire \c0.n17538 ;
    wire \c0.n9355 ;
    wire n2568_cascade_;
    wire \c0.n17541 ;
    wire \c0.n21_cascade_ ;
    wire \c0.n25 ;
    wire \c0.n27_cascade_ ;
    wire \c0.n5_adj_2438 ;
    wire \c0.data_in_frame_6_7 ;
    wire \c0.n4_adj_2548 ;
    wire data_in_frame_8_4;
    wire n19_adj_2651;
    wire data_in_frame_8_3;
    wire n9380;
    wire n9054;
    wire n6_adj_2604_cascade_;
    wire data_in_frame_7_0;
    wire \c0.data_in_frame_1_7 ;
    wire \c0.data_in_frame_3_5 ;
    wire \c0.n17614 ;
    wire \c0.n8666 ;
    wire data_out_frame2_14_1;
    wire n18104;
    wire n18097;
    wire n18103;
    wire data_in_7_3;
    wire n18054;
    wire data_out_frame2_10_4;
    wire data_out_frame2_11_4;
    wire data_out_frame2_14_5;
    wire \c0.data_in_frame_10_0 ;
    wire \c0.n14631 ;
    wire data_out_frame2_12_3;
    wire data_in_20_2;
    wire \c0.n17815 ;
    wire \c0.n17818 ;
    wire \c0.n6_adj_2432 ;
    wire \c0.n18372_cascade_ ;
    wire \c0.n18375_cascade_ ;
    wire \c0.tx2.r_Tx_Data_3 ;
    wire data_out_frame2_18_3;
    wire \c0.data_out_frame2_19_3 ;
    wire data_out_frame2_16_3;
    wire \c0.n18510_cascade_ ;
    wire data_out_frame2_17_3;
    wire \c0.data_out_frame2_20_3 ;
    wire \c0.n18513_cascade_ ;
    wire \c0.n22_adj_2527 ;
    wire n9652;
    wire n9922;
    wire r_Bit_Index_2_adj_2635;
    wire \c0.n17559 ;
    wire n9135;
    wire \c0.data_out_frame2_0_3 ;
    wire \c0.n18082 ;
    wire r_Bit_Index_1_adj_2636;
    wire r_Bit_Index_0_adj_2637;
    wire n4980;
    wire bfn_6_30_0_;
    wire n225;
    wire \c0.rx.n16365 ;
    wire \c0.rx.n16366 ;
    wire \c0.rx.n16367 ;
    wire \c0.rx.n16368 ;
    wire \c0.rx.n16369 ;
    wire \c0.rx.n16370 ;
    wire \c0.rx.n16371 ;
    wire n224;
    wire n226;
    wire n221;
    wire n223;
    wire \c0.rx.n17999 ;
    wire \c0.n18444 ;
    wire \c0.n9 ;
    wire data_out_frame2_18_4;
    wire \c0.data_out_frame2_19_4 ;
    wire data_out_frame2_16_4;
    wire \c0.n18528_cascade_ ;
    wire data_out_frame2_17_4;
    wire \c0.n134 ;
    wire \c0.n18531_cascade_ ;
    wire data_out_frame2_5_4;
    wire \c0.n17955_cascade_ ;
    wire \c0.byte_transmit_counter2_2 ;
    wire \c0.data_out_frame2_0_4 ;
    wire \c0.n18456_cascade_ ;
    wire \c0.n18447 ;
    wire \c0.n18459_cascade_ ;
    wire \c0.n22_adj_2525 ;
    wire \c0.byte_transmit_counter2_3 ;
    wire \c0.n15_cascade_ ;
    wire \c0.byte_transmit_counter2_4 ;
    wire \c0.tx2.r_Tx_Data_4 ;
    wire \c0.tx2.n7727 ;
    wire data_in_2_7;
    wire data_in_4_7;
    wire data_in_4_5;
    wire data_in_3_5;
    wire \c0.n28_adj_2475_cascade_ ;
    wire \c0.n8_adj_2474 ;
    wire \c0.n8559 ;
    wire \c0.data_in_2_0 ;
    wire data_in_0_1;
    wire data_in_1_7;
    wire data_in_2_5;
    wire \c0.n17_adj_2486 ;
    wire \c0.data_in_1_3 ;
    wire \c0.data_in_0_3 ;
    wire data_in_4_3;
    wire data_in_3_3;
    wire \c0.data_in_frame_7_4 ;
    wire n2587;
    wire \c0.data_in_7_4 ;
    wire \c0.data_in_6_4 ;
    wire data_in_5_4;
    wire \c0.data_in_4_4 ;
    wire n17952;
    wire data_in_2_4;
    wire \c0.data_in_3_4 ;
    wire \c0.n17743 ;
    wire data_in_4_0;
    wire \c0.data_in_3_0 ;
    wire data_in_1_6;
    wire data_in_0_6;
    wire data_in_2_6;
    wire data_in_3_1;
    wire data_in_9_1;
    wire \c0.data_in_frame_7_5 ;
    wire data_in_frame_8_6;
    wire \c0.n17473 ;
    wire \c0.data_in_4_6 ;
    wire data_in_frame_5_7;
    wire \c0.n9368 ;
    wire \c0.n9365 ;
    wire \c0.n2600_cascade_ ;
    wire \c0.n9334 ;
    wire \c0.n10_adj_2493 ;
    wire data_in_3_6;
    wire data_in_1_2;
    wire \c0.n8572 ;
    wire data_in_frame_6_5;
    wire \c0.n4_adj_2512 ;
    wire n2594;
    wire n2573_cascade_;
    wire n17481;
    wire \c0.n9043 ;
    wire \c0.n8886 ;
    wire \c0.n15927 ;
    wire \c0.n17594 ;
    wire \c0.n17412 ;
    wire n2565_cascade_;
    wire n2574;
    wire n17547;
    wire \c0.n23_cascade_ ;
    wire \c0.n17536 ;
    wire \c0.n28 ;
    wire data_in_frame_8_0;
    wire data_in_frame_1_1;
    wire \c0.data_in_frame_10_4 ;
    wire n2563;
    wire \c0.data_in_frame_7_2 ;
    wire \c0.n8062 ;
    wire n2563_cascade_;
    wire \c0.n9204 ;
    wire \c0.n8890 ;
    wire \c0.n17592_cascade_ ;
    wire \c0.n26 ;
    wire data_in_10_1;
    wire \c0.n17544 ;
    wire \c0.n8056 ;
    wire n2566_cascade_;
    wire n2561;
    wire \c0.n19 ;
    wire data_in_9_0;
    wire \c0.data_in_frame_9_0 ;
    wire n2575;
    wire \c0.n17504 ;
    wire \c0.n6_adj_2541_cascade_ ;
    wire \c0.n17591 ;
    wire \c0.data_out_frame2_20_4 ;
    wire \c0.n17488 ;
    wire data_in_frame_9_6;
    wire n17479;
    wire n9051;
    wire n6_adj_2583;
    wire \c0.data_out_frame2_19_2 ;
    wire \c0.data_in_frame_0_1 ;
    wire \c0.data_in_frame_3_6 ;
    wire \c0.data_in_frame_2_1 ;
    wire \c0.data_in_frame_0_2 ;
    wire \c0.n10_adj_2536 ;
    wire n18101;
    wire data_in_8_3;
    wire n8517_cascade_;
    wire n17366;
    wire data_in_9_3;
    wire r_Clock_Count_0;
    wire r_Clock_Count_5;
    wire r_Clock_Count_3;
    wire r_Clock_Count_4;
    wire \c0.tx.n10_cascade_ ;
    wire r_Clock_Count_1;
    wire data_in_5_5;
    wire data_in_19_0;
    wire data_in_10_0;
    wire rx_data_4;
    wire data_in_15_2;
    wire data_in_14_2;
    wire data_in_4_2;
    wire data_in_9_7;
    wire data_in_8_7;
    wire data_out_frame2_13_0;
    wire data_in_18_5;
    wire n8562_cascade_;
    wire rx_data_2;
    wire \c0.rx.n2_cascade_ ;
    wire \c0.rx.n2 ;
    wire r_Clock_Count_0_adj_2624;
    wire r_Clock_Count_1_adj_2623;
    wire \c0.rx.n79 ;
    wire \c0.rx.n18597 ;
    wire \c0.rx.r_Rx_Data_R ;
    wire \c0.rx.n13537 ;
    wire \c0.rx.n4_adj_2424 ;
    wire \c0.rx.n17381 ;
    wire \c0.rx.n18003_cascade_ ;
    wire n13880_cascade_;
    wire \c0.rx.n10193 ;
    wire r_Clock_Count_2_adj_2622;
    wire \c0.rx.n124 ;
    wire r_Clock_Count_3_adj_2621;
    wire \c0.rx.n97_cascade_ ;
    wire \c0.rx.n17345 ;
    wire n13880;
    wire n222;
    wire r_Clock_Count_4_adj_2620;
    wire n3;
    wire \c0.rx.n18001 ;
    wire n17856_cascade_;
    wire n17855;
    wire LED_c;
    wire \c0.rx.n112 ;
    wire data_out_frame2_7_4;
    wire data_out_frame2_6_4;
    wire \c0.n5_adj_2425 ;
    wire data_out_frame2_9_4;
    wire data_out_frame2_8_4;
    wire \c0.n8 ;
    wire \c0.data_out_frame2_0_1 ;
    wire \c0.byte_transmit_counter2_1 ;
    wire \c0.byte_transmit_counter2_0 ;
    wire \c0.n18086 ;
    wire data_in_10_7;
    wire data_in_11_7;
    wire data_in_12_7;
    wire data_in_13_7;
    wire data_in_14_7;
    wire data_in_16_7;
    wire data_in_15_7;
    wire n2564;
    wire data_in_14_1;
    wire data_in_2_1;
    wire data_in_1_1;
    wire data_in_13_1;
    wire data_in_12_1;
    wire data_in_11_1;
    wire data_in_6_6;
    wire data_in_5_6;
    wire n9606;
    wire data_out_frame2_7_7;
    wire \c0.data_in_frame_9_7 ;
    wire \c0.n17433 ;
    wire data_in_7_7;
    wire n2573;
    wire \c0.data_in_frame_9_2 ;
    wire n2565;
    wire \c0.data_in_frame_10_2 ;
    wire n2566;
    wire n1396;
    wire n2571;
    wire \c0.data_in_frame_9_4 ;
    wire data_in_17_7;
    wire n7364;
    wire data_in_6_2;
    wire data_in_5_2;
    wire \c0.data_in_frame_10_5 ;
    wire n2562;
    wire data_in_10_5;
    wire data_in_9_5;
    wire data_in_12_5;
    wire data_in_11_5;
    wire n18098;
    wire \c0.n142 ;
    wire \c0.n1 ;
    wire FRAME_MATCHER_next_state_1;
    wire \c0.FRAME_MATCHER_state_0 ;
    wire \c0.n1_adj_2437 ;
    wire r_SM_Main_2_N_2323_1_cascade_;
    wire n17757_cascade_;
    wire \c0.FRAME_MATCHER_state_2 ;
    wire \c0.FRAME_MATCHER_state_1 ;
    wire \c0.n157 ;
    wire n18010;
    wire n9390;
    wire n9390_cascade_;
    wire n17681_cascade_;
    wire n16466;
    wire n17356;
    wire n18102;
    wire r_Clock_Count_2;
    wire n13601;
    wire data_in_7_2;
    wire n13597;
    wire rx_data_6;
    wire data_in_16_2;
    wire n4;
    wire rx_data_3;
    wire n4_adj_2582;
    wire data_in_20_6;
    wire data_in_8_2;
    wire n8567;
    wire data_in_11_2;
    wire data_in_13_2;
    wire data_in_12_2;
    wire FRAME_MATCHER_next_state_31_N_2026_1;
    wire n63_adj_2642;
    wire n63;
    wire FRAME_MATCHER_next_state_0;
    wire data_in_17_5;
    wire \c0.rx.r_SM_Main_2_N_2386_0 ;
    wire \c0.rx.n18066 ;
    wire rand_data_0;
    wire bfn_9_29_0_;
    wire rand_data_1;
    wire n16412;
    wire rand_data_2;
    wire n16413;
    wire rand_data_3;
    wire n16414;
    wire rand_data_4;
    wire n16415;
    wire rand_data_5;
    wire n16416;
    wire rand_data_6;
    wire rand_setpoint_6;
    wire n16417;
    wire rand_data_7;
    wire rand_setpoint_7;
    wire n16418;
    wire n16419;
    wire rand_data_8;
    wire bfn_9_30_0_;
    wire rand_data_9;
    wire n16420;
    wire rand_data_10;
    wire n16421;
    wire rand_data_11;
    wire n16422;
    wire rand_data_12;
    wire n16423;
    wire rand_data_13;
    wire n16424;
    wire rand_data_14;
    wire n16425;
    wire rand_data_15;
    wire n16426;
    wire n16427;
    wire rand_data_16;
    wire bfn_9_31_0_;
    wire rand_data_17;
    wire n16428;
    wire rand_data_18;
    wire n16429;
    wire rand_data_19;
    wire n16430;
    wire rand_data_20;
    wire n16431;
    wire rand_data_21;
    wire n16432;
    wire rand_data_22;
    wire n16433;
    wire rand_data_23;
    wire n16434;
    wire n16435;
    wire rand_data_24;
    wire bfn_9_32_0_;
    wire rand_data_25;
    wire n16436;
    wire rand_data_26;
    wire n16437;
    wire rand_data_27;
    wire n16438;
    wire rand_data_28;
    wire n16439;
    wire rand_data_29;
    wire n16440;
    wire rand_data_30;
    wire n16441;
    wire rand_data_31;
    wire n16442;
    wire data_in_1_5;
    wire data_in_7_5;
    wire data_in_6_5;
    wire data_in_8_1;
    wire \c0.data_in_7_1 ;
    wire data_in_10_3;
    wire data_in_6_7;
    wire data_in_5_7;
    wire \c0.data_in_frame_10_1 ;
    wire \c0.data_in_frame_10_3 ;
    wire \c0.n6 ;
    wire data_in_11_0;
    wire n7086;
    wire data_in_15_1;
    wire \c0.data_in_frame_9_1 ;
    wire \c0.data_in_frame_10_7 ;
    wire \c0.data_in_frame_9_5 ;
    wire \c0.data_in_frame_9_3 ;
    wire \c0.n8989 ;
    wire data_in_10_2;
    wire data_in_9_2;
    wire data_in_18_7;
    wire rx_data_7;
    wire data_in_16_3;
    wire data_in_15_3;
    wire data_in_20_7;
    wire data_in_19_7;
    wire n12123;
    wire n7080;
    wire n17767;
    wire \c0.tx.n17 ;
    wire r_Tx_Data_2;
    wire r_Clock_Count_6;
    wire r_Clock_Count_7;
    wire n1_cascade_;
    wire n3_adj_2650_cascade_;
    wire tx_o_adj_2584;
    wire \c0.n17556_cascade_ ;
    wire data_in_1_4;
    wire data_in_0_5;
    wire data_in_2_3;
    wire data_in_3_2;
    wire \c0.n16_adj_2513 ;
    wire data_in_18_0;
    wire n9796;
    wire r_Tx_Data_7;
    wire r_Bit_Index_2;
    wire n12_adj_2618;
    wire n22;
    wire n17950;
    wire r_Clock_Count_8;
    wire \c0.n6_adj_2448 ;
    wire data_in_19_6;
    wire data_in_18_6;
    wire rx_data_1;
    wire rand_setpoint_2;
    wire data_in_19_5;
    wire rx_data_5;
    wire data_in_20_5;
    wire \c0.n17911 ;
    wire \c0.n5_adj_2488 ;
    wire \c0.n18498 ;
    wire \c0.n2_adj_2487_cascade_ ;
    wire n4_adj_2649;
    wire n8562;
    wire n4_adj_2649_cascade_;
    wire r_Rx_Data;
    wire rx_data_0;
    wire data_in_20_0;
    wire data_in_17_6;
    wire data_in_16_6;
    wire rand_setpoint_4;
    wire data_in_15_6;
    wire rand_setpoint_11;
    wire rand_setpoint_25;
    wire rand_setpoint_30;
    wire rand_setpoint_31;
    wire rand_setpoint_10;
    wire r_Clock_Count_5_adj_2619;
    wire \c0.rx.r_Clock_Count_7 ;
    wire \c0.rx.n97 ;
    wire \c0.rx.r_Clock_Count_6 ;
    wire \c0.rx.r_SM_Main_2_N_2380_2_cascade_ ;
    wire \c0.rx.n18000_cascade_ ;
    wire \c0.rx.n18594 ;
    wire rand_setpoint_27;
    wire \c0.n17966_cascade_ ;
    wire rand_setpoint_29;
    wire \c0.n17970_cascade_ ;
    wire rand_setpoint_24;
    wire \c0.n17957_cascade_ ;
    wire rand_setpoint_22;
    wire data_in_19_2;
    wire data_in_20_4;
    wire data_in_19_4;
    wire data_in_18_4;
    wire data_in_18_2;
    wire data_in_17_2;
    wire data_in_8_4;
    wire data_in_9_4;
    wire data_in_10_4;
    wire data_in_11_4;
    wire data_in_12_4;
    wire data_in_13_4;
    wire data_in_14_4;
    wire data_in_11_3;
    wire data_in_15_4;
    wire data_in_17_4;
    wire data_in_16_4;
    wire data_in_4_1;
    wire \c0.n18089_cascade_ ;
    wire \c0.n18429_cascade_ ;
    wire tx_data_7_N_keep;
    wire \c0.n18017_cascade_ ;
    wire \c0.n18426 ;
    wire data_in_17_3;
    wire \c0.n5_adj_2499 ;
    wire \c0.n18378_cascade_ ;
    wire \c0.n18381_cascade_ ;
    wire tx_data_2_N_keep;
    wire data_in_20_3;
    wire data_in_13_5;
    wire data_in_19_3;
    wire data_in_18_3;
    wire data_in_12_0;
    wire data_in_12_3;
    wire n18462;
    wire n18465;
    wire data_in_9_6;
    wire data_in_8_6;
    wire data_in_16_5;
    wire data_in_14_3;
    wire data_in_13_3;
    wire n17737_cascade_;
    wire n17312;
    wire n17312_cascade_;
    wire n14_adj_2615_cascade_;
    wire data_in_17_1;
    wire data_in_16_1;
    wire n17757;
    wire r_Bit_Index_0;
    wire data_in_18_1;
    wire n18438;
    wire r_Bit_Index_1;
    wire n18441;
    wire data_in_13_0;
    wire r_Tx_Data_3;
    wire data_in_20_1;
    wire data_in_19_1;
    wire data_in_17_0;
    wire data_in_16_0;
    wire \c0.n18501 ;
    wire tx_data_0_N_keep_cascade_;
    wire r_Tx_Data_0;
    wire data_in_15_5;
    wire data_in_14_5;
    wire n4958;
    wire r_Bit_Index_2_adj_2625;
    wire n4958_cascade_;
    wire n9920_cascade_;
    wire r_Bit_Index_1_adj_2626;
    wire data_in_15_0;
    wire data_in_14_0;
    wire rand_setpoint_1;
    wire rand_setpoint_0;
    wire \c0.n8953_cascade_ ;
    wire rand_setpoint_5;
    wire \c0.n5 ;
    wire \c0.n17972 ;
    wire \c0.rx.r_SM_Main_2_N_2380_2 ;
    wire \c0.rx.n17351 ;
    wire \c0.rx.r_SM_Main_0 ;
    wire \c0.rx.n17376 ;
    wire \c0.data_out_6__2__N_803_cascade_ ;
    wire rand_setpoint_18;
    wire \c0.n2216_cascade_ ;
    wire \c0.data_out_6_2 ;
    wire rand_setpoint_26;
    wire \c0.data_out_6__2__N_803 ;
    wire \c0.n17964_cascade_ ;
    wire \c0.n17525_cascade_ ;
    wire \c0.rx.n9553 ;
    wire \c0.rx.r_SM_Main_2 ;
    wire \c0.rx.r_SM_Main_1 ;
    wire \c0.data_in_6_1 ;
    wire data_in_5_1;
    wire data_in_10_6;
    wire data_in_11_6;
    wire \c0.n17755 ;
    wire \c0.n25_adj_2517 ;
    wire \c0.n1314_cascade_ ;
    wire bfn_12_24_0_;
    wire \c0.n16305 ;
    wire \c0.n7273 ;
    wire \c0.n16306 ;
    wire \c0.n7272 ;
    wire \c0.n16307 ;
    wire \c0.n16308 ;
    wire \c0.n16309 ;
    wire \c0.n7269 ;
    wire \c0.n16310 ;
    wire \c0.n16311 ;
    wire \c0.n16312 ;
    wire \c0.n18011 ;
    wire bfn_12_25_0_;
    wire \c0.n7266 ;
    wire \c0.n16313 ;
    wire \c0.n7265 ;
    wire \c0.n16314 ;
    wire \c0.n16315 ;
    wire \c0.n16316 ;
    wire \c0.n16317 ;
    wire \c0.n16318 ;
    wire r_SM_Main_2_N_2323_1;
    wire n4_adj_2653_cascade_;
    wire r_SM_Main_2;
    wire r_SM_Main_0;
    wire r_SM_Main_1;
    wire \c0.tx_active_prev ;
    wire \c0.n17349 ;
    wire \c0.n17937 ;
    wire \c0.n18390_cascade_ ;
    wire \c0.n18393_cascade_ ;
    wire tx_data_3_N_keep;
    wire \c0.n18095 ;
    wire n9646;
    wire n9920;
    wire r_Bit_Index_0_adj_2627;
    wire \c0.data_out_6__7__N_675_cascade_ ;
    wire rand_setpoint_15;
    wire \c0.n17928_cascade_ ;
    wire rand_setpoint_14;
    wire \c0.n17465 ;
    wire \c0.n17906_cascade_ ;
    wire \c0.n17921 ;
    wire \c0.data_out_10_6 ;
    wire \c0.n2_adj_2483 ;
    wire \c0.n17389 ;
    wire \c0.n17389_cascade_ ;
    wire \c0.n17600_cascade_ ;
    wire \c0.n9658 ;
    wire \c0.n17398_cascade_ ;
    wire rand_setpoint_20;
    wire \c0.n2146_cascade_ ;
    wire \c0.data_out_5__3__N_964 ;
    wire \c0.data_out_5__3__N_964_cascade_ ;
    wire \c0.data_out_6__3__N_785_cascade_ ;
    wire rand_setpoint_19;
    wire \c0.n2181_cascade_ ;
    wire data_out_6__6__N_729;
    wire data_out_2_0;
    wire data_out_6__7__N_678;
    wire n96_cascade_;
    wire n47_cascade_;
    wire n2615;
    wire n41_cascade_;
    wire n17958;
    wire n43;
    wire \c0.n7271 ;
    wire \c0.n18105 ;
    wire \c0.n18012 ;
    wire \c0.n17936 ;
    wire \c0.n7275 ;
    wire \c0.n7274 ;
    wire \c0.n18008 ;
    wire \c0.delay_counter_3 ;
    wire \c0.delay_counter_1 ;
    wire \c0.delay_counter_2 ;
    wire \c0.delay_counter_4 ;
    wire delay_counter_0;
    wire delay_counter_13;
    wire delay_counter_14;
    wire \c0.n7264 ;
    wire n29_cascade_;
    wire data_in_12_6;
    wire \c0.n149_cascade_ ;
    wire \c0.n93 ;
    wire n8529_cascade_;
    wire \c0.n8550_cascade_ ;
    wire n121_adj_2606;
    wire n8529;
    wire n121_adj_2606_cascade_;
    wire n13_adj_2652;
    wire \c0.n251 ;
    wire bfn_13_26_0_;
    wire \c0.n16350 ;
    wire \c0.n16351 ;
    wire \c0.n16352 ;
    wire \c0.n16353 ;
    wire byte_transmit_counter_5;
    wire tx_transmit_N_2239_5;
    wire \c0.n16354 ;
    wire \c0.n16355 ;
    wire byte_transmit_counter_7;
    wire \c0.n16356 ;
    wire tx_transmit_N_2239_7;
    wire data_out_3_4;
    wire \c0.n18093_cascade_ ;
    wire \c0.n18399_cascade_ ;
    wire tx_transmit_N_2239_4;
    wire \c0.n5_adj_2447 ;
    wire \c0.n17941_cascade_ ;
    wire \c0.n18396 ;
    wire \c0.n18068 ;
    wire \c0.n5_adj_2490 ;
    wire \c0.data_out_10_4 ;
    wire \c0.n18067 ;
    wire \c0.n18092 ;
    wire \c0.n18094 ;
    wire \c0.n18096 ;
    wire \c0.n18088 ;
    wire \c0.n8634 ;
    wire \c0.n9276_cascade_ ;
    wire \c0.data_out_7__1__N_626 ;
    wire \c0.n17623_cascade_ ;
    wire rand_setpoint_8;
    wire \c0.n17916_cascade_ ;
    wire \c0.data_out_7_0 ;
    wire \c0.n8486 ;
    wire \c0.n8486_cascade_ ;
    wire \c0.n16450 ;
    wire n4_adj_2612;
    wire rand_setpoint_13;
    wire \c0.n17925_cascade_ ;
    wire rand_setpoint_12;
    wire \c0.n17931_cascade_ ;
    wire \c0.n17400 ;
    wire \c0.data_out_7__4__N_550 ;
    wire \c0.data_out_7_4 ;
    wire data_out_5__4__N_959;
    wire rand_setpoint_28;
    wire \c0.n17967_cascade_ ;
    wire \c0.n6_adj_2467 ;
    wire \c0.n9276 ;
    wire \c0.n17662_cascade_ ;
    wire rand_setpoint_23;
    wire \c0.n2041_cascade_ ;
    wire \c0.n17974 ;
    wire rand_setpoint_16;
    wire \c0.n17693_cascade_ ;
    wire \c0.data_out_6_0 ;
    wire data_out_1_7;
    wire \c0.n17578 ;
    wire \c0.delay_counter_10 ;
    wire n96;
    wire n6878;
    wire n17672_cascade_;
    wire \c0.n113 ;
    wire n17364;
    wire \c0.n18009 ;
    wire \c0.delay_counter_12 ;
    wire n119;
    wire UART_TRANSMITTER_state_7_N_1749_2_cascade_;
    wire n18032;
    wire n8488;
    wire n17709;
    wire \c0.delay_counter_6 ;
    wire \c0.delay_counter_9 ;
    wire \c0.n17753 ;
    wire n29;
    wire \c0.n7268 ;
    wire \c0.n1314 ;
    wire \c0.delay_counter_7 ;
    wire \c0.delay_counter_11 ;
    wire \c0.delay_counter_8 ;
    wire \c0.delay_counter_5 ;
    wire \c0.n10_adj_2532_cascade_ ;
    wire \c0.n14_adj_2533 ;
    wire n17306;
    wire n17306_cascade_;
    wire \c0.n17387 ;
    wire \c0.n6_adj_2534 ;
    wire tx_data_4_N_keep;
    wire r_Tx_Data_4;
    wire \c0.n16_adj_2445_cascade_ ;
    wire \c0.n19_adj_2446_cascade_ ;
    wire \c0.n8550 ;
    wire \c0.n2650 ;
    wire \c0.tx_transmit_N_2239_0 ;
    wire \c0.tx_transmit_N_2239_1 ;
    wire tx_transmit_N_2239_2;
    wire \c0.n97 ;
    wire \c0.tx_transmit ;
    wire tx_active;
    wire n13415;
    wire tx_transmit_N_2239_3;
    wire r_Tx_Data_5;
    wire n16485;
    wire \c0.n7428 ;
    wire n14_adj_2615;
    wire n9631;
    wire tx_transmit_N_2239_6;
    wire byte_transmit_counter_6;
    wire \c0.n149 ;
    wire \c0.n17741 ;
    wire r_Tx_Data_1;
    wire \c0.n18071 ;
    wire \c0.n8_adj_2526_cascade_ ;
    wire \c0.n18072 ;
    wire \c0.n17644 ;
    wire \c0.data_out_7__2__N_574 ;
    wire \c0.data_out_7__2__N_574_cascade_ ;
    wire \c0.data_out_10_2 ;
    wire \c0.data_out_9_2 ;
    wire \c0.data_out_9_3 ;
    wire \c0.n18073_cascade_ ;
    wire rand_setpoint_3;
    wire data_out_8_2;
    wire \c0.data_out_6_4 ;
    wire \c0.n9091_cascade_ ;
    wire \c0.n17566_cascade_ ;
    wire \c0.data_out_6_3 ;
    wire \c0.n9195_cascade_ ;
    wire \c0.data_out_7__4__N_556 ;
    wire \c0.n18015 ;
    wire \c0.n8_adj_2516 ;
    wire \c0.data_out_6_7 ;
    wire \c0.n9195 ;
    wire \c0.n17668_cascade_ ;
    wire \c0.n8812 ;
    wire \c0.n8_adj_2511_cascade_ ;
    wire \c0.n17623 ;
    wire \c0.n8950 ;
    wire \c0.data_out_9_0 ;
    wire \c0.data_out_10_0 ;
    wire \c0.n18016 ;
    wire \c0.data_out_2_3 ;
    wire \c0.n4_adj_2543_cascade_ ;
    wire rand_setpoint_21;
    wire \c0.n9656_cascade_ ;
    wire rand_setpoint_17;
    wire \c0.n2251_cascade_ ;
    wire \c0.n17962 ;
    wire \c0.data_out_6__1__N_849 ;
    wire \c0.data_out_1_1 ;
    wire data_out_1_2;
    wire \c0.n8767_cascade_ ;
    wire \c0.n17525 ;
    wire \c0.n17641 ;
    wire \c0.n17457_cascade_ ;
    wire \c0.n8964 ;
    wire \c0.n17415 ;
    wire \c0.data_out_6__3__N_788 ;
    wire \c0.n17415_cascade_ ;
    wire \c0.data_out_5_2 ;
    wire rand_setpoint_9;
    wire \c0.n9518 ;
    wire data_out_6__2__N_804;
    wire \c0.n17457 ;
    wire \c0.n17654 ;
    wire \c0.n18061 ;
    wire \c0.data_out_7__5__N_543 ;
    wire data_out_6__1__N_850;
    wire \c0.n2 ;
    wire \c0.n18060 ;
    wire data_out_0_5;
    wire \c0.n18065_cascade_ ;
    wire tx_data_5_N_keep;
    wire \c0.n18014 ;
    wire tx_data_1_N_keep;
    wire \c0.n17943 ;
    wire \c0.n5_adj_2481_cascade_ ;
    wire \c0.n18091 ;
    wire \c0.n18402_cascade_ ;
    wire \c0.n2_adj_2476 ;
    wire \c0.n18405 ;
    wire \c0.data_out_5_1 ;
    wire \c0.n45_adj_2518_cascade_ ;
    wire \c0.n1_adj_2522 ;
    wire \c0.n46_cascade_ ;
    wire \c0.n44_adj_2524 ;
    wire \c0.n8_adj_2531 ;
    wire \c0.n18069_cascade_ ;
    wire \c0.n18070 ;
    wire rx_data_ready;
    wire data_in_14_6;
    wire data_in_13_6;
    wire \c0.n17445 ;
    wire \c0.n17510 ;
    wire \c0.data_out_9_1 ;
    wire data_out_8_1;
    wire \c0.n8_adj_2519 ;
    wire \c0.n8_adj_2535 ;
    wire \c0.n17398 ;
    wire \c0.n9091 ;
    wire \c0.data_out_9_4 ;
    wire \c0.data_out_6_1 ;
    wire \c0.n17499 ;
    wire \c0.n6_adj_2451 ;
    wire \c0.data_out_10_5 ;
    wire \c0.n18064 ;
    wire \c0.n17668 ;
    wire \c0.n9087 ;
    wire \c0.n8_adj_2528_cascade_ ;
    wire \c0.data_out_10_1 ;
    wire \c0.n17556 ;
    wire \c0.data_out_6__7__N_675 ;
    wire \c0.data_out_10_7 ;
    wire \c0.n8600 ;
    wire \c0.data_out_5_3 ;
    wire \c0.n17635_cascade_ ;
    wire \c0.n17922 ;
    wire \c0.data_out_7__7__N_519 ;
    wire \c0.data_out_7_5 ;
    wire \c0.n17492 ;
    wire \c0.n17635 ;
    wire \c0.n17492_cascade_ ;
    wire \c0.data_out_10_3 ;
    wire \c0.data_out_7_2 ;
    wire \c0.n17600 ;
    wire \c0.data_out_9_6 ;
    wire \c0.data_out_7_1 ;
    wire \c0.n17454 ;
    wire \c0.data_out_6_5 ;
    wire \c0.data_out_6__5__N_752 ;
    wire \c0.n17454_cascade_ ;
    wire \c0.data_out_9_5 ;
    wire \c0.n8_adj_2537 ;
    wire \c0.n17626 ;
    wire \c0.n17608 ;
    wire \c0.n8970 ;
    wire \c0.n17662 ;
    wire data_out_8_6;
    wire \c0.n17665 ;
    wire \c0.n12_adj_2482_cascade_ ;
    wire \c0.data_out_7_3 ;
    wire data_out_10__7__N_114;
    wire \c0.data_out_9_7 ;
    wire data_out_8_7;
    wire \c0.n8_adj_2538 ;
    wire \c0.data_out_0_6 ;
    wire data_out_0_3;
    wire data_out_0_1;
    wire data_out_0_0;
    wire \c0.n8926 ;
    wire \c0.n8767 ;
    wire \c0.n8926_cascade_ ;
    wire n2720;
    wire UART_TRANSMITTER_state_0;
    wire n4430;
    wire data_out_1_6;
    wire data_out_3_5;
    wire UART_TRANSMITTER_state_1;
    wire n9519;
    wire data_out_5__7__N_931;
    wire \c0.data_out_6__4__N_765 ;
    wire \c0.n1_adj_2484 ;
    wire \c0.n18414_cascade_ ;
    wire byte_transmit_counter_4;
    wire \c0.n18417_cascade_ ;
    wire byte_transmit_counter_3;
    wire n7734;
    wire tx_data_6_N_keep_cascade_;
    wire r_Tx_Data_6;
    wire \c0.data_out_7__6__N_530 ;
    wire \c0.n17949 ;
    wire data_out_3_6;
    wire \c0.n18090 ;
    wire \c0.byte_transmit_counter_0 ;
    wire \c0.data_out_7_6 ;
    wire \c0.n5_adj_2444 ;
    wire \c0.n8_adj_2539 ;
    wire byte_transmit_counter_2;
    wire \c0.n18062 ;
    wire \c0.byte_transmit_counter_1 ;
    wire \c0.n18063 ;
    wire data_out_8_0;
    wire \c0.data_out_7_7 ;
    wire \c0.n17638 ;
    wire n26;
    wire bfn_16_29_0_;
    wire n25;
    wire n16380;
    wire n24;
    wire n16381;
    wire n23;
    wire n16382;
    wire n22_adj_2655;
    wire n16383;
    wire n21;
    wire n16384;
    wire n20;
    wire n16385;
    wire n19;
    wire n16386;
    wire n16387;
    wire n18;
    wire bfn_16_30_0_;
    wire n17;
    wire n16388;
    wire n16;
    wire n16389;
    wire n15;
    wire n16390;
    wire n14;
    wire n16391;
    wire n13;
    wire n16392;
    wire n12;
    wire n16393;
    wire n11;
    wire n16394;
    wire n16395;
    wire n10;
    wire bfn_16_31_0_;
    wire n9;
    wire n16396;
    wire n8_adj_2617;
    wire n16397;
    wire n7;
    wire n16398;
    wire n6;
    wire n16399;
    wire blink_counter_21;
    wire n16400;
    wire blink_counter_22;
    wire n16401;
    wire blink_counter_23;
    wire n16402;
    wire n16403;
    wire blink_counter_24;
    wire bfn_16_32_0_;
    wire n16404;
    wire blink_counter_25;
    wire CLK_c;
    wire \c0.data_out_5__5__N_950 ;
    wire \c0.n17438 ;
    wire \c0.data_out_6__3__N_781 ;
    wire \c0.n17653 ;
    wire \c0.n17976 ;
    wire \c0.n8953 ;
    wire data_out_8_5;
    wire \c0.data_out_6_6 ;
    wire \c0.n8922 ;
    wire data_out_8_4;
    wire data_out_8_3;
    wire \c0.n17620 ;
    wire \c0.n17611 ;
    wire \c0.n17659 ;
    wire \c0.n8777 ;
    wire UART_TRANSMITTER_state_2;
    wire \c0.n17918 ;
    wire _gnd_net_;

    defparam LED_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam LED_pad_iopad.PULLUP=1'b0;
    IO_PAD LED_pad_iopad (
            .OE(N__50526),
            .DIN(N__50525),
            .DOUT(N__50524),
            .PACKAGEPIN(LED));
    defparam LED_pad_preio.PIN_TYPE=6'b011001;
    defparam LED_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO LED_pad_preio (
            .PADOEN(N__50526),
            .PADOUT(N__50525),
            .PADIN(N__50524),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__30263),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam USBPU_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam USBPU_pad_iopad.PULLUP=1'b0;
    IO_PAD USBPU_pad_iopad (
            .OE(N__50517),
            .DIN(N__50516),
            .DOUT(N__50515),
            .PACKAGEPIN(USBPU));
    defparam USBPU_pad_preio.PIN_TYPE=6'b011001;
    defparam USBPU_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO USBPU_pad_preio (
            .PADOEN(N__50517),
            .PADOUT(N__50516),
            .PADIN(N__50515),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam rx_input_iopad.IO_STANDARD="SB_LVCMOS";
    defparam rx_input_iopad.PULLUP=1'b1;
    IO_PAD rx_input_iopad (
            .OE(N__50508),
            .DIN(N__50507),
            .DOUT(N__50506),
            .PACKAGEPIN(PIN_2));
    defparam rx_input_preio.PIN_TYPE=6'b000000;
    defparam rx_input_preio.NEG_TRIGGER=1'b0;
    PRE_IO rx_input_preio (
            .PADOEN(N__50508),
            .PADOUT(N__50507),
            .PADIN(N__50506),
            .CLOCKENABLE(VCCG0),
            .DIN0(\c0.rx.r_Rx_Data_R ),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(GNDG0),
            .INPUTCLK(N__50364),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam tx2_output_iopad.IO_STANDARD="SB_LVCMOS";
    defparam tx2_output_iopad.PULLUP=1'b1;
    IO_PAD tx2_output_iopad (
            .OE(N__50499),
            .DIN(N__50498),
            .DOUT(N__50497),
            .PACKAGEPIN(PIN_3));
    defparam tx2_output_preio.PIN_TYPE=6'b101001;
    defparam tx2_output_preio.NEG_TRIGGER=1'b0;
    PRE_IO tx2_output_preio (
            .PADOEN(N__50499),
            .PADOUT(N__50498),
            .PADIN(N__50497),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__21152),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__21122));
    defparam tx_output_iopad.IO_STANDARD="SB_LVCMOS";
    defparam tx_output_iopad.PULLUP=1'b1;
    IO_PAD tx_output_iopad (
            .OE(N__50490),
            .DIN(N__50489),
            .DOUT(N__50488),
            .PACKAGEPIN(PIN_1));
    defparam tx_output_preio.PIN_TYPE=6'b101001;
    defparam tx_output_preio.NEG_TRIGGER=1'b0;
    PRE_IO tx_output_preio (
            .PADOEN(N__50490),
            .PADOUT(N__50489),
            .PADIN(N__50488),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__37175),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__21161));
    defparam CLK_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam CLK_pad_iopad.PULLUP=1'b0;
    IO_PAD CLK_pad_iopad (
            .OE(N__50481),
            .DIN(N__50480),
            .DOUT(N__50479),
            .PACKAGEPIN(CLK));
    defparam CLK_pad_preio.PIN_TYPE=6'b000001;
    defparam CLK_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO CLK_pad_preio (
            .PADOEN(N__50481),
            .PADOUT(N__50480),
            .PADIN(N__50479),
            .CLOCKENABLE(),
            .DIN0(CLK_pad_gb_input),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    InMux I__12591 (
            .O(N__50462),
            .I(n16404));
    InMux I__12590 (
            .O(N__50459),
            .I(N__50456));
    LocalMux I__12589 (
            .O(N__50456),
            .I(N__50453));
    Span4Mux_v I__12588 (
            .O(N__50453),
            .I(N__50450));
    Span4Mux_h I__12587 (
            .O(N__50450),
            .I(N__50447));
    Span4Mux_h I__12586 (
            .O(N__50447),
            .I(N__50443));
    InMux I__12585 (
            .O(N__50446),
            .I(N__50440));
    Odrv4 I__12584 (
            .O(N__50443),
            .I(blink_counter_25));
    LocalMux I__12583 (
            .O(N__50440),
            .I(blink_counter_25));
    ClkMux I__12582 (
            .O(N__50435),
            .I(N__49880));
    ClkMux I__12581 (
            .O(N__50434),
            .I(N__49880));
    ClkMux I__12580 (
            .O(N__50433),
            .I(N__49880));
    ClkMux I__12579 (
            .O(N__50432),
            .I(N__49880));
    ClkMux I__12578 (
            .O(N__50431),
            .I(N__49880));
    ClkMux I__12577 (
            .O(N__50430),
            .I(N__49880));
    ClkMux I__12576 (
            .O(N__50429),
            .I(N__49880));
    ClkMux I__12575 (
            .O(N__50428),
            .I(N__49880));
    ClkMux I__12574 (
            .O(N__50427),
            .I(N__49880));
    ClkMux I__12573 (
            .O(N__50426),
            .I(N__49880));
    ClkMux I__12572 (
            .O(N__50425),
            .I(N__49880));
    ClkMux I__12571 (
            .O(N__50424),
            .I(N__49880));
    ClkMux I__12570 (
            .O(N__50423),
            .I(N__49880));
    ClkMux I__12569 (
            .O(N__50422),
            .I(N__49880));
    ClkMux I__12568 (
            .O(N__50421),
            .I(N__49880));
    ClkMux I__12567 (
            .O(N__50420),
            .I(N__49880));
    ClkMux I__12566 (
            .O(N__50419),
            .I(N__49880));
    ClkMux I__12565 (
            .O(N__50418),
            .I(N__49880));
    ClkMux I__12564 (
            .O(N__50417),
            .I(N__49880));
    ClkMux I__12563 (
            .O(N__50416),
            .I(N__49880));
    ClkMux I__12562 (
            .O(N__50415),
            .I(N__49880));
    ClkMux I__12561 (
            .O(N__50414),
            .I(N__49880));
    ClkMux I__12560 (
            .O(N__50413),
            .I(N__49880));
    ClkMux I__12559 (
            .O(N__50412),
            .I(N__49880));
    ClkMux I__12558 (
            .O(N__50411),
            .I(N__49880));
    ClkMux I__12557 (
            .O(N__50410),
            .I(N__49880));
    ClkMux I__12556 (
            .O(N__50409),
            .I(N__49880));
    ClkMux I__12555 (
            .O(N__50408),
            .I(N__49880));
    ClkMux I__12554 (
            .O(N__50407),
            .I(N__49880));
    ClkMux I__12553 (
            .O(N__50406),
            .I(N__49880));
    ClkMux I__12552 (
            .O(N__50405),
            .I(N__49880));
    ClkMux I__12551 (
            .O(N__50404),
            .I(N__49880));
    ClkMux I__12550 (
            .O(N__50403),
            .I(N__49880));
    ClkMux I__12549 (
            .O(N__50402),
            .I(N__49880));
    ClkMux I__12548 (
            .O(N__50401),
            .I(N__49880));
    ClkMux I__12547 (
            .O(N__50400),
            .I(N__49880));
    ClkMux I__12546 (
            .O(N__50399),
            .I(N__49880));
    ClkMux I__12545 (
            .O(N__50398),
            .I(N__49880));
    ClkMux I__12544 (
            .O(N__50397),
            .I(N__49880));
    ClkMux I__12543 (
            .O(N__50396),
            .I(N__49880));
    ClkMux I__12542 (
            .O(N__50395),
            .I(N__49880));
    ClkMux I__12541 (
            .O(N__50394),
            .I(N__49880));
    ClkMux I__12540 (
            .O(N__50393),
            .I(N__49880));
    ClkMux I__12539 (
            .O(N__50392),
            .I(N__49880));
    ClkMux I__12538 (
            .O(N__50391),
            .I(N__49880));
    ClkMux I__12537 (
            .O(N__50390),
            .I(N__49880));
    ClkMux I__12536 (
            .O(N__50389),
            .I(N__49880));
    ClkMux I__12535 (
            .O(N__50388),
            .I(N__49880));
    ClkMux I__12534 (
            .O(N__50387),
            .I(N__49880));
    ClkMux I__12533 (
            .O(N__50386),
            .I(N__49880));
    ClkMux I__12532 (
            .O(N__50385),
            .I(N__49880));
    ClkMux I__12531 (
            .O(N__50384),
            .I(N__49880));
    ClkMux I__12530 (
            .O(N__50383),
            .I(N__49880));
    ClkMux I__12529 (
            .O(N__50382),
            .I(N__49880));
    ClkMux I__12528 (
            .O(N__50381),
            .I(N__49880));
    ClkMux I__12527 (
            .O(N__50380),
            .I(N__49880));
    ClkMux I__12526 (
            .O(N__50379),
            .I(N__49880));
    ClkMux I__12525 (
            .O(N__50378),
            .I(N__49880));
    ClkMux I__12524 (
            .O(N__50377),
            .I(N__49880));
    ClkMux I__12523 (
            .O(N__50376),
            .I(N__49880));
    ClkMux I__12522 (
            .O(N__50375),
            .I(N__49880));
    ClkMux I__12521 (
            .O(N__50374),
            .I(N__49880));
    ClkMux I__12520 (
            .O(N__50373),
            .I(N__49880));
    ClkMux I__12519 (
            .O(N__50372),
            .I(N__49880));
    ClkMux I__12518 (
            .O(N__50371),
            .I(N__49880));
    ClkMux I__12517 (
            .O(N__50370),
            .I(N__49880));
    ClkMux I__12516 (
            .O(N__50369),
            .I(N__49880));
    ClkMux I__12515 (
            .O(N__50368),
            .I(N__49880));
    ClkMux I__12514 (
            .O(N__50367),
            .I(N__49880));
    ClkMux I__12513 (
            .O(N__50366),
            .I(N__49880));
    ClkMux I__12512 (
            .O(N__50365),
            .I(N__49880));
    ClkMux I__12511 (
            .O(N__50364),
            .I(N__49880));
    ClkMux I__12510 (
            .O(N__50363),
            .I(N__49880));
    ClkMux I__12509 (
            .O(N__50362),
            .I(N__49880));
    ClkMux I__12508 (
            .O(N__50361),
            .I(N__49880));
    ClkMux I__12507 (
            .O(N__50360),
            .I(N__49880));
    ClkMux I__12506 (
            .O(N__50359),
            .I(N__49880));
    ClkMux I__12505 (
            .O(N__50358),
            .I(N__49880));
    ClkMux I__12504 (
            .O(N__50357),
            .I(N__49880));
    ClkMux I__12503 (
            .O(N__50356),
            .I(N__49880));
    ClkMux I__12502 (
            .O(N__50355),
            .I(N__49880));
    ClkMux I__12501 (
            .O(N__50354),
            .I(N__49880));
    ClkMux I__12500 (
            .O(N__50353),
            .I(N__49880));
    ClkMux I__12499 (
            .O(N__50352),
            .I(N__49880));
    ClkMux I__12498 (
            .O(N__50351),
            .I(N__49880));
    ClkMux I__12497 (
            .O(N__50350),
            .I(N__49880));
    ClkMux I__12496 (
            .O(N__50349),
            .I(N__49880));
    ClkMux I__12495 (
            .O(N__50348),
            .I(N__49880));
    ClkMux I__12494 (
            .O(N__50347),
            .I(N__49880));
    ClkMux I__12493 (
            .O(N__50346),
            .I(N__49880));
    ClkMux I__12492 (
            .O(N__50345),
            .I(N__49880));
    ClkMux I__12491 (
            .O(N__50344),
            .I(N__49880));
    ClkMux I__12490 (
            .O(N__50343),
            .I(N__49880));
    ClkMux I__12489 (
            .O(N__50342),
            .I(N__49880));
    ClkMux I__12488 (
            .O(N__50341),
            .I(N__49880));
    ClkMux I__12487 (
            .O(N__50340),
            .I(N__49880));
    ClkMux I__12486 (
            .O(N__50339),
            .I(N__49880));
    ClkMux I__12485 (
            .O(N__50338),
            .I(N__49880));
    ClkMux I__12484 (
            .O(N__50337),
            .I(N__49880));
    ClkMux I__12483 (
            .O(N__50336),
            .I(N__49880));
    ClkMux I__12482 (
            .O(N__50335),
            .I(N__49880));
    ClkMux I__12481 (
            .O(N__50334),
            .I(N__49880));
    ClkMux I__12480 (
            .O(N__50333),
            .I(N__49880));
    ClkMux I__12479 (
            .O(N__50332),
            .I(N__49880));
    ClkMux I__12478 (
            .O(N__50331),
            .I(N__49880));
    ClkMux I__12477 (
            .O(N__50330),
            .I(N__49880));
    ClkMux I__12476 (
            .O(N__50329),
            .I(N__49880));
    ClkMux I__12475 (
            .O(N__50328),
            .I(N__49880));
    ClkMux I__12474 (
            .O(N__50327),
            .I(N__49880));
    ClkMux I__12473 (
            .O(N__50326),
            .I(N__49880));
    ClkMux I__12472 (
            .O(N__50325),
            .I(N__49880));
    ClkMux I__12471 (
            .O(N__50324),
            .I(N__49880));
    ClkMux I__12470 (
            .O(N__50323),
            .I(N__49880));
    ClkMux I__12469 (
            .O(N__50322),
            .I(N__49880));
    ClkMux I__12468 (
            .O(N__50321),
            .I(N__49880));
    ClkMux I__12467 (
            .O(N__50320),
            .I(N__49880));
    ClkMux I__12466 (
            .O(N__50319),
            .I(N__49880));
    ClkMux I__12465 (
            .O(N__50318),
            .I(N__49880));
    ClkMux I__12464 (
            .O(N__50317),
            .I(N__49880));
    ClkMux I__12463 (
            .O(N__50316),
            .I(N__49880));
    ClkMux I__12462 (
            .O(N__50315),
            .I(N__49880));
    ClkMux I__12461 (
            .O(N__50314),
            .I(N__49880));
    ClkMux I__12460 (
            .O(N__50313),
            .I(N__49880));
    ClkMux I__12459 (
            .O(N__50312),
            .I(N__49880));
    ClkMux I__12458 (
            .O(N__50311),
            .I(N__49880));
    ClkMux I__12457 (
            .O(N__50310),
            .I(N__49880));
    ClkMux I__12456 (
            .O(N__50309),
            .I(N__49880));
    ClkMux I__12455 (
            .O(N__50308),
            .I(N__49880));
    ClkMux I__12454 (
            .O(N__50307),
            .I(N__49880));
    ClkMux I__12453 (
            .O(N__50306),
            .I(N__49880));
    ClkMux I__12452 (
            .O(N__50305),
            .I(N__49880));
    ClkMux I__12451 (
            .O(N__50304),
            .I(N__49880));
    ClkMux I__12450 (
            .O(N__50303),
            .I(N__49880));
    ClkMux I__12449 (
            .O(N__50302),
            .I(N__49880));
    ClkMux I__12448 (
            .O(N__50301),
            .I(N__49880));
    ClkMux I__12447 (
            .O(N__50300),
            .I(N__49880));
    ClkMux I__12446 (
            .O(N__50299),
            .I(N__49880));
    ClkMux I__12445 (
            .O(N__50298),
            .I(N__49880));
    ClkMux I__12444 (
            .O(N__50297),
            .I(N__49880));
    ClkMux I__12443 (
            .O(N__50296),
            .I(N__49880));
    ClkMux I__12442 (
            .O(N__50295),
            .I(N__49880));
    ClkMux I__12441 (
            .O(N__50294),
            .I(N__49880));
    ClkMux I__12440 (
            .O(N__50293),
            .I(N__49880));
    ClkMux I__12439 (
            .O(N__50292),
            .I(N__49880));
    ClkMux I__12438 (
            .O(N__50291),
            .I(N__49880));
    ClkMux I__12437 (
            .O(N__50290),
            .I(N__49880));
    ClkMux I__12436 (
            .O(N__50289),
            .I(N__49880));
    ClkMux I__12435 (
            .O(N__50288),
            .I(N__49880));
    ClkMux I__12434 (
            .O(N__50287),
            .I(N__49880));
    ClkMux I__12433 (
            .O(N__50286),
            .I(N__49880));
    ClkMux I__12432 (
            .O(N__50285),
            .I(N__49880));
    ClkMux I__12431 (
            .O(N__50284),
            .I(N__49880));
    ClkMux I__12430 (
            .O(N__50283),
            .I(N__49880));
    ClkMux I__12429 (
            .O(N__50282),
            .I(N__49880));
    ClkMux I__12428 (
            .O(N__50281),
            .I(N__49880));
    ClkMux I__12427 (
            .O(N__50280),
            .I(N__49880));
    ClkMux I__12426 (
            .O(N__50279),
            .I(N__49880));
    ClkMux I__12425 (
            .O(N__50278),
            .I(N__49880));
    ClkMux I__12424 (
            .O(N__50277),
            .I(N__49880));
    ClkMux I__12423 (
            .O(N__50276),
            .I(N__49880));
    ClkMux I__12422 (
            .O(N__50275),
            .I(N__49880));
    ClkMux I__12421 (
            .O(N__50274),
            .I(N__49880));
    ClkMux I__12420 (
            .O(N__50273),
            .I(N__49880));
    ClkMux I__12419 (
            .O(N__50272),
            .I(N__49880));
    ClkMux I__12418 (
            .O(N__50271),
            .I(N__49880));
    ClkMux I__12417 (
            .O(N__50270),
            .I(N__49880));
    ClkMux I__12416 (
            .O(N__50269),
            .I(N__49880));
    ClkMux I__12415 (
            .O(N__50268),
            .I(N__49880));
    ClkMux I__12414 (
            .O(N__50267),
            .I(N__49880));
    ClkMux I__12413 (
            .O(N__50266),
            .I(N__49880));
    ClkMux I__12412 (
            .O(N__50265),
            .I(N__49880));
    ClkMux I__12411 (
            .O(N__50264),
            .I(N__49880));
    ClkMux I__12410 (
            .O(N__50263),
            .I(N__49880));
    ClkMux I__12409 (
            .O(N__50262),
            .I(N__49880));
    ClkMux I__12408 (
            .O(N__50261),
            .I(N__49880));
    ClkMux I__12407 (
            .O(N__50260),
            .I(N__49880));
    ClkMux I__12406 (
            .O(N__50259),
            .I(N__49880));
    ClkMux I__12405 (
            .O(N__50258),
            .I(N__49880));
    ClkMux I__12404 (
            .O(N__50257),
            .I(N__49880));
    ClkMux I__12403 (
            .O(N__50256),
            .I(N__49880));
    ClkMux I__12402 (
            .O(N__50255),
            .I(N__49880));
    ClkMux I__12401 (
            .O(N__50254),
            .I(N__49880));
    ClkMux I__12400 (
            .O(N__50253),
            .I(N__49880));
    ClkMux I__12399 (
            .O(N__50252),
            .I(N__49880));
    ClkMux I__12398 (
            .O(N__50251),
            .I(N__49880));
    GlobalMux I__12397 (
            .O(N__49880),
            .I(N__49877));
    gio2CtrlBuf I__12396 (
            .O(N__49877),
            .I(CLK_c));
    InMux I__12395 (
            .O(N__49874),
            .I(N__49869));
    InMux I__12394 (
            .O(N__49873),
            .I(N__49863));
    InMux I__12393 (
            .O(N__49872),
            .I(N__49860));
    LocalMux I__12392 (
            .O(N__49869),
            .I(N__49857));
    InMux I__12391 (
            .O(N__49868),
            .I(N__49854));
    InMux I__12390 (
            .O(N__49867),
            .I(N__49850));
    InMux I__12389 (
            .O(N__49866),
            .I(N__49847));
    LocalMux I__12388 (
            .O(N__49863),
            .I(N__49843));
    LocalMux I__12387 (
            .O(N__49860),
            .I(N__49836));
    Span4Mux_h I__12386 (
            .O(N__49857),
            .I(N__49836));
    LocalMux I__12385 (
            .O(N__49854),
            .I(N__49836));
    InMux I__12384 (
            .O(N__49853),
            .I(N__49833));
    LocalMux I__12383 (
            .O(N__49850),
            .I(N__49830));
    LocalMux I__12382 (
            .O(N__49847),
            .I(N__49827));
    InMux I__12381 (
            .O(N__49846),
            .I(N__49824));
    Span4Mux_h I__12380 (
            .O(N__49843),
            .I(N__49819));
    Span4Mux_v I__12379 (
            .O(N__49836),
            .I(N__49819));
    LocalMux I__12378 (
            .O(N__49833),
            .I(\c0.data_out_5__5__N_950 ));
    Odrv4 I__12377 (
            .O(N__49830),
            .I(\c0.data_out_5__5__N_950 ));
    Odrv4 I__12376 (
            .O(N__49827),
            .I(\c0.data_out_5__5__N_950 ));
    LocalMux I__12375 (
            .O(N__49824),
            .I(\c0.data_out_5__5__N_950 ));
    Odrv4 I__12374 (
            .O(N__49819),
            .I(\c0.data_out_5__5__N_950 ));
    InMux I__12373 (
            .O(N__49808),
            .I(N__49804));
    InMux I__12372 (
            .O(N__49807),
            .I(N__49801));
    LocalMux I__12371 (
            .O(N__49804),
            .I(N__49798));
    LocalMux I__12370 (
            .O(N__49801),
            .I(\c0.n17438 ));
    Odrv4 I__12369 (
            .O(N__49798),
            .I(\c0.n17438 ));
    CascadeMux I__12368 (
            .O(N__49793),
            .I(N__49787));
    InMux I__12367 (
            .O(N__49792),
            .I(N__49784));
    InMux I__12366 (
            .O(N__49791),
            .I(N__49780));
    InMux I__12365 (
            .O(N__49790),
            .I(N__49777));
    InMux I__12364 (
            .O(N__49787),
            .I(N__49774));
    LocalMux I__12363 (
            .O(N__49784),
            .I(N__49771));
    InMux I__12362 (
            .O(N__49783),
            .I(N__49768));
    LocalMux I__12361 (
            .O(N__49780),
            .I(N__49763));
    LocalMux I__12360 (
            .O(N__49777),
            .I(N__49763));
    LocalMux I__12359 (
            .O(N__49774),
            .I(N__49760));
    Span4Mux_h I__12358 (
            .O(N__49771),
            .I(N__49755));
    LocalMux I__12357 (
            .O(N__49768),
            .I(N__49755));
    Odrv12 I__12356 (
            .O(N__49763),
            .I(\c0.data_out_6__3__N_781 ));
    Odrv4 I__12355 (
            .O(N__49760),
            .I(\c0.data_out_6__3__N_781 ));
    Odrv4 I__12354 (
            .O(N__49755),
            .I(\c0.data_out_6__3__N_781 ));
    InMux I__12353 (
            .O(N__49748),
            .I(N__49745));
    LocalMux I__12352 (
            .O(N__49745),
            .I(N__49741));
    InMux I__12351 (
            .O(N__49744),
            .I(N__49738));
    Span4Mux_h I__12350 (
            .O(N__49741),
            .I(N__49733));
    LocalMux I__12349 (
            .O(N__49738),
            .I(N__49733));
    Odrv4 I__12348 (
            .O(N__49733),
            .I(\c0.n17653 ));
    InMux I__12347 (
            .O(N__49730),
            .I(N__49727));
    LocalMux I__12346 (
            .O(N__49727),
            .I(N__49724));
    Odrv4 I__12345 (
            .O(N__49724),
            .I(\c0.n17976 ));
    InMux I__12344 (
            .O(N__49721),
            .I(N__49718));
    LocalMux I__12343 (
            .O(N__49718),
            .I(N__49715));
    Span4Mux_h I__12342 (
            .O(N__49715),
            .I(N__49712));
    Odrv4 I__12341 (
            .O(N__49712),
            .I(\c0.n8953 ));
    CascadeMux I__12340 (
            .O(N__49709),
            .I(N__49703));
    InMux I__12339 (
            .O(N__49708),
            .I(N__49698));
    InMux I__12338 (
            .O(N__49707),
            .I(N__49698));
    InMux I__12337 (
            .O(N__49706),
            .I(N__49694));
    InMux I__12336 (
            .O(N__49703),
            .I(N__49691));
    LocalMux I__12335 (
            .O(N__49698),
            .I(N__49688));
    InMux I__12334 (
            .O(N__49697),
            .I(N__49685));
    LocalMux I__12333 (
            .O(N__49694),
            .I(N__49682));
    LocalMux I__12332 (
            .O(N__49691),
            .I(N__49679));
    Span4Mux_s3_v I__12331 (
            .O(N__49688),
            .I(N__49676));
    LocalMux I__12330 (
            .O(N__49685),
            .I(data_out_8_5));
    Odrv4 I__12329 (
            .O(N__49682),
            .I(data_out_8_5));
    Odrv12 I__12328 (
            .O(N__49679),
            .I(data_out_8_5));
    Odrv4 I__12327 (
            .O(N__49676),
            .I(data_out_8_5));
    InMux I__12326 (
            .O(N__49667),
            .I(N__49664));
    LocalMux I__12325 (
            .O(N__49664),
            .I(N__49660));
    InMux I__12324 (
            .O(N__49663),
            .I(N__49657));
    Span4Mux_v I__12323 (
            .O(N__49660),
            .I(N__49652));
    LocalMux I__12322 (
            .O(N__49657),
            .I(N__49652));
    Span4Mux_h I__12321 (
            .O(N__49652),
            .I(N__49648));
    InMux I__12320 (
            .O(N__49651),
            .I(N__49645));
    Span4Mux_v I__12319 (
            .O(N__49648),
            .I(N__49642));
    LocalMux I__12318 (
            .O(N__49645),
            .I(\c0.data_out_6_6 ));
    Odrv4 I__12317 (
            .O(N__49642),
            .I(\c0.data_out_6_6 ));
    InMux I__12316 (
            .O(N__49637),
            .I(N__49634));
    LocalMux I__12315 (
            .O(N__49634),
            .I(N__49630));
    InMux I__12314 (
            .O(N__49633),
            .I(N__49627));
    Span12Mux_h I__12313 (
            .O(N__49630),
            .I(N__49624));
    LocalMux I__12312 (
            .O(N__49627),
            .I(N__49621));
    Odrv12 I__12311 (
            .O(N__49624),
            .I(\c0.n8922 ));
    Odrv4 I__12310 (
            .O(N__49621),
            .I(\c0.n8922 ));
    InMux I__12309 (
            .O(N__49616),
            .I(N__49612));
    InMux I__12308 (
            .O(N__49615),
            .I(N__49607));
    LocalMux I__12307 (
            .O(N__49612),
            .I(N__49604));
    InMux I__12306 (
            .O(N__49611),
            .I(N__49598));
    InMux I__12305 (
            .O(N__49610),
            .I(N__49598));
    LocalMux I__12304 (
            .O(N__49607),
            .I(N__49595));
    Span4Mux_h I__12303 (
            .O(N__49604),
            .I(N__49592));
    InMux I__12302 (
            .O(N__49603),
            .I(N__49589));
    LocalMux I__12301 (
            .O(N__49598),
            .I(N__49586));
    Span4Mux_h I__12300 (
            .O(N__49595),
            .I(N__49581));
    Span4Mux_h I__12299 (
            .O(N__49592),
            .I(N__49581));
    LocalMux I__12298 (
            .O(N__49589),
            .I(data_out_8_4));
    Odrv12 I__12297 (
            .O(N__49586),
            .I(data_out_8_4));
    Odrv4 I__12296 (
            .O(N__49581),
            .I(data_out_8_4));
    InMux I__12295 (
            .O(N__49574),
            .I(N__49571));
    LocalMux I__12294 (
            .O(N__49571),
            .I(N__49568));
    Span4Mux_h I__12293 (
            .O(N__49568),
            .I(N__49562));
    InMux I__12292 (
            .O(N__49567),
            .I(N__49555));
    InMux I__12291 (
            .O(N__49566),
            .I(N__49555));
    InMux I__12290 (
            .O(N__49565),
            .I(N__49555));
    Odrv4 I__12289 (
            .O(N__49562),
            .I(data_out_8_3));
    LocalMux I__12288 (
            .O(N__49555),
            .I(data_out_8_3));
    InMux I__12287 (
            .O(N__49550),
            .I(N__49546));
    InMux I__12286 (
            .O(N__49549),
            .I(N__49543));
    LocalMux I__12285 (
            .O(N__49546),
            .I(N__49540));
    LocalMux I__12284 (
            .O(N__49543),
            .I(N__49537));
    Span4Mux_s3_v I__12283 (
            .O(N__49540),
            .I(N__49534));
    Span4Mux_h I__12282 (
            .O(N__49537),
            .I(N__49531));
    Odrv4 I__12281 (
            .O(N__49534),
            .I(\c0.n17620 ));
    Odrv4 I__12280 (
            .O(N__49531),
            .I(\c0.n17620 ));
    InMux I__12279 (
            .O(N__49526),
            .I(N__49523));
    LocalMux I__12278 (
            .O(N__49523),
            .I(N__49520));
    Span4Mux_h I__12277 (
            .O(N__49520),
            .I(N__49516));
    InMux I__12276 (
            .O(N__49519),
            .I(N__49513));
    Span4Mux_h I__12275 (
            .O(N__49516),
            .I(N__49510));
    LocalMux I__12274 (
            .O(N__49513),
            .I(\c0.n17611 ));
    Odrv4 I__12273 (
            .O(N__49510),
            .I(\c0.n17611 ));
    InMux I__12272 (
            .O(N__49505),
            .I(N__49501));
    InMux I__12271 (
            .O(N__49504),
            .I(N__49498));
    LocalMux I__12270 (
            .O(N__49501),
            .I(N__49493));
    LocalMux I__12269 (
            .O(N__49498),
            .I(N__49493));
    Span4Mux_h I__12268 (
            .O(N__49493),
            .I(N__49490));
    Odrv4 I__12267 (
            .O(N__49490),
            .I(\c0.n17659 ));
    CascadeMux I__12266 (
            .O(N__49487),
            .I(N__49483));
    CascadeMux I__12265 (
            .O(N__49486),
            .I(N__49480));
    InMux I__12264 (
            .O(N__49483),
            .I(N__49477));
    InMux I__12263 (
            .O(N__49480),
            .I(N__49473));
    LocalMux I__12262 (
            .O(N__49477),
            .I(N__49470));
    InMux I__12261 (
            .O(N__49476),
            .I(N__49467));
    LocalMux I__12260 (
            .O(N__49473),
            .I(N__49464));
    Span4Mux_h I__12259 (
            .O(N__49470),
            .I(N__49461));
    LocalMux I__12258 (
            .O(N__49467),
            .I(N__49456));
    Span4Mux_h I__12257 (
            .O(N__49464),
            .I(N__49456));
    Odrv4 I__12256 (
            .O(N__49461),
            .I(\c0.n8777 ));
    Odrv4 I__12255 (
            .O(N__49456),
            .I(\c0.n8777 ));
    InMux I__12254 (
            .O(N__49451),
            .I(N__49437));
    InMux I__12253 (
            .O(N__49450),
            .I(N__49437));
    CascadeMux I__12252 (
            .O(N__49449),
            .I(N__49432));
    InMux I__12251 (
            .O(N__49448),
            .I(N__49427));
    InMux I__12250 (
            .O(N__49447),
            .I(N__49427));
    InMux I__12249 (
            .O(N__49446),
            .I(N__49424));
    CascadeMux I__12248 (
            .O(N__49445),
            .I(N__49411));
    InMux I__12247 (
            .O(N__49444),
            .I(N__49404));
    InMux I__12246 (
            .O(N__49443),
            .I(N__49404));
    InMux I__12245 (
            .O(N__49442),
            .I(N__49404));
    LocalMux I__12244 (
            .O(N__49437),
            .I(N__49401));
    InMux I__12243 (
            .O(N__49436),
            .I(N__49398));
    InMux I__12242 (
            .O(N__49435),
            .I(N__49392));
    InMux I__12241 (
            .O(N__49432),
            .I(N__49392));
    LocalMux I__12240 (
            .O(N__49427),
            .I(N__49389));
    LocalMux I__12239 (
            .O(N__49424),
            .I(N__49386));
    InMux I__12238 (
            .O(N__49423),
            .I(N__49378));
    InMux I__12237 (
            .O(N__49422),
            .I(N__49378));
    InMux I__12236 (
            .O(N__49421),
            .I(N__49371));
    InMux I__12235 (
            .O(N__49420),
            .I(N__49371));
    InMux I__12234 (
            .O(N__49419),
            .I(N__49371));
    InMux I__12233 (
            .O(N__49418),
            .I(N__49368));
    InMux I__12232 (
            .O(N__49417),
            .I(N__49365));
    InMux I__12231 (
            .O(N__49416),
            .I(N__49356));
    InMux I__12230 (
            .O(N__49415),
            .I(N__49356));
    InMux I__12229 (
            .O(N__49414),
            .I(N__49356));
    InMux I__12228 (
            .O(N__49411),
            .I(N__49353));
    LocalMux I__12227 (
            .O(N__49404),
            .I(N__49350));
    Span4Mux_s3_v I__12226 (
            .O(N__49401),
            .I(N__49347));
    LocalMux I__12225 (
            .O(N__49398),
            .I(N__49344));
    InMux I__12224 (
            .O(N__49397),
            .I(N__49341));
    LocalMux I__12223 (
            .O(N__49392),
            .I(N__49334));
    Span4Mux_s3_v I__12222 (
            .O(N__49389),
            .I(N__49334));
    Span4Mux_s3_v I__12221 (
            .O(N__49386),
            .I(N__49334));
    InMux I__12220 (
            .O(N__49385),
            .I(N__49329));
    InMux I__12219 (
            .O(N__49384),
            .I(N__49329));
    InMux I__12218 (
            .O(N__49383),
            .I(N__49318));
    LocalMux I__12217 (
            .O(N__49378),
            .I(N__49309));
    LocalMux I__12216 (
            .O(N__49371),
            .I(N__49309));
    LocalMux I__12215 (
            .O(N__49368),
            .I(N__49309));
    LocalMux I__12214 (
            .O(N__49365),
            .I(N__49309));
    CascadeMux I__12213 (
            .O(N__49364),
            .I(N__49305));
    CascadeMux I__12212 (
            .O(N__49363),
            .I(N__49301));
    LocalMux I__12211 (
            .O(N__49356),
            .I(N__49298));
    LocalMux I__12210 (
            .O(N__49353),
            .I(N__49295));
    Span4Mux_s3_v I__12209 (
            .O(N__49350),
            .I(N__49292));
    Span4Mux_h I__12208 (
            .O(N__49347),
            .I(N__49282));
    Span4Mux_h I__12207 (
            .O(N__49344),
            .I(N__49282));
    LocalMux I__12206 (
            .O(N__49341),
            .I(N__49282));
    Span4Mux_h I__12205 (
            .O(N__49334),
            .I(N__49277));
    LocalMux I__12204 (
            .O(N__49329),
            .I(N__49277));
    InMux I__12203 (
            .O(N__49328),
            .I(N__49272));
    InMux I__12202 (
            .O(N__49327),
            .I(N__49272));
    InMux I__12201 (
            .O(N__49326),
            .I(N__49267));
    InMux I__12200 (
            .O(N__49325),
            .I(N__49267));
    InMux I__12199 (
            .O(N__49324),
            .I(N__49264));
    InMux I__12198 (
            .O(N__49323),
            .I(N__49257));
    InMux I__12197 (
            .O(N__49322),
            .I(N__49257));
    InMux I__12196 (
            .O(N__49321),
            .I(N__49257));
    LocalMux I__12195 (
            .O(N__49318),
            .I(N__49248));
    Span4Mux_s3_v I__12194 (
            .O(N__49309),
            .I(N__49248));
    CascadeMux I__12193 (
            .O(N__49308),
            .I(N__49245));
    InMux I__12192 (
            .O(N__49305),
            .I(N__49237));
    InMux I__12191 (
            .O(N__49304),
            .I(N__49237));
    InMux I__12190 (
            .O(N__49301),
            .I(N__49237));
    Span4Mux_s3_v I__12189 (
            .O(N__49298),
            .I(N__49230));
    Span4Mux_s3_v I__12188 (
            .O(N__49295),
            .I(N__49230));
    Span4Mux_h I__12187 (
            .O(N__49292),
            .I(N__49230));
    InMux I__12186 (
            .O(N__49291),
            .I(N__49223));
    InMux I__12185 (
            .O(N__49290),
            .I(N__49223));
    InMux I__12184 (
            .O(N__49289),
            .I(N__49223));
    Sp12to4 I__12183 (
            .O(N__49282),
            .I(N__49218));
    Sp12to4 I__12182 (
            .O(N__49277),
            .I(N__49218));
    LocalMux I__12181 (
            .O(N__49272),
            .I(N__49209));
    LocalMux I__12180 (
            .O(N__49267),
            .I(N__49209));
    LocalMux I__12179 (
            .O(N__49264),
            .I(N__49209));
    LocalMux I__12178 (
            .O(N__49257),
            .I(N__49209));
    InMux I__12177 (
            .O(N__49256),
            .I(N__49204));
    InMux I__12176 (
            .O(N__49255),
            .I(N__49204));
    InMux I__12175 (
            .O(N__49254),
            .I(N__49199));
    InMux I__12174 (
            .O(N__49253),
            .I(N__49199));
    Span4Mux_v I__12173 (
            .O(N__49248),
            .I(N__49196));
    InMux I__12172 (
            .O(N__49245),
            .I(N__49191));
    InMux I__12171 (
            .O(N__49244),
            .I(N__49191));
    LocalMux I__12170 (
            .O(N__49237),
            .I(N__49184));
    Span4Mux_v I__12169 (
            .O(N__49230),
            .I(N__49184));
    LocalMux I__12168 (
            .O(N__49223),
            .I(N__49184));
    Span12Mux_s10_v I__12167 (
            .O(N__49218),
            .I(N__49181));
    Span12Mux_s5_v I__12166 (
            .O(N__49209),
            .I(N__49176));
    LocalMux I__12165 (
            .O(N__49204),
            .I(N__49176));
    LocalMux I__12164 (
            .O(N__49199),
            .I(UART_TRANSMITTER_state_2));
    Odrv4 I__12163 (
            .O(N__49196),
            .I(UART_TRANSMITTER_state_2));
    LocalMux I__12162 (
            .O(N__49191),
            .I(UART_TRANSMITTER_state_2));
    Odrv4 I__12161 (
            .O(N__49184),
            .I(UART_TRANSMITTER_state_2));
    Odrv12 I__12160 (
            .O(N__49181),
            .I(UART_TRANSMITTER_state_2));
    Odrv12 I__12159 (
            .O(N__49176),
            .I(UART_TRANSMITTER_state_2));
    InMux I__12158 (
            .O(N__49163),
            .I(N__49160));
    LocalMux I__12157 (
            .O(N__49160),
            .I(N__49157));
    Span4Mux_h I__12156 (
            .O(N__49157),
            .I(N__49154));
    Odrv4 I__12155 (
            .O(N__49154),
            .I(\c0.n17918 ));
    InMux I__12154 (
            .O(N__49151),
            .I(bfn_16_31_0_));
    InMux I__12153 (
            .O(N__49148),
            .I(N__49145));
    LocalMux I__12152 (
            .O(N__49145),
            .I(n9));
    InMux I__12151 (
            .O(N__49142),
            .I(n16396));
    InMux I__12150 (
            .O(N__49139),
            .I(N__49136));
    LocalMux I__12149 (
            .O(N__49136),
            .I(n8_adj_2617));
    InMux I__12148 (
            .O(N__49133),
            .I(n16397));
    InMux I__12147 (
            .O(N__49130),
            .I(N__49127));
    LocalMux I__12146 (
            .O(N__49127),
            .I(n7));
    InMux I__12145 (
            .O(N__49124),
            .I(n16398));
    InMux I__12144 (
            .O(N__49121),
            .I(N__49118));
    LocalMux I__12143 (
            .O(N__49118),
            .I(n6));
    InMux I__12142 (
            .O(N__49115),
            .I(n16399));
    CascadeMux I__12141 (
            .O(N__49112),
            .I(N__49108));
    InMux I__12140 (
            .O(N__49111),
            .I(N__49103));
    InMux I__12139 (
            .O(N__49108),
            .I(N__49103));
    LocalMux I__12138 (
            .O(N__49103),
            .I(N__49099));
    InMux I__12137 (
            .O(N__49102),
            .I(N__49096));
    Odrv12 I__12136 (
            .O(N__49099),
            .I(blink_counter_21));
    LocalMux I__12135 (
            .O(N__49096),
            .I(blink_counter_21));
    InMux I__12134 (
            .O(N__49091),
            .I(n16400));
    InMux I__12133 (
            .O(N__49088),
            .I(N__49082));
    InMux I__12132 (
            .O(N__49087),
            .I(N__49082));
    LocalMux I__12131 (
            .O(N__49082),
            .I(N__49079));
    Span12Mux_h I__12130 (
            .O(N__49079),
            .I(N__49075));
    InMux I__12129 (
            .O(N__49078),
            .I(N__49072));
    Odrv12 I__12128 (
            .O(N__49075),
            .I(blink_counter_22));
    LocalMux I__12127 (
            .O(N__49072),
            .I(blink_counter_22));
    InMux I__12126 (
            .O(N__49067),
            .I(n16401));
    InMux I__12125 (
            .O(N__49064),
            .I(N__49058));
    InMux I__12124 (
            .O(N__49063),
            .I(N__49058));
    LocalMux I__12123 (
            .O(N__49058),
            .I(N__49054));
    InMux I__12122 (
            .O(N__49057),
            .I(N__49051));
    Odrv12 I__12121 (
            .O(N__49054),
            .I(blink_counter_23));
    LocalMux I__12120 (
            .O(N__49051),
            .I(blink_counter_23));
    InMux I__12119 (
            .O(N__49046),
            .I(n16402));
    CascadeMux I__12118 (
            .O(N__49043),
            .I(N__49040));
    InMux I__12117 (
            .O(N__49040),
            .I(N__49034));
    InMux I__12116 (
            .O(N__49039),
            .I(N__49034));
    LocalMux I__12115 (
            .O(N__49034),
            .I(N__49031));
    Span4Mux_v I__12114 (
            .O(N__49031),
            .I(N__49028));
    Span4Mux_h I__12113 (
            .O(N__49028),
            .I(N__49025));
    Span4Mux_h I__12112 (
            .O(N__49025),
            .I(N__49021));
    InMux I__12111 (
            .O(N__49024),
            .I(N__49018));
    Odrv4 I__12110 (
            .O(N__49021),
            .I(blink_counter_24));
    LocalMux I__12109 (
            .O(N__49018),
            .I(blink_counter_24));
    InMux I__12108 (
            .O(N__49013),
            .I(bfn_16_32_0_));
    InMux I__12107 (
            .O(N__49010),
            .I(N__49007));
    LocalMux I__12106 (
            .O(N__49007),
            .I(n18));
    InMux I__12105 (
            .O(N__49004),
            .I(bfn_16_30_0_));
    InMux I__12104 (
            .O(N__49001),
            .I(N__48998));
    LocalMux I__12103 (
            .O(N__48998),
            .I(n17));
    InMux I__12102 (
            .O(N__48995),
            .I(n16388));
    InMux I__12101 (
            .O(N__48992),
            .I(N__48989));
    LocalMux I__12100 (
            .O(N__48989),
            .I(n16));
    InMux I__12099 (
            .O(N__48986),
            .I(n16389));
    InMux I__12098 (
            .O(N__48983),
            .I(N__48980));
    LocalMux I__12097 (
            .O(N__48980),
            .I(n15));
    InMux I__12096 (
            .O(N__48977),
            .I(n16390));
    InMux I__12095 (
            .O(N__48974),
            .I(N__48971));
    LocalMux I__12094 (
            .O(N__48971),
            .I(n14));
    InMux I__12093 (
            .O(N__48968),
            .I(n16391));
    InMux I__12092 (
            .O(N__48965),
            .I(N__48962));
    LocalMux I__12091 (
            .O(N__48962),
            .I(n13));
    InMux I__12090 (
            .O(N__48959),
            .I(n16392));
    InMux I__12089 (
            .O(N__48956),
            .I(N__48953));
    LocalMux I__12088 (
            .O(N__48953),
            .I(n12));
    InMux I__12087 (
            .O(N__48950),
            .I(n16393));
    InMux I__12086 (
            .O(N__48947),
            .I(N__48944));
    LocalMux I__12085 (
            .O(N__48944),
            .I(n11));
    InMux I__12084 (
            .O(N__48941),
            .I(n16394));
    InMux I__12083 (
            .O(N__48938),
            .I(N__48935));
    LocalMux I__12082 (
            .O(N__48935),
            .I(n10));
    InMux I__12081 (
            .O(N__48932),
            .I(N__48929));
    LocalMux I__12080 (
            .O(N__48929),
            .I(n26));
    InMux I__12079 (
            .O(N__48926),
            .I(bfn_16_29_0_));
    InMux I__12078 (
            .O(N__48923),
            .I(N__48920));
    LocalMux I__12077 (
            .O(N__48920),
            .I(n25));
    InMux I__12076 (
            .O(N__48917),
            .I(n16380));
    InMux I__12075 (
            .O(N__48914),
            .I(N__48911));
    LocalMux I__12074 (
            .O(N__48911),
            .I(n24));
    InMux I__12073 (
            .O(N__48908),
            .I(n16381));
    InMux I__12072 (
            .O(N__48905),
            .I(N__48902));
    LocalMux I__12071 (
            .O(N__48902),
            .I(n23));
    InMux I__12070 (
            .O(N__48899),
            .I(n16382));
    InMux I__12069 (
            .O(N__48896),
            .I(N__48893));
    LocalMux I__12068 (
            .O(N__48893),
            .I(n22_adj_2655));
    InMux I__12067 (
            .O(N__48890),
            .I(n16383));
    InMux I__12066 (
            .O(N__48887),
            .I(N__48884));
    LocalMux I__12065 (
            .O(N__48884),
            .I(n21));
    InMux I__12064 (
            .O(N__48881),
            .I(n16384));
    InMux I__12063 (
            .O(N__48878),
            .I(N__48875));
    LocalMux I__12062 (
            .O(N__48875),
            .I(n20));
    InMux I__12061 (
            .O(N__48872),
            .I(n16385));
    InMux I__12060 (
            .O(N__48869),
            .I(N__48866));
    LocalMux I__12059 (
            .O(N__48866),
            .I(n19));
    InMux I__12058 (
            .O(N__48863),
            .I(n16386));
    InMux I__12057 (
            .O(N__48860),
            .I(N__48857));
    LocalMux I__12056 (
            .O(N__48857),
            .I(N__48854));
    Span4Mux_v I__12055 (
            .O(N__48854),
            .I(N__48851));
    Odrv4 I__12054 (
            .O(N__48851),
            .I(\c0.n1_adj_2484 ));
    CascadeMux I__12053 (
            .O(N__48848),
            .I(\c0.n18414_cascade_ ));
    InMux I__12052 (
            .O(N__48845),
            .I(N__48841));
    InMux I__12051 (
            .O(N__48844),
            .I(N__48834));
    LocalMux I__12050 (
            .O(N__48841),
            .I(N__48830));
    InMux I__12049 (
            .O(N__48840),
            .I(N__48825));
    InMux I__12048 (
            .O(N__48839),
            .I(N__48825));
    InMux I__12047 (
            .O(N__48838),
            .I(N__48822));
    InMux I__12046 (
            .O(N__48837),
            .I(N__48819));
    LocalMux I__12045 (
            .O(N__48834),
            .I(N__48816));
    CascadeMux I__12044 (
            .O(N__48833),
            .I(N__48812));
    Span4Mux_h I__12043 (
            .O(N__48830),
            .I(N__48808));
    LocalMux I__12042 (
            .O(N__48825),
            .I(N__48805));
    LocalMux I__12041 (
            .O(N__48822),
            .I(N__48801));
    LocalMux I__12040 (
            .O(N__48819),
            .I(N__48798));
    Span4Mux_h I__12039 (
            .O(N__48816),
            .I(N__48795));
    InMux I__12038 (
            .O(N__48815),
            .I(N__48792));
    InMux I__12037 (
            .O(N__48812),
            .I(N__48787));
    InMux I__12036 (
            .O(N__48811),
            .I(N__48787));
    Span4Mux_v I__12035 (
            .O(N__48808),
            .I(N__48782));
    Span4Mux_h I__12034 (
            .O(N__48805),
            .I(N__48782));
    InMux I__12033 (
            .O(N__48804),
            .I(N__48779));
    Odrv4 I__12032 (
            .O(N__48801),
            .I(byte_transmit_counter_4));
    Odrv4 I__12031 (
            .O(N__48798),
            .I(byte_transmit_counter_4));
    Odrv4 I__12030 (
            .O(N__48795),
            .I(byte_transmit_counter_4));
    LocalMux I__12029 (
            .O(N__48792),
            .I(byte_transmit_counter_4));
    LocalMux I__12028 (
            .O(N__48787),
            .I(byte_transmit_counter_4));
    Odrv4 I__12027 (
            .O(N__48782),
            .I(byte_transmit_counter_4));
    LocalMux I__12026 (
            .O(N__48779),
            .I(byte_transmit_counter_4));
    CascadeMux I__12025 (
            .O(N__48764),
            .I(\c0.n18417_cascade_ ));
    CascadeMux I__12024 (
            .O(N__48761),
            .I(N__48756));
    InMux I__12023 (
            .O(N__48760),
            .I(N__48751));
    InMux I__12022 (
            .O(N__48759),
            .I(N__48748));
    InMux I__12021 (
            .O(N__48756),
            .I(N__48745));
    InMux I__12020 (
            .O(N__48755),
            .I(N__48742));
    InMux I__12019 (
            .O(N__48754),
            .I(N__48739));
    LocalMux I__12018 (
            .O(N__48751),
            .I(N__48733));
    LocalMux I__12017 (
            .O(N__48748),
            .I(N__48730));
    LocalMux I__12016 (
            .O(N__48745),
            .I(N__48725));
    LocalMux I__12015 (
            .O(N__48742),
            .I(N__48725));
    LocalMux I__12014 (
            .O(N__48739),
            .I(N__48721));
    InMux I__12013 (
            .O(N__48738),
            .I(N__48717));
    InMux I__12012 (
            .O(N__48737),
            .I(N__48712));
    InMux I__12011 (
            .O(N__48736),
            .I(N__48712));
    Span4Mux_h I__12010 (
            .O(N__48733),
            .I(N__48705));
    Span4Mux_h I__12009 (
            .O(N__48730),
            .I(N__48705));
    Span4Mux_h I__12008 (
            .O(N__48725),
            .I(N__48705));
    InMux I__12007 (
            .O(N__48724),
            .I(N__48702));
    Span4Mux_h I__12006 (
            .O(N__48721),
            .I(N__48699));
    InMux I__12005 (
            .O(N__48720),
            .I(N__48696));
    LocalMux I__12004 (
            .O(N__48717),
            .I(byte_transmit_counter_3));
    LocalMux I__12003 (
            .O(N__48712),
            .I(byte_transmit_counter_3));
    Odrv4 I__12002 (
            .O(N__48705),
            .I(byte_transmit_counter_3));
    LocalMux I__12001 (
            .O(N__48702),
            .I(byte_transmit_counter_3));
    Odrv4 I__12000 (
            .O(N__48699),
            .I(byte_transmit_counter_3));
    LocalMux I__11999 (
            .O(N__48696),
            .I(byte_transmit_counter_3));
    InMux I__11998 (
            .O(N__48683),
            .I(N__48679));
    InMux I__11997 (
            .O(N__48682),
            .I(N__48676));
    LocalMux I__11996 (
            .O(N__48679),
            .I(N__48671));
    LocalMux I__11995 (
            .O(N__48676),
            .I(N__48668));
    InMux I__11994 (
            .O(N__48675),
            .I(N__48665));
    InMux I__11993 (
            .O(N__48674),
            .I(N__48662));
    Span4Mux_h I__11992 (
            .O(N__48671),
            .I(N__48657));
    Span4Mux_v I__11991 (
            .O(N__48668),
            .I(N__48652));
    LocalMux I__11990 (
            .O(N__48665),
            .I(N__48652));
    LocalMux I__11989 (
            .O(N__48662),
            .I(N__48649));
    InMux I__11988 (
            .O(N__48661),
            .I(N__48643));
    InMux I__11987 (
            .O(N__48660),
            .I(N__48643));
    Span4Mux_v I__11986 (
            .O(N__48657),
            .I(N__48635));
    Span4Mux_h I__11985 (
            .O(N__48652),
            .I(N__48635));
    Span4Mux_h I__11984 (
            .O(N__48649),
            .I(N__48635));
    InMux I__11983 (
            .O(N__48648),
            .I(N__48632));
    LocalMux I__11982 (
            .O(N__48643),
            .I(N__48629));
    InMux I__11981 (
            .O(N__48642),
            .I(N__48626));
    Odrv4 I__11980 (
            .O(N__48635),
            .I(n7734));
    LocalMux I__11979 (
            .O(N__48632),
            .I(n7734));
    Odrv12 I__11978 (
            .O(N__48629),
            .I(n7734));
    LocalMux I__11977 (
            .O(N__48626),
            .I(n7734));
    CascadeMux I__11976 (
            .O(N__48617),
            .I(tx_data_6_N_keep_cascade_));
    InMux I__11975 (
            .O(N__48614),
            .I(N__48611));
    LocalMux I__11974 (
            .O(N__48611),
            .I(N__48608));
    Span4Mux_h I__11973 (
            .O(N__48608),
            .I(N__48604));
    InMux I__11972 (
            .O(N__48607),
            .I(N__48601));
    Span4Mux_h I__11971 (
            .O(N__48604),
            .I(N__48598));
    LocalMux I__11970 (
            .O(N__48601),
            .I(r_Tx_Data_6));
    Odrv4 I__11969 (
            .O(N__48598),
            .I(r_Tx_Data_6));
    InMux I__11968 (
            .O(N__48593),
            .I(N__48586));
    InMux I__11967 (
            .O(N__48592),
            .I(N__48583));
    InMux I__11966 (
            .O(N__48591),
            .I(N__48580));
    InMux I__11965 (
            .O(N__48590),
            .I(N__48577));
    InMux I__11964 (
            .O(N__48589),
            .I(N__48574));
    LocalMux I__11963 (
            .O(N__48586),
            .I(N__48571));
    LocalMux I__11962 (
            .O(N__48583),
            .I(N__48564));
    LocalMux I__11961 (
            .O(N__48580),
            .I(N__48564));
    LocalMux I__11960 (
            .O(N__48577),
            .I(N__48561));
    LocalMux I__11959 (
            .O(N__48574),
            .I(N__48556));
    Span4Mux_h I__11958 (
            .O(N__48571),
            .I(N__48556));
    InMux I__11957 (
            .O(N__48570),
            .I(N__48553));
    InMux I__11956 (
            .O(N__48569),
            .I(N__48550));
    Span4Mux_h I__11955 (
            .O(N__48564),
            .I(N__48547));
    Span4Mux_h I__11954 (
            .O(N__48561),
            .I(N__48542));
    Span4Mux_h I__11953 (
            .O(N__48556),
            .I(N__48542));
    LocalMux I__11952 (
            .O(N__48553),
            .I(\c0.data_out_7__6__N_530 ));
    LocalMux I__11951 (
            .O(N__48550),
            .I(\c0.data_out_7__6__N_530 ));
    Odrv4 I__11950 (
            .O(N__48547),
            .I(\c0.data_out_7__6__N_530 ));
    Odrv4 I__11949 (
            .O(N__48542),
            .I(\c0.data_out_7__6__N_530 ));
    InMux I__11948 (
            .O(N__48533),
            .I(N__48530));
    LocalMux I__11947 (
            .O(N__48530),
            .I(\c0.n17949 ));
    CascadeMux I__11946 (
            .O(N__48527),
            .I(N__48523));
    InMux I__11945 (
            .O(N__48526),
            .I(N__48519));
    InMux I__11944 (
            .O(N__48523),
            .I(N__48516));
    InMux I__11943 (
            .O(N__48522),
            .I(N__48513));
    LocalMux I__11942 (
            .O(N__48519),
            .I(N__48510));
    LocalMux I__11941 (
            .O(N__48516),
            .I(N__48507));
    LocalMux I__11940 (
            .O(N__48513),
            .I(N__48504));
    Span4Mux_v I__11939 (
            .O(N__48510),
            .I(N__48496));
    Span4Mux_v I__11938 (
            .O(N__48507),
            .I(N__48496));
    Span4Mux_v I__11937 (
            .O(N__48504),
            .I(N__48493));
    InMux I__11936 (
            .O(N__48503),
            .I(N__48486));
    InMux I__11935 (
            .O(N__48502),
            .I(N__48486));
    InMux I__11934 (
            .O(N__48501),
            .I(N__48486));
    Odrv4 I__11933 (
            .O(N__48496),
            .I(data_out_3_6));
    Odrv4 I__11932 (
            .O(N__48493),
            .I(data_out_3_6));
    LocalMux I__11931 (
            .O(N__48486),
            .I(data_out_3_6));
    InMux I__11930 (
            .O(N__48479),
            .I(N__48476));
    LocalMux I__11929 (
            .O(N__48476),
            .I(\c0.n18090 ));
    InMux I__11928 (
            .O(N__48473),
            .I(N__48470));
    LocalMux I__11927 (
            .O(N__48470),
            .I(N__48454));
    InMux I__11926 (
            .O(N__48469),
            .I(N__48447));
    InMux I__11925 (
            .O(N__48468),
            .I(N__48447));
    InMux I__11924 (
            .O(N__48467),
            .I(N__48447));
    InMux I__11923 (
            .O(N__48466),
            .I(N__48440));
    InMux I__11922 (
            .O(N__48465),
            .I(N__48440));
    InMux I__11921 (
            .O(N__48464),
            .I(N__48440));
    InMux I__11920 (
            .O(N__48463),
            .I(N__48433));
    InMux I__11919 (
            .O(N__48462),
            .I(N__48433));
    InMux I__11918 (
            .O(N__48461),
            .I(N__48433));
    InMux I__11917 (
            .O(N__48460),
            .I(N__48422));
    InMux I__11916 (
            .O(N__48459),
            .I(N__48404));
    InMux I__11915 (
            .O(N__48458),
            .I(N__48404));
    InMux I__11914 (
            .O(N__48457),
            .I(N__48404));
    Span4Mux_s3_v I__11913 (
            .O(N__48454),
            .I(N__48385));
    LocalMux I__11912 (
            .O(N__48447),
            .I(N__48385));
    LocalMux I__11911 (
            .O(N__48440),
            .I(N__48385));
    LocalMux I__11910 (
            .O(N__48433),
            .I(N__48385));
    InMux I__11909 (
            .O(N__48432),
            .I(N__48378));
    InMux I__11908 (
            .O(N__48431),
            .I(N__48378));
    InMux I__11907 (
            .O(N__48430),
            .I(N__48378));
    InMux I__11906 (
            .O(N__48429),
            .I(N__48373));
    InMux I__11905 (
            .O(N__48428),
            .I(N__48368));
    InMux I__11904 (
            .O(N__48427),
            .I(N__48368));
    InMux I__11903 (
            .O(N__48426),
            .I(N__48365));
    InMux I__11902 (
            .O(N__48425),
            .I(N__48362));
    LocalMux I__11901 (
            .O(N__48422),
            .I(N__48359));
    InMux I__11900 (
            .O(N__48421),
            .I(N__48354));
    InMux I__11899 (
            .O(N__48420),
            .I(N__48354));
    InMux I__11898 (
            .O(N__48419),
            .I(N__48349));
    InMux I__11897 (
            .O(N__48418),
            .I(N__48349));
    InMux I__11896 (
            .O(N__48417),
            .I(N__48344));
    InMux I__11895 (
            .O(N__48416),
            .I(N__48344));
    InMux I__11894 (
            .O(N__48415),
            .I(N__48333));
    InMux I__11893 (
            .O(N__48414),
            .I(N__48333));
    InMux I__11892 (
            .O(N__48413),
            .I(N__48333));
    InMux I__11891 (
            .O(N__48412),
            .I(N__48333));
    InMux I__11890 (
            .O(N__48411),
            .I(N__48333));
    LocalMux I__11889 (
            .O(N__48404),
            .I(N__48330));
    InMux I__11888 (
            .O(N__48403),
            .I(N__48325));
    InMux I__11887 (
            .O(N__48402),
            .I(N__48325));
    InMux I__11886 (
            .O(N__48401),
            .I(N__48318));
    InMux I__11885 (
            .O(N__48400),
            .I(N__48318));
    InMux I__11884 (
            .O(N__48399),
            .I(N__48318));
    CascadeMux I__11883 (
            .O(N__48398),
            .I(N__48315));
    InMux I__11882 (
            .O(N__48397),
            .I(N__48307));
    InMux I__11881 (
            .O(N__48396),
            .I(N__48307));
    InMux I__11880 (
            .O(N__48395),
            .I(N__48303));
    InMux I__11879 (
            .O(N__48394),
            .I(N__48300));
    Span4Mux_v I__11878 (
            .O(N__48385),
            .I(N__48295));
    LocalMux I__11877 (
            .O(N__48378),
            .I(N__48295));
    InMux I__11876 (
            .O(N__48377),
            .I(N__48292));
    InMux I__11875 (
            .O(N__48376),
            .I(N__48289));
    LocalMux I__11874 (
            .O(N__48373),
            .I(N__48284));
    LocalMux I__11873 (
            .O(N__48368),
            .I(N__48284));
    LocalMux I__11872 (
            .O(N__48365),
            .I(N__48281));
    LocalMux I__11871 (
            .O(N__48362),
            .I(N__48274));
    Span4Mux_h I__11870 (
            .O(N__48359),
            .I(N__48274));
    LocalMux I__11869 (
            .O(N__48354),
            .I(N__48274));
    LocalMux I__11868 (
            .O(N__48349),
            .I(N__48261));
    LocalMux I__11867 (
            .O(N__48344),
            .I(N__48261));
    LocalMux I__11866 (
            .O(N__48333),
            .I(N__48261));
    Span4Mux_h I__11865 (
            .O(N__48330),
            .I(N__48261));
    LocalMux I__11864 (
            .O(N__48325),
            .I(N__48261));
    LocalMux I__11863 (
            .O(N__48318),
            .I(N__48261));
    InMux I__11862 (
            .O(N__48315),
            .I(N__48258));
    InMux I__11861 (
            .O(N__48314),
            .I(N__48255));
    InMux I__11860 (
            .O(N__48313),
            .I(N__48250));
    InMux I__11859 (
            .O(N__48312),
            .I(N__48250));
    LocalMux I__11858 (
            .O(N__48307),
            .I(N__48247));
    InMux I__11857 (
            .O(N__48306),
            .I(N__48244));
    LocalMux I__11856 (
            .O(N__48303),
            .I(N__48237));
    LocalMux I__11855 (
            .O(N__48300),
            .I(N__48237));
    Span4Mux_h I__11854 (
            .O(N__48295),
            .I(N__48237));
    LocalMux I__11853 (
            .O(N__48292),
            .I(N__48222));
    LocalMux I__11852 (
            .O(N__48289),
            .I(N__48222));
    Span4Mux_h I__11851 (
            .O(N__48284),
            .I(N__48222));
    Span4Mux_v I__11850 (
            .O(N__48281),
            .I(N__48222));
    Span4Mux_v I__11849 (
            .O(N__48274),
            .I(N__48222));
    Span4Mux_v I__11848 (
            .O(N__48261),
            .I(N__48222));
    LocalMux I__11847 (
            .O(N__48258),
            .I(N__48222));
    LocalMux I__11846 (
            .O(N__48255),
            .I(\c0.byte_transmit_counter_0 ));
    LocalMux I__11845 (
            .O(N__48250),
            .I(\c0.byte_transmit_counter_0 ));
    Odrv12 I__11844 (
            .O(N__48247),
            .I(\c0.byte_transmit_counter_0 ));
    LocalMux I__11843 (
            .O(N__48244),
            .I(\c0.byte_transmit_counter_0 ));
    Odrv4 I__11842 (
            .O(N__48237),
            .I(\c0.byte_transmit_counter_0 ));
    Odrv4 I__11841 (
            .O(N__48222),
            .I(\c0.byte_transmit_counter_0 ));
    InMux I__11840 (
            .O(N__48209),
            .I(N__48205));
    InMux I__11839 (
            .O(N__48208),
            .I(N__48202));
    LocalMux I__11838 (
            .O(N__48205),
            .I(N__48199));
    LocalMux I__11837 (
            .O(N__48202),
            .I(N__48195));
    Span4Mux_h I__11836 (
            .O(N__48199),
            .I(N__48192));
    InMux I__11835 (
            .O(N__48198),
            .I(N__48189));
    Odrv4 I__11834 (
            .O(N__48195),
            .I(\c0.data_out_7_6 ));
    Odrv4 I__11833 (
            .O(N__48192),
            .I(\c0.data_out_7_6 ));
    LocalMux I__11832 (
            .O(N__48189),
            .I(\c0.data_out_7_6 ));
    CascadeMux I__11831 (
            .O(N__48182),
            .I(N__48179));
    InMux I__11830 (
            .O(N__48179),
            .I(N__48176));
    LocalMux I__11829 (
            .O(N__48176),
            .I(\c0.n5_adj_2444 ));
    InMux I__11828 (
            .O(N__48173),
            .I(N__48170));
    LocalMux I__11827 (
            .O(N__48170),
            .I(N__48167));
    Odrv4 I__11826 (
            .O(N__48167),
            .I(\c0.n8_adj_2539 ));
    CascadeMux I__11825 (
            .O(N__48164),
            .I(N__48160));
    InMux I__11824 (
            .O(N__48163),
            .I(N__48152));
    InMux I__11823 (
            .O(N__48160),
            .I(N__48145));
    InMux I__11822 (
            .O(N__48159),
            .I(N__48140));
    InMux I__11821 (
            .O(N__48158),
            .I(N__48140));
    InMux I__11820 (
            .O(N__48157),
            .I(N__48137));
    CascadeMux I__11819 (
            .O(N__48156),
            .I(N__48130));
    InMux I__11818 (
            .O(N__48155),
            .I(N__48126));
    LocalMux I__11817 (
            .O(N__48152),
            .I(N__48123));
    InMux I__11816 (
            .O(N__48151),
            .I(N__48116));
    InMux I__11815 (
            .O(N__48150),
            .I(N__48116));
    InMux I__11814 (
            .O(N__48149),
            .I(N__48116));
    InMux I__11813 (
            .O(N__48148),
            .I(N__48113));
    LocalMux I__11812 (
            .O(N__48145),
            .I(N__48103));
    LocalMux I__11811 (
            .O(N__48140),
            .I(N__48100));
    LocalMux I__11810 (
            .O(N__48137),
            .I(N__48097));
    InMux I__11809 (
            .O(N__48136),
            .I(N__48092));
    InMux I__11808 (
            .O(N__48135),
            .I(N__48092));
    InMux I__11807 (
            .O(N__48134),
            .I(N__48089));
    InMux I__11806 (
            .O(N__48133),
            .I(N__48082));
    InMux I__11805 (
            .O(N__48130),
            .I(N__48082));
    InMux I__11804 (
            .O(N__48129),
            .I(N__48082));
    LocalMux I__11803 (
            .O(N__48126),
            .I(N__48077));
    Span4Mux_v I__11802 (
            .O(N__48123),
            .I(N__48072));
    LocalMux I__11801 (
            .O(N__48116),
            .I(N__48072));
    LocalMux I__11800 (
            .O(N__48113),
            .I(N__48069));
    InMux I__11799 (
            .O(N__48112),
            .I(N__48066));
    InMux I__11798 (
            .O(N__48111),
            .I(N__48061));
    InMux I__11797 (
            .O(N__48110),
            .I(N__48061));
    InMux I__11796 (
            .O(N__48109),
            .I(N__48056));
    InMux I__11795 (
            .O(N__48108),
            .I(N__48056));
    InMux I__11794 (
            .O(N__48107),
            .I(N__48051));
    InMux I__11793 (
            .O(N__48106),
            .I(N__48051));
    Span4Mux_v I__11792 (
            .O(N__48103),
            .I(N__48038));
    Span4Mux_h I__11791 (
            .O(N__48100),
            .I(N__48038));
    Span4Mux_v I__11790 (
            .O(N__48097),
            .I(N__48038));
    LocalMux I__11789 (
            .O(N__48092),
            .I(N__48038));
    LocalMux I__11788 (
            .O(N__48089),
            .I(N__48038));
    LocalMux I__11787 (
            .O(N__48082),
            .I(N__48038));
    InMux I__11786 (
            .O(N__48081),
            .I(N__48033));
    InMux I__11785 (
            .O(N__48080),
            .I(N__48033));
    Span4Mux_v I__11784 (
            .O(N__48077),
            .I(N__48024));
    Span4Mux_h I__11783 (
            .O(N__48072),
            .I(N__48024));
    Span4Mux_v I__11782 (
            .O(N__48069),
            .I(N__48024));
    LocalMux I__11781 (
            .O(N__48066),
            .I(N__48024));
    LocalMux I__11780 (
            .O(N__48061),
            .I(N__48021));
    LocalMux I__11779 (
            .O(N__48056),
            .I(N__48018));
    LocalMux I__11778 (
            .O(N__48051),
            .I(N__48013));
    Span4Mux_h I__11777 (
            .O(N__48038),
            .I(N__48013));
    LocalMux I__11776 (
            .O(N__48033),
            .I(N__48008));
    Span4Mux_h I__11775 (
            .O(N__48024),
            .I(N__48008));
    Odrv4 I__11774 (
            .O(N__48021),
            .I(byte_transmit_counter_2));
    Odrv12 I__11773 (
            .O(N__48018),
            .I(byte_transmit_counter_2));
    Odrv4 I__11772 (
            .O(N__48013),
            .I(byte_transmit_counter_2));
    Odrv4 I__11771 (
            .O(N__48008),
            .I(byte_transmit_counter_2));
    CascadeMux I__11770 (
            .O(N__47999),
            .I(N__47996));
    InMux I__11769 (
            .O(N__47996),
            .I(N__47993));
    LocalMux I__11768 (
            .O(N__47993),
            .I(N__47990));
    Odrv12 I__11767 (
            .O(N__47990),
            .I(\c0.n18062 ));
    InMux I__11766 (
            .O(N__47987),
            .I(N__47978));
    InMux I__11765 (
            .O(N__47986),
            .I(N__47975));
    InMux I__11764 (
            .O(N__47985),
            .I(N__47964));
    InMux I__11763 (
            .O(N__47984),
            .I(N__47961));
    InMux I__11762 (
            .O(N__47983),
            .I(N__47958));
    InMux I__11761 (
            .O(N__47982),
            .I(N__47953));
    InMux I__11760 (
            .O(N__47981),
            .I(N__47950));
    LocalMux I__11759 (
            .O(N__47978),
            .I(N__47947));
    LocalMux I__11758 (
            .O(N__47975),
            .I(N__47944));
    InMux I__11757 (
            .O(N__47974),
            .I(N__47941));
    InMux I__11756 (
            .O(N__47973),
            .I(N__47934));
    InMux I__11755 (
            .O(N__47972),
            .I(N__47934));
    InMux I__11754 (
            .O(N__47971),
            .I(N__47934));
    InMux I__11753 (
            .O(N__47970),
            .I(N__47931));
    CascadeMux I__11752 (
            .O(N__47969),
            .I(N__47927));
    InMux I__11751 (
            .O(N__47968),
            .I(N__47922));
    InMux I__11750 (
            .O(N__47967),
            .I(N__47922));
    LocalMux I__11749 (
            .O(N__47964),
            .I(N__47919));
    LocalMux I__11748 (
            .O(N__47961),
            .I(N__47916));
    LocalMux I__11747 (
            .O(N__47958),
            .I(N__47913));
    InMux I__11746 (
            .O(N__47957),
            .I(N__47908));
    InMux I__11745 (
            .O(N__47956),
            .I(N__47908));
    LocalMux I__11744 (
            .O(N__47953),
            .I(N__47903));
    LocalMux I__11743 (
            .O(N__47950),
            .I(N__47903));
    Span4Mux_h I__11742 (
            .O(N__47947),
            .I(N__47894));
    Span4Mux_v I__11741 (
            .O(N__47944),
            .I(N__47894));
    LocalMux I__11740 (
            .O(N__47941),
            .I(N__47894));
    LocalMux I__11739 (
            .O(N__47934),
            .I(N__47894));
    LocalMux I__11738 (
            .O(N__47931),
            .I(N__47891));
    InMux I__11737 (
            .O(N__47930),
            .I(N__47887));
    InMux I__11736 (
            .O(N__47927),
            .I(N__47884));
    LocalMux I__11735 (
            .O(N__47922),
            .I(N__47881));
    Span4Mux_h I__11734 (
            .O(N__47919),
            .I(N__47876));
    Span4Mux_h I__11733 (
            .O(N__47916),
            .I(N__47876));
    Span4Mux_h I__11732 (
            .O(N__47913),
            .I(N__47871));
    LocalMux I__11731 (
            .O(N__47908),
            .I(N__47871));
    Span4Mux_v I__11730 (
            .O(N__47903),
            .I(N__47864));
    Span4Mux_h I__11729 (
            .O(N__47894),
            .I(N__47864));
    Span4Mux_h I__11728 (
            .O(N__47891),
            .I(N__47864));
    InMux I__11727 (
            .O(N__47890),
            .I(N__47861));
    LocalMux I__11726 (
            .O(N__47887),
            .I(\c0.byte_transmit_counter_1 ));
    LocalMux I__11725 (
            .O(N__47884),
            .I(\c0.byte_transmit_counter_1 ));
    Odrv12 I__11724 (
            .O(N__47881),
            .I(\c0.byte_transmit_counter_1 ));
    Odrv4 I__11723 (
            .O(N__47876),
            .I(\c0.byte_transmit_counter_1 ));
    Odrv4 I__11722 (
            .O(N__47871),
            .I(\c0.byte_transmit_counter_1 ));
    Odrv4 I__11721 (
            .O(N__47864),
            .I(\c0.byte_transmit_counter_1 ));
    LocalMux I__11720 (
            .O(N__47861),
            .I(\c0.byte_transmit_counter_1 ));
    InMux I__11719 (
            .O(N__47846),
            .I(N__47843));
    LocalMux I__11718 (
            .O(N__47843),
            .I(\c0.n18063 ));
    InMux I__11717 (
            .O(N__47840),
            .I(N__47837));
    LocalMux I__11716 (
            .O(N__47837),
            .I(N__47834));
    Span4Mux_h I__11715 (
            .O(N__47834),
            .I(N__47830));
    InMux I__11714 (
            .O(N__47833),
            .I(N__47827));
    Span4Mux_h I__11713 (
            .O(N__47830),
            .I(N__47822));
    LocalMux I__11712 (
            .O(N__47827),
            .I(N__47819));
    InMux I__11711 (
            .O(N__47826),
            .I(N__47814));
    InMux I__11710 (
            .O(N__47825),
            .I(N__47814));
    Odrv4 I__11709 (
            .O(N__47822),
            .I(data_out_8_0));
    Odrv4 I__11708 (
            .O(N__47819),
            .I(data_out_8_0));
    LocalMux I__11707 (
            .O(N__47814),
            .I(data_out_8_0));
    InMux I__11706 (
            .O(N__47807),
            .I(N__47804));
    LocalMux I__11705 (
            .O(N__47804),
            .I(N__47801));
    Span4Mux_h I__11704 (
            .O(N__47801),
            .I(N__47796));
    InMux I__11703 (
            .O(N__47800),
            .I(N__47793));
    InMux I__11702 (
            .O(N__47799),
            .I(N__47790));
    Odrv4 I__11701 (
            .O(N__47796),
            .I(\c0.data_out_7_7 ));
    LocalMux I__11700 (
            .O(N__47793),
            .I(\c0.data_out_7_7 ));
    LocalMux I__11699 (
            .O(N__47790),
            .I(\c0.data_out_7_7 ));
    CascadeMux I__11698 (
            .O(N__47783),
            .I(N__47780));
    InMux I__11697 (
            .O(N__47780),
            .I(N__47774));
    InMux I__11696 (
            .O(N__47779),
            .I(N__47774));
    LocalMux I__11695 (
            .O(N__47774),
            .I(\c0.n17638 ));
    InMux I__11694 (
            .O(N__47771),
            .I(N__47763));
    InMux I__11693 (
            .O(N__47770),
            .I(N__47760));
    InMux I__11692 (
            .O(N__47769),
            .I(N__47757));
    InMux I__11691 (
            .O(N__47768),
            .I(N__47754));
    InMux I__11690 (
            .O(N__47767),
            .I(N__47750));
    InMux I__11689 (
            .O(N__47766),
            .I(N__47747));
    LocalMux I__11688 (
            .O(N__47763),
            .I(N__47744));
    LocalMux I__11687 (
            .O(N__47760),
            .I(N__47741));
    LocalMux I__11686 (
            .O(N__47757),
            .I(N__47736));
    LocalMux I__11685 (
            .O(N__47754),
            .I(N__47736));
    InMux I__11684 (
            .O(N__47753),
            .I(N__47733));
    LocalMux I__11683 (
            .O(N__47750),
            .I(N__47730));
    LocalMux I__11682 (
            .O(N__47747),
            .I(N__47723));
    Span4Mux_v I__11681 (
            .O(N__47744),
            .I(N__47723));
    Span4Mux_v I__11680 (
            .O(N__47741),
            .I(N__47723));
    Span4Mux_v I__11679 (
            .O(N__47736),
            .I(N__47720));
    LocalMux I__11678 (
            .O(N__47733),
            .I(\c0.data_out_0_6 ));
    Odrv4 I__11677 (
            .O(N__47730),
            .I(\c0.data_out_0_6 ));
    Odrv4 I__11676 (
            .O(N__47723),
            .I(\c0.data_out_0_6 ));
    Odrv4 I__11675 (
            .O(N__47720),
            .I(\c0.data_out_0_6 ));
    CascadeMux I__11674 (
            .O(N__47711),
            .I(N__47708));
    InMux I__11673 (
            .O(N__47708),
            .I(N__47705));
    LocalMux I__11672 (
            .O(N__47705),
            .I(N__47700));
    InMux I__11671 (
            .O(N__47704),
            .I(N__47697));
    InMux I__11670 (
            .O(N__47703),
            .I(N__47692));
    Span4Mux_v I__11669 (
            .O(N__47700),
            .I(N__47687));
    LocalMux I__11668 (
            .O(N__47697),
            .I(N__47687));
    InMux I__11667 (
            .O(N__47696),
            .I(N__47684));
    InMux I__11666 (
            .O(N__47695),
            .I(N__47681));
    LocalMux I__11665 (
            .O(N__47692),
            .I(N__47674));
    Span4Mux_h I__11664 (
            .O(N__47687),
            .I(N__47674));
    LocalMux I__11663 (
            .O(N__47684),
            .I(N__47674));
    LocalMux I__11662 (
            .O(N__47681),
            .I(N__47671));
    Span4Mux_v I__11661 (
            .O(N__47674),
            .I(N__47664));
    Span4Mux_h I__11660 (
            .O(N__47671),
            .I(N__47664));
    InMux I__11659 (
            .O(N__47670),
            .I(N__47661));
    InMux I__11658 (
            .O(N__47669),
            .I(N__47658));
    Span4Mux_h I__11657 (
            .O(N__47664),
            .I(N__47655));
    LocalMux I__11656 (
            .O(N__47661),
            .I(data_out_0_3));
    LocalMux I__11655 (
            .O(N__47658),
            .I(data_out_0_3));
    Odrv4 I__11654 (
            .O(N__47655),
            .I(data_out_0_3));
    InMux I__11653 (
            .O(N__47648),
            .I(N__47645));
    LocalMux I__11652 (
            .O(N__47645),
            .I(N__47641));
    InMux I__11651 (
            .O(N__47644),
            .I(N__47637));
    Span4Mux_v I__11650 (
            .O(N__47641),
            .I(N__47632));
    InMux I__11649 (
            .O(N__47640),
            .I(N__47629));
    LocalMux I__11648 (
            .O(N__47637),
            .I(N__47626));
    InMux I__11647 (
            .O(N__47636),
            .I(N__47623));
    InMux I__11646 (
            .O(N__47635),
            .I(N__47620));
    Span4Mux_h I__11645 (
            .O(N__47632),
            .I(N__47616));
    LocalMux I__11644 (
            .O(N__47629),
            .I(N__47613));
    Span4Mux_v I__11643 (
            .O(N__47626),
            .I(N__47610));
    LocalMux I__11642 (
            .O(N__47623),
            .I(N__47605));
    LocalMux I__11641 (
            .O(N__47620),
            .I(N__47605));
    InMux I__11640 (
            .O(N__47619),
            .I(N__47602));
    Span4Mux_v I__11639 (
            .O(N__47616),
            .I(N__47599));
    Span4Mux_v I__11638 (
            .O(N__47613),
            .I(N__47596));
    Span4Mux_v I__11637 (
            .O(N__47610),
            .I(N__47591));
    Span4Mux_v I__11636 (
            .O(N__47605),
            .I(N__47591));
    LocalMux I__11635 (
            .O(N__47602),
            .I(N__47584));
    Span4Mux_h I__11634 (
            .O(N__47599),
            .I(N__47584));
    Span4Mux_v I__11633 (
            .O(N__47596),
            .I(N__47584));
    Odrv4 I__11632 (
            .O(N__47591),
            .I(data_out_0_1));
    Odrv4 I__11631 (
            .O(N__47584),
            .I(data_out_0_1));
    InMux I__11630 (
            .O(N__47579),
            .I(N__47574));
    InMux I__11629 (
            .O(N__47578),
            .I(N__47571));
    InMux I__11628 (
            .O(N__47577),
            .I(N__47568));
    LocalMux I__11627 (
            .O(N__47574),
            .I(N__47565));
    LocalMux I__11626 (
            .O(N__47571),
            .I(N__47562));
    LocalMux I__11625 (
            .O(N__47568),
            .I(N__47558));
    Span4Mux_s2_v I__11624 (
            .O(N__47565),
            .I(N__47553));
    Span4Mux_s2_v I__11623 (
            .O(N__47562),
            .I(N__47553));
    InMux I__11622 (
            .O(N__47561),
            .I(N__47550));
    Span4Mux_v I__11621 (
            .O(N__47558),
            .I(N__47547));
    Span4Mux_h I__11620 (
            .O(N__47553),
            .I(N__47544));
    LocalMux I__11619 (
            .O(N__47550),
            .I(data_out_0_0));
    Odrv4 I__11618 (
            .O(N__47547),
            .I(data_out_0_0));
    Odrv4 I__11617 (
            .O(N__47544),
            .I(data_out_0_0));
    CascadeMux I__11616 (
            .O(N__47537),
            .I(N__47534));
    InMux I__11615 (
            .O(N__47534),
            .I(N__47530));
    InMux I__11614 (
            .O(N__47533),
            .I(N__47526));
    LocalMux I__11613 (
            .O(N__47530),
            .I(N__47523));
    InMux I__11612 (
            .O(N__47529),
            .I(N__47520));
    LocalMux I__11611 (
            .O(N__47526),
            .I(N__47513));
    Span4Mux_s1_v I__11610 (
            .O(N__47523),
            .I(N__47513));
    LocalMux I__11609 (
            .O(N__47520),
            .I(N__47513));
    Span4Mux_v I__11608 (
            .O(N__47513),
            .I(N__47510));
    Odrv4 I__11607 (
            .O(N__47510),
            .I(\c0.n8926 ));
    InMux I__11606 (
            .O(N__47507),
            .I(N__47504));
    LocalMux I__11605 (
            .O(N__47504),
            .I(\c0.n8767 ));
    CascadeMux I__11604 (
            .O(N__47501),
            .I(\c0.n8926_cascade_ ));
    CascadeMux I__11603 (
            .O(N__47498),
            .I(N__47495));
    InMux I__11602 (
            .O(N__47495),
            .I(N__47489));
    InMux I__11601 (
            .O(N__47494),
            .I(N__47489));
    LocalMux I__11600 (
            .O(N__47489),
            .I(N__47485));
    InMux I__11599 (
            .O(N__47488),
            .I(N__47482));
    Span4Mux_h I__11598 (
            .O(N__47485),
            .I(N__47477));
    LocalMux I__11597 (
            .O(N__47482),
            .I(N__47477));
    Span4Mux_h I__11596 (
            .O(N__47477),
            .I(N__47473));
    InMux I__11595 (
            .O(N__47476),
            .I(N__47470));
    Odrv4 I__11594 (
            .O(N__47473),
            .I(n2720));
    LocalMux I__11593 (
            .O(N__47470),
            .I(n2720));
    CascadeMux I__11592 (
            .O(N__47465),
            .I(N__47462));
    InMux I__11591 (
            .O(N__47462),
            .I(N__47458));
    CascadeMux I__11590 (
            .O(N__47461),
            .I(N__47455));
    LocalMux I__11589 (
            .O(N__47458),
            .I(N__47431));
    InMux I__11588 (
            .O(N__47455),
            .I(N__47428));
    InMux I__11587 (
            .O(N__47454),
            .I(N__47421));
    InMux I__11586 (
            .O(N__47453),
            .I(N__47421));
    InMux I__11585 (
            .O(N__47452),
            .I(N__47421));
    InMux I__11584 (
            .O(N__47451),
            .I(N__47416));
    InMux I__11583 (
            .O(N__47450),
            .I(N__47416));
    CascadeMux I__11582 (
            .O(N__47449),
            .I(N__47406));
    InMux I__11581 (
            .O(N__47448),
            .I(N__47386));
    InMux I__11580 (
            .O(N__47447),
            .I(N__47386));
    InMux I__11579 (
            .O(N__47446),
            .I(N__47386));
    InMux I__11578 (
            .O(N__47445),
            .I(N__47386));
    InMux I__11577 (
            .O(N__47444),
            .I(N__47386));
    InMux I__11576 (
            .O(N__47443),
            .I(N__47375));
    InMux I__11575 (
            .O(N__47442),
            .I(N__47375));
    InMux I__11574 (
            .O(N__47441),
            .I(N__47375));
    InMux I__11573 (
            .O(N__47440),
            .I(N__47375));
    InMux I__11572 (
            .O(N__47439),
            .I(N__47375));
    InMux I__11571 (
            .O(N__47438),
            .I(N__47368));
    InMux I__11570 (
            .O(N__47437),
            .I(N__47368));
    InMux I__11569 (
            .O(N__47436),
            .I(N__47368));
    InMux I__11568 (
            .O(N__47435),
            .I(N__47363));
    InMux I__11567 (
            .O(N__47434),
            .I(N__47363));
    Span4Mux_v I__11566 (
            .O(N__47431),
            .I(N__47356));
    LocalMux I__11565 (
            .O(N__47428),
            .I(N__47356));
    LocalMux I__11564 (
            .O(N__47421),
            .I(N__47356));
    LocalMux I__11563 (
            .O(N__47416),
            .I(N__47353));
    InMux I__11562 (
            .O(N__47415),
            .I(N__47348));
    InMux I__11561 (
            .O(N__47414),
            .I(N__47348));
    InMux I__11560 (
            .O(N__47413),
            .I(N__47343));
    InMux I__11559 (
            .O(N__47412),
            .I(N__47343));
    InMux I__11558 (
            .O(N__47411),
            .I(N__47338));
    InMux I__11557 (
            .O(N__47410),
            .I(N__47333));
    InMux I__11556 (
            .O(N__47409),
            .I(N__47333));
    InMux I__11555 (
            .O(N__47406),
            .I(N__47330));
    InMux I__11554 (
            .O(N__47405),
            .I(N__47327));
    InMux I__11553 (
            .O(N__47404),
            .I(N__47322));
    InMux I__11552 (
            .O(N__47403),
            .I(N__47322));
    InMux I__11551 (
            .O(N__47402),
            .I(N__47317));
    InMux I__11550 (
            .O(N__47401),
            .I(N__47317));
    InMux I__11549 (
            .O(N__47400),
            .I(N__47312));
    InMux I__11548 (
            .O(N__47399),
            .I(N__47312));
    InMux I__11547 (
            .O(N__47398),
            .I(N__47307));
    InMux I__11546 (
            .O(N__47397),
            .I(N__47307));
    LocalMux I__11545 (
            .O(N__47386),
            .I(N__47302));
    LocalMux I__11544 (
            .O(N__47375),
            .I(N__47302));
    LocalMux I__11543 (
            .O(N__47368),
            .I(N__47284));
    LocalMux I__11542 (
            .O(N__47363),
            .I(N__47284));
    Span4Mux_s1_v I__11541 (
            .O(N__47356),
            .I(N__47284));
    Span4Mux_s1_v I__11540 (
            .O(N__47353),
            .I(N__47284));
    LocalMux I__11539 (
            .O(N__47348),
            .I(N__47284));
    LocalMux I__11538 (
            .O(N__47343),
            .I(N__47280));
    InMux I__11537 (
            .O(N__47342),
            .I(N__47277));
    InMux I__11536 (
            .O(N__47341),
            .I(N__47272));
    LocalMux I__11535 (
            .O(N__47338),
            .I(N__47259));
    LocalMux I__11534 (
            .O(N__47333),
            .I(N__47259));
    LocalMux I__11533 (
            .O(N__47330),
            .I(N__47259));
    LocalMux I__11532 (
            .O(N__47327),
            .I(N__47259));
    LocalMux I__11531 (
            .O(N__47322),
            .I(N__47259));
    LocalMux I__11530 (
            .O(N__47317),
            .I(N__47259));
    LocalMux I__11529 (
            .O(N__47312),
            .I(N__47252));
    LocalMux I__11528 (
            .O(N__47307),
            .I(N__47252));
    Span4Mux_s3_v I__11527 (
            .O(N__47302),
            .I(N__47252));
    InMux I__11526 (
            .O(N__47301),
            .I(N__47243));
    InMux I__11525 (
            .O(N__47300),
            .I(N__47243));
    InMux I__11524 (
            .O(N__47299),
            .I(N__47243));
    InMux I__11523 (
            .O(N__47298),
            .I(N__47243));
    InMux I__11522 (
            .O(N__47297),
            .I(N__47237));
    InMux I__11521 (
            .O(N__47296),
            .I(N__47230));
    InMux I__11520 (
            .O(N__47295),
            .I(N__47230));
    Span4Mux_v I__11519 (
            .O(N__47284),
            .I(N__47226));
    InMux I__11518 (
            .O(N__47283),
            .I(N__47223));
    Span4Mux_v I__11517 (
            .O(N__47280),
            .I(N__47220));
    LocalMux I__11516 (
            .O(N__47277),
            .I(N__47217));
    InMux I__11515 (
            .O(N__47276),
            .I(N__47212));
    InMux I__11514 (
            .O(N__47275),
            .I(N__47212));
    LocalMux I__11513 (
            .O(N__47272),
            .I(N__47203));
    Span4Mux_s3_v I__11512 (
            .O(N__47259),
            .I(N__47203));
    Span4Mux_h I__11511 (
            .O(N__47252),
            .I(N__47203));
    LocalMux I__11510 (
            .O(N__47243),
            .I(N__47203));
    InMux I__11509 (
            .O(N__47242),
            .I(N__47200));
    InMux I__11508 (
            .O(N__47241),
            .I(N__47197));
    InMux I__11507 (
            .O(N__47240),
            .I(N__47194));
    LocalMux I__11506 (
            .O(N__47237),
            .I(N__47191));
    InMux I__11505 (
            .O(N__47236),
            .I(N__47188));
    InMux I__11504 (
            .O(N__47235),
            .I(N__47185));
    LocalMux I__11503 (
            .O(N__47230),
            .I(N__47182));
    InMux I__11502 (
            .O(N__47229),
            .I(N__47179));
    Span4Mux_v I__11501 (
            .O(N__47226),
            .I(N__47170));
    LocalMux I__11500 (
            .O(N__47223),
            .I(N__47170));
    Span4Mux_v I__11499 (
            .O(N__47220),
            .I(N__47170));
    Span4Mux_v I__11498 (
            .O(N__47217),
            .I(N__47170));
    LocalMux I__11497 (
            .O(N__47212),
            .I(N__47163));
    Span4Mux_v I__11496 (
            .O(N__47203),
            .I(N__47163));
    LocalMux I__11495 (
            .O(N__47200),
            .I(N__47163));
    LocalMux I__11494 (
            .O(N__47197),
            .I(UART_TRANSMITTER_state_0));
    LocalMux I__11493 (
            .O(N__47194),
            .I(UART_TRANSMITTER_state_0));
    Odrv12 I__11492 (
            .O(N__47191),
            .I(UART_TRANSMITTER_state_0));
    LocalMux I__11491 (
            .O(N__47188),
            .I(UART_TRANSMITTER_state_0));
    LocalMux I__11490 (
            .O(N__47185),
            .I(UART_TRANSMITTER_state_0));
    Odrv4 I__11489 (
            .O(N__47182),
            .I(UART_TRANSMITTER_state_0));
    LocalMux I__11488 (
            .O(N__47179),
            .I(UART_TRANSMITTER_state_0));
    Odrv4 I__11487 (
            .O(N__47170),
            .I(UART_TRANSMITTER_state_0));
    Odrv4 I__11486 (
            .O(N__47163),
            .I(UART_TRANSMITTER_state_0));
    SRMux I__11485 (
            .O(N__47144),
            .I(N__47138));
    CascadeMux I__11484 (
            .O(N__47143),
            .I(N__47131));
    CascadeMux I__11483 (
            .O(N__47142),
            .I(N__47128));
    CascadeMux I__11482 (
            .O(N__47141),
            .I(N__47123));
    LocalMux I__11481 (
            .O(N__47138),
            .I(N__47119));
    InMux I__11480 (
            .O(N__47137),
            .I(N__47112));
    InMux I__11479 (
            .O(N__47136),
            .I(N__47112));
    InMux I__11478 (
            .O(N__47135),
            .I(N__47112));
    CascadeMux I__11477 (
            .O(N__47134),
            .I(N__47107));
    InMux I__11476 (
            .O(N__47131),
            .I(N__47103));
    InMux I__11475 (
            .O(N__47128),
            .I(N__47100));
    CascadeMux I__11474 (
            .O(N__47127),
            .I(N__47097));
    InMux I__11473 (
            .O(N__47126),
            .I(N__47094));
    InMux I__11472 (
            .O(N__47123),
            .I(N__47089));
    InMux I__11471 (
            .O(N__47122),
            .I(N__47089));
    Span4Mux_h I__11470 (
            .O(N__47119),
            .I(N__47086));
    LocalMux I__11469 (
            .O(N__47112),
            .I(N__47083));
    CascadeMux I__11468 (
            .O(N__47111),
            .I(N__47080));
    InMux I__11467 (
            .O(N__47110),
            .I(N__47074));
    InMux I__11466 (
            .O(N__47107),
            .I(N__47071));
    InMux I__11465 (
            .O(N__47106),
            .I(N__47068));
    LocalMux I__11464 (
            .O(N__47103),
            .I(N__47065));
    LocalMux I__11463 (
            .O(N__47100),
            .I(N__47062));
    InMux I__11462 (
            .O(N__47097),
            .I(N__47059));
    LocalMux I__11461 (
            .O(N__47094),
            .I(N__47054));
    LocalMux I__11460 (
            .O(N__47089),
            .I(N__47054));
    Span4Mux_v I__11459 (
            .O(N__47086),
            .I(N__47049));
    Span4Mux_s3_v I__11458 (
            .O(N__47083),
            .I(N__47049));
    InMux I__11457 (
            .O(N__47080),
            .I(N__47044));
    InMux I__11456 (
            .O(N__47079),
            .I(N__47044));
    CascadeMux I__11455 (
            .O(N__47078),
            .I(N__47041));
    CascadeMux I__11454 (
            .O(N__47077),
            .I(N__47036));
    LocalMux I__11453 (
            .O(N__47074),
            .I(N__47033));
    LocalMux I__11452 (
            .O(N__47071),
            .I(N__47030));
    LocalMux I__11451 (
            .O(N__47068),
            .I(N__47027));
    Span4Mux_h I__11450 (
            .O(N__47065),
            .I(N__47022));
    Span4Mux_h I__11449 (
            .O(N__47062),
            .I(N__47022));
    LocalMux I__11448 (
            .O(N__47059),
            .I(N__47019));
    Span4Mux_s2_v I__11447 (
            .O(N__47054),
            .I(N__47016));
    Sp12to4 I__11446 (
            .O(N__47049),
            .I(N__47011));
    LocalMux I__11445 (
            .O(N__47044),
            .I(N__47011));
    InMux I__11444 (
            .O(N__47041),
            .I(N__47004));
    InMux I__11443 (
            .O(N__47040),
            .I(N__47004));
    InMux I__11442 (
            .O(N__47039),
            .I(N__47004));
    InMux I__11441 (
            .O(N__47036),
            .I(N__47001));
    Span4Mux_s1_v I__11440 (
            .O(N__47033),
            .I(N__46992));
    Span4Mux_h I__11439 (
            .O(N__47030),
            .I(N__46992));
    Span4Mux_h I__11438 (
            .O(N__47027),
            .I(N__46992));
    Span4Mux_v I__11437 (
            .O(N__47022),
            .I(N__46992));
    Odrv12 I__11436 (
            .O(N__47019),
            .I(n4430));
    Odrv4 I__11435 (
            .O(N__47016),
            .I(n4430));
    Odrv12 I__11434 (
            .O(N__47011),
            .I(n4430));
    LocalMux I__11433 (
            .O(N__47004),
            .I(n4430));
    LocalMux I__11432 (
            .O(N__47001),
            .I(n4430));
    Odrv4 I__11431 (
            .O(N__46992),
            .I(n4430));
    InMux I__11430 (
            .O(N__46979),
            .I(N__46973));
    InMux I__11429 (
            .O(N__46978),
            .I(N__46970));
    InMux I__11428 (
            .O(N__46977),
            .I(N__46965));
    InMux I__11427 (
            .O(N__46976),
            .I(N__46965));
    LocalMux I__11426 (
            .O(N__46973),
            .I(N__46962));
    LocalMux I__11425 (
            .O(N__46970),
            .I(data_out_1_6));
    LocalMux I__11424 (
            .O(N__46965),
            .I(data_out_1_6));
    Odrv12 I__11423 (
            .O(N__46962),
            .I(data_out_1_6));
    InMux I__11422 (
            .O(N__46955),
            .I(N__46951));
    InMux I__11421 (
            .O(N__46954),
            .I(N__46946));
    LocalMux I__11420 (
            .O(N__46951),
            .I(N__46943));
    InMux I__11419 (
            .O(N__46950),
            .I(N__46940));
    InMux I__11418 (
            .O(N__46949),
            .I(N__46937));
    LocalMux I__11417 (
            .O(N__46946),
            .I(N__46934));
    Span4Mux_h I__11416 (
            .O(N__46943),
            .I(N__46931));
    LocalMux I__11415 (
            .O(N__46940),
            .I(N__46928));
    LocalMux I__11414 (
            .O(N__46937),
            .I(data_out_3_5));
    Odrv4 I__11413 (
            .O(N__46934),
            .I(data_out_3_5));
    Odrv4 I__11412 (
            .O(N__46931),
            .I(data_out_3_5));
    Odrv4 I__11411 (
            .O(N__46928),
            .I(data_out_3_5));
    CascadeMux I__11410 (
            .O(N__46919),
            .I(N__46911));
    CascadeMux I__11409 (
            .O(N__46918),
            .I(N__46908));
    CascadeMux I__11408 (
            .O(N__46917),
            .I(N__46904));
    CascadeMux I__11407 (
            .O(N__46916),
            .I(N__46885));
    CascadeMux I__11406 (
            .O(N__46915),
            .I(N__46874));
    InMux I__11405 (
            .O(N__46914),
            .I(N__46866));
    InMux I__11404 (
            .O(N__46911),
            .I(N__46863));
    InMux I__11403 (
            .O(N__46908),
            .I(N__46858));
    InMux I__11402 (
            .O(N__46907),
            .I(N__46858));
    InMux I__11401 (
            .O(N__46904),
            .I(N__46855));
    InMux I__11400 (
            .O(N__46903),
            .I(N__46848));
    InMux I__11399 (
            .O(N__46902),
            .I(N__46848));
    InMux I__11398 (
            .O(N__46901),
            .I(N__46848));
    InMux I__11397 (
            .O(N__46900),
            .I(N__46845));
    InMux I__11396 (
            .O(N__46899),
            .I(N__46842));
    InMux I__11395 (
            .O(N__46898),
            .I(N__46837));
    InMux I__11394 (
            .O(N__46897),
            .I(N__46837));
    InMux I__11393 (
            .O(N__46896),
            .I(N__46830));
    InMux I__11392 (
            .O(N__46895),
            .I(N__46830));
    InMux I__11391 (
            .O(N__46894),
            .I(N__46830));
    InMux I__11390 (
            .O(N__46893),
            .I(N__46825));
    InMux I__11389 (
            .O(N__46892),
            .I(N__46825));
    InMux I__11388 (
            .O(N__46891),
            .I(N__46820));
    InMux I__11387 (
            .O(N__46890),
            .I(N__46820));
    InMux I__11386 (
            .O(N__46889),
            .I(N__46815));
    InMux I__11385 (
            .O(N__46888),
            .I(N__46815));
    InMux I__11384 (
            .O(N__46885),
            .I(N__46812));
    InMux I__11383 (
            .O(N__46884),
            .I(N__46805));
    InMux I__11382 (
            .O(N__46883),
            .I(N__46805));
    InMux I__11381 (
            .O(N__46882),
            .I(N__46805));
    CascadeMux I__11380 (
            .O(N__46881),
            .I(N__46801));
    InMux I__11379 (
            .O(N__46880),
            .I(N__46796));
    CascadeMux I__11378 (
            .O(N__46879),
            .I(N__46790));
    InMux I__11377 (
            .O(N__46878),
            .I(N__46780));
    InMux I__11376 (
            .O(N__46877),
            .I(N__46780));
    InMux I__11375 (
            .O(N__46874),
            .I(N__46773));
    InMux I__11374 (
            .O(N__46873),
            .I(N__46773));
    InMux I__11373 (
            .O(N__46872),
            .I(N__46773));
    InMux I__11372 (
            .O(N__46871),
            .I(N__46766));
    InMux I__11371 (
            .O(N__46870),
            .I(N__46766));
    InMux I__11370 (
            .O(N__46869),
            .I(N__46766));
    LocalMux I__11369 (
            .O(N__46866),
            .I(N__46759));
    LocalMux I__11368 (
            .O(N__46863),
            .I(N__46759));
    LocalMux I__11367 (
            .O(N__46858),
            .I(N__46759));
    LocalMux I__11366 (
            .O(N__46855),
            .I(N__46756));
    LocalMux I__11365 (
            .O(N__46848),
            .I(N__46753));
    LocalMux I__11364 (
            .O(N__46845),
            .I(N__46744));
    LocalMux I__11363 (
            .O(N__46842),
            .I(N__46744));
    LocalMux I__11362 (
            .O(N__46837),
            .I(N__46744));
    LocalMux I__11361 (
            .O(N__46830),
            .I(N__46744));
    LocalMux I__11360 (
            .O(N__46825),
            .I(N__46733));
    LocalMux I__11359 (
            .O(N__46820),
            .I(N__46733));
    LocalMux I__11358 (
            .O(N__46815),
            .I(N__46733));
    LocalMux I__11357 (
            .O(N__46812),
            .I(N__46733));
    LocalMux I__11356 (
            .O(N__46805),
            .I(N__46733));
    InMux I__11355 (
            .O(N__46804),
            .I(N__46730));
    InMux I__11354 (
            .O(N__46801),
            .I(N__46725));
    InMux I__11353 (
            .O(N__46800),
            .I(N__46725));
    InMux I__11352 (
            .O(N__46799),
            .I(N__46720));
    LocalMux I__11351 (
            .O(N__46796),
            .I(N__46717));
    InMux I__11350 (
            .O(N__46795),
            .I(N__46714));
    InMux I__11349 (
            .O(N__46794),
            .I(N__46711));
    InMux I__11348 (
            .O(N__46793),
            .I(N__46706));
    InMux I__11347 (
            .O(N__46790),
            .I(N__46706));
    InMux I__11346 (
            .O(N__46789),
            .I(N__46703));
    InMux I__11345 (
            .O(N__46788),
            .I(N__46698));
    InMux I__11344 (
            .O(N__46787),
            .I(N__46698));
    InMux I__11343 (
            .O(N__46786),
            .I(N__46691));
    InMux I__11342 (
            .O(N__46785),
            .I(N__46688));
    LocalMux I__11341 (
            .O(N__46780),
            .I(N__46673));
    LocalMux I__11340 (
            .O(N__46773),
            .I(N__46673));
    LocalMux I__11339 (
            .O(N__46766),
            .I(N__46673));
    Span4Mux_s2_v I__11338 (
            .O(N__46759),
            .I(N__46673));
    Span4Mux_h I__11337 (
            .O(N__46756),
            .I(N__46673));
    Span4Mux_h I__11336 (
            .O(N__46753),
            .I(N__46673));
    Span4Mux_s2_v I__11335 (
            .O(N__46744),
            .I(N__46673));
    Span4Mux_s3_v I__11334 (
            .O(N__46733),
            .I(N__46667));
    LocalMux I__11333 (
            .O(N__46730),
            .I(N__46662));
    LocalMux I__11332 (
            .O(N__46725),
            .I(N__46662));
    InMux I__11331 (
            .O(N__46724),
            .I(N__46657));
    InMux I__11330 (
            .O(N__46723),
            .I(N__46657));
    LocalMux I__11329 (
            .O(N__46720),
            .I(N__46654));
    Span4Mux_v I__11328 (
            .O(N__46717),
            .I(N__46647));
    LocalMux I__11327 (
            .O(N__46714),
            .I(N__46647));
    LocalMux I__11326 (
            .O(N__46711),
            .I(N__46647));
    LocalMux I__11325 (
            .O(N__46706),
            .I(N__46642));
    LocalMux I__11324 (
            .O(N__46703),
            .I(N__46637));
    LocalMux I__11323 (
            .O(N__46698),
            .I(N__46637));
    InMux I__11322 (
            .O(N__46697),
            .I(N__46628));
    InMux I__11321 (
            .O(N__46696),
            .I(N__46628));
    InMux I__11320 (
            .O(N__46695),
            .I(N__46628));
    InMux I__11319 (
            .O(N__46694),
            .I(N__46628));
    LocalMux I__11318 (
            .O(N__46691),
            .I(N__46624));
    LocalMux I__11317 (
            .O(N__46688),
            .I(N__46621));
    Span4Mux_v I__11316 (
            .O(N__46673),
            .I(N__46618));
    InMux I__11315 (
            .O(N__46672),
            .I(N__46611));
    InMux I__11314 (
            .O(N__46671),
            .I(N__46611));
    InMux I__11313 (
            .O(N__46670),
            .I(N__46611));
    Span4Mux_h I__11312 (
            .O(N__46667),
            .I(N__46606));
    Span4Mux_s3_v I__11311 (
            .O(N__46662),
            .I(N__46606));
    LocalMux I__11310 (
            .O(N__46657),
            .I(N__46599));
    Span4Mux_v I__11309 (
            .O(N__46654),
            .I(N__46599));
    Span4Mux_h I__11308 (
            .O(N__46647),
            .I(N__46599));
    InMux I__11307 (
            .O(N__46646),
            .I(N__46594));
    InMux I__11306 (
            .O(N__46645),
            .I(N__46594));
    Span4Mux_h I__11305 (
            .O(N__46642),
            .I(N__46587));
    Span4Mux_v I__11304 (
            .O(N__46637),
            .I(N__46587));
    LocalMux I__11303 (
            .O(N__46628),
            .I(N__46587));
    InMux I__11302 (
            .O(N__46627),
            .I(N__46584));
    Odrv12 I__11301 (
            .O(N__46624),
            .I(UART_TRANSMITTER_state_1));
    Odrv12 I__11300 (
            .O(N__46621),
            .I(UART_TRANSMITTER_state_1));
    Odrv4 I__11299 (
            .O(N__46618),
            .I(UART_TRANSMITTER_state_1));
    LocalMux I__11298 (
            .O(N__46611),
            .I(UART_TRANSMITTER_state_1));
    Odrv4 I__11297 (
            .O(N__46606),
            .I(UART_TRANSMITTER_state_1));
    Odrv4 I__11296 (
            .O(N__46599),
            .I(UART_TRANSMITTER_state_1));
    LocalMux I__11295 (
            .O(N__46594),
            .I(UART_TRANSMITTER_state_1));
    Odrv4 I__11294 (
            .O(N__46587),
            .I(UART_TRANSMITTER_state_1));
    LocalMux I__11293 (
            .O(N__46584),
            .I(UART_TRANSMITTER_state_1));
    CEMux I__11292 (
            .O(N__46565),
            .I(N__46561));
    CEMux I__11291 (
            .O(N__46564),
            .I(N__46558));
    LocalMux I__11290 (
            .O(N__46561),
            .I(N__46554));
    LocalMux I__11289 (
            .O(N__46558),
            .I(N__46551));
    CEMux I__11288 (
            .O(N__46557),
            .I(N__46548));
    Span4Mux_s1_v I__11287 (
            .O(N__46554),
            .I(N__46539));
    Span4Mux_h I__11286 (
            .O(N__46551),
            .I(N__46539));
    LocalMux I__11285 (
            .O(N__46548),
            .I(N__46539));
    CEMux I__11284 (
            .O(N__46547),
            .I(N__46535));
    CEMux I__11283 (
            .O(N__46546),
            .I(N__46532));
    Span4Mux_h I__11282 (
            .O(N__46539),
            .I(N__46528));
    CEMux I__11281 (
            .O(N__46538),
            .I(N__46525));
    LocalMux I__11280 (
            .O(N__46535),
            .I(N__46520));
    LocalMux I__11279 (
            .O(N__46532),
            .I(N__46517));
    InMux I__11278 (
            .O(N__46531),
            .I(N__46513));
    Span4Mux_h I__11277 (
            .O(N__46528),
            .I(N__46508));
    LocalMux I__11276 (
            .O(N__46525),
            .I(N__46508));
    InMux I__11275 (
            .O(N__46524),
            .I(N__46503));
    InMux I__11274 (
            .O(N__46523),
            .I(N__46503));
    Span4Mux_v I__11273 (
            .O(N__46520),
            .I(N__46499));
    Span4Mux_v I__11272 (
            .O(N__46517),
            .I(N__46496));
    CEMux I__11271 (
            .O(N__46516),
            .I(N__46493));
    LocalMux I__11270 (
            .O(N__46513),
            .I(N__46490));
    Span4Mux_h I__11269 (
            .O(N__46508),
            .I(N__46485));
    LocalMux I__11268 (
            .O(N__46503),
            .I(N__46485));
    CascadeMux I__11267 (
            .O(N__46502),
            .I(N__46481));
    Span4Mux_h I__11266 (
            .O(N__46499),
            .I(N__46478));
    Sp12to4 I__11265 (
            .O(N__46496),
            .I(N__46475));
    LocalMux I__11264 (
            .O(N__46493),
            .I(N__46472));
    Span4Mux_h I__11263 (
            .O(N__46490),
            .I(N__46467));
    Span4Mux_s1_v I__11262 (
            .O(N__46485),
            .I(N__46467));
    InMux I__11261 (
            .O(N__46484),
            .I(N__46462));
    InMux I__11260 (
            .O(N__46481),
            .I(N__46462));
    Odrv4 I__11259 (
            .O(N__46478),
            .I(n9519));
    Odrv12 I__11258 (
            .O(N__46475),
            .I(n9519));
    Odrv4 I__11257 (
            .O(N__46472),
            .I(n9519));
    Odrv4 I__11256 (
            .O(N__46467),
            .I(n9519));
    LocalMux I__11255 (
            .O(N__46462),
            .I(n9519));
    InMux I__11254 (
            .O(N__46451),
            .I(N__46442));
    InMux I__11253 (
            .O(N__46450),
            .I(N__46442));
    InMux I__11252 (
            .O(N__46449),
            .I(N__46435));
    InMux I__11251 (
            .O(N__46448),
            .I(N__46435));
    InMux I__11250 (
            .O(N__46447),
            .I(N__46432));
    LocalMux I__11249 (
            .O(N__46442),
            .I(N__46429));
    InMux I__11248 (
            .O(N__46441),
            .I(N__46426));
    InMux I__11247 (
            .O(N__46440),
            .I(N__46423));
    LocalMux I__11246 (
            .O(N__46435),
            .I(N__46416));
    LocalMux I__11245 (
            .O(N__46432),
            .I(N__46416));
    Span4Mux_s2_v I__11244 (
            .O(N__46429),
            .I(N__46416));
    LocalMux I__11243 (
            .O(N__46426),
            .I(N__46413));
    LocalMux I__11242 (
            .O(N__46423),
            .I(N__46409));
    Span4Mux_h I__11241 (
            .O(N__46416),
            .I(N__46406));
    Span4Mux_h I__11240 (
            .O(N__46413),
            .I(N__46403));
    InMux I__11239 (
            .O(N__46412),
            .I(N__46400));
    Span12Mux_h I__11238 (
            .O(N__46409),
            .I(N__46397));
    Span4Mux_v I__11237 (
            .O(N__46406),
            .I(N__46394));
    Span4Mux_v I__11236 (
            .O(N__46403),
            .I(N__46391));
    LocalMux I__11235 (
            .O(N__46400),
            .I(data_out_5__7__N_931));
    Odrv12 I__11234 (
            .O(N__46397),
            .I(data_out_5__7__N_931));
    Odrv4 I__11233 (
            .O(N__46394),
            .I(data_out_5__7__N_931));
    Odrv4 I__11232 (
            .O(N__46391),
            .I(data_out_5__7__N_931));
    InMux I__11231 (
            .O(N__46382),
            .I(N__46379));
    LocalMux I__11230 (
            .O(N__46379),
            .I(N__46375));
    InMux I__11229 (
            .O(N__46378),
            .I(N__46372));
    Odrv4 I__11228 (
            .O(N__46375),
            .I(\c0.data_out_6__4__N_765 ));
    LocalMux I__11227 (
            .O(N__46372),
            .I(\c0.data_out_6__4__N_765 ));
    InMux I__11226 (
            .O(N__46367),
            .I(N__46361));
    InMux I__11225 (
            .O(N__46366),
            .I(N__46358));
    CascadeMux I__11224 (
            .O(N__46365),
            .I(N__46355));
    InMux I__11223 (
            .O(N__46364),
            .I(N__46352));
    LocalMux I__11222 (
            .O(N__46361),
            .I(N__46349));
    LocalMux I__11221 (
            .O(N__46358),
            .I(N__46346));
    InMux I__11220 (
            .O(N__46355),
            .I(N__46343));
    LocalMux I__11219 (
            .O(N__46352),
            .I(N__46340));
    Span4Mux_h I__11218 (
            .O(N__46349),
            .I(N__46335));
    Span4Mux_h I__11217 (
            .O(N__46346),
            .I(N__46335));
    LocalMux I__11216 (
            .O(N__46343),
            .I(\c0.data_out_7_2 ));
    Odrv12 I__11215 (
            .O(N__46340),
            .I(\c0.data_out_7_2 ));
    Odrv4 I__11214 (
            .O(N__46335),
            .I(\c0.data_out_7_2 ));
    CascadeMux I__11213 (
            .O(N__46328),
            .I(N__46325));
    InMux I__11212 (
            .O(N__46325),
            .I(N__46322));
    LocalMux I__11211 (
            .O(N__46322),
            .I(N__46319));
    Odrv12 I__11210 (
            .O(N__46319),
            .I(\c0.n17600 ));
    InMux I__11209 (
            .O(N__46316),
            .I(N__46313));
    LocalMux I__11208 (
            .O(N__46313),
            .I(\c0.data_out_9_6 ));
    InMux I__11207 (
            .O(N__46310),
            .I(N__46306));
    InMux I__11206 (
            .O(N__46309),
            .I(N__46303));
    LocalMux I__11205 (
            .O(N__46306),
            .I(N__46297));
    LocalMux I__11204 (
            .O(N__46303),
            .I(N__46297));
    InMux I__11203 (
            .O(N__46302),
            .I(N__46294));
    Span4Mux_h I__11202 (
            .O(N__46297),
            .I(N__46291));
    LocalMux I__11201 (
            .O(N__46294),
            .I(\c0.data_out_7_1 ));
    Odrv4 I__11200 (
            .O(N__46291),
            .I(\c0.data_out_7_1 ));
    InMux I__11199 (
            .O(N__46286),
            .I(N__46283));
    LocalMux I__11198 (
            .O(N__46283),
            .I(\c0.n17454 ));
    InMux I__11197 (
            .O(N__46280),
            .I(N__46276));
    InMux I__11196 (
            .O(N__46279),
            .I(N__46272));
    LocalMux I__11195 (
            .O(N__46276),
            .I(N__46269));
    InMux I__11194 (
            .O(N__46275),
            .I(N__46266));
    LocalMux I__11193 (
            .O(N__46272),
            .I(N__46261));
    Span4Mux_h I__11192 (
            .O(N__46269),
            .I(N__46261));
    LocalMux I__11191 (
            .O(N__46266),
            .I(\c0.data_out_6_5 ));
    Odrv4 I__11190 (
            .O(N__46261),
            .I(\c0.data_out_6_5 ));
    InMux I__11189 (
            .O(N__46256),
            .I(N__46252));
    InMux I__11188 (
            .O(N__46255),
            .I(N__46249));
    LocalMux I__11187 (
            .O(N__46252),
            .I(\c0.data_out_6__5__N_752 ));
    LocalMux I__11186 (
            .O(N__46249),
            .I(\c0.data_out_6__5__N_752 ));
    CascadeMux I__11185 (
            .O(N__46244),
            .I(\c0.n17454_cascade_ ));
    InMux I__11184 (
            .O(N__46241),
            .I(N__46238));
    LocalMux I__11183 (
            .O(N__46238),
            .I(\c0.data_out_9_5 ));
    InMux I__11182 (
            .O(N__46235),
            .I(N__46232));
    LocalMux I__11181 (
            .O(N__46232),
            .I(N__46229));
    Span4Mux_h I__11180 (
            .O(N__46229),
            .I(N__46226));
    Odrv4 I__11179 (
            .O(N__46226),
            .I(\c0.n8_adj_2537 ));
    InMux I__11178 (
            .O(N__46223),
            .I(N__46220));
    LocalMux I__11177 (
            .O(N__46220),
            .I(N__46216));
    CascadeMux I__11176 (
            .O(N__46219),
            .I(N__46213));
    Span4Mux_s3_v I__11175 (
            .O(N__46216),
            .I(N__46210));
    InMux I__11174 (
            .O(N__46213),
            .I(N__46207));
    Span4Mux_h I__11173 (
            .O(N__46210),
            .I(N__46204));
    LocalMux I__11172 (
            .O(N__46207),
            .I(\c0.n17626 ));
    Odrv4 I__11171 (
            .O(N__46204),
            .I(\c0.n17626 ));
    InMux I__11170 (
            .O(N__46199),
            .I(N__46195));
    InMux I__11169 (
            .O(N__46198),
            .I(N__46192));
    LocalMux I__11168 (
            .O(N__46195),
            .I(N__46189));
    LocalMux I__11167 (
            .O(N__46192),
            .I(\c0.n17608 ));
    Odrv4 I__11166 (
            .O(N__46189),
            .I(\c0.n17608 ));
    CascadeMux I__11165 (
            .O(N__46184),
            .I(N__46180));
    InMux I__11164 (
            .O(N__46183),
            .I(N__46177));
    InMux I__11163 (
            .O(N__46180),
            .I(N__46174));
    LocalMux I__11162 (
            .O(N__46177),
            .I(N__46169));
    LocalMux I__11161 (
            .O(N__46174),
            .I(N__46169));
    Span4Mux_h I__11160 (
            .O(N__46169),
            .I(N__46166));
    Odrv4 I__11159 (
            .O(N__46166),
            .I(\c0.n8970 ));
    InMux I__11158 (
            .O(N__46163),
            .I(N__46160));
    LocalMux I__11157 (
            .O(N__46160),
            .I(N__46157));
    Span4Mux_h I__11156 (
            .O(N__46157),
            .I(N__46154));
    Odrv4 I__11155 (
            .O(N__46154),
            .I(\c0.n17662 ));
    InMux I__11154 (
            .O(N__46151),
            .I(N__46143));
    InMux I__11153 (
            .O(N__46150),
            .I(N__46143));
    InMux I__11152 (
            .O(N__46149),
            .I(N__46138));
    InMux I__11151 (
            .O(N__46148),
            .I(N__46138));
    LocalMux I__11150 (
            .O(N__46143),
            .I(N__46135));
    LocalMux I__11149 (
            .O(N__46138),
            .I(N__46131));
    Span4Mux_h I__11148 (
            .O(N__46135),
            .I(N__46128));
    InMux I__11147 (
            .O(N__46134),
            .I(N__46125));
    Span4Mux_v I__11146 (
            .O(N__46131),
            .I(N__46122));
    Span4Mux_h I__11145 (
            .O(N__46128),
            .I(N__46119));
    LocalMux I__11144 (
            .O(N__46125),
            .I(data_out_8_6));
    Odrv4 I__11143 (
            .O(N__46122),
            .I(data_out_8_6));
    Odrv4 I__11142 (
            .O(N__46119),
            .I(data_out_8_6));
    InMux I__11141 (
            .O(N__46112),
            .I(N__46109));
    LocalMux I__11140 (
            .O(N__46109),
            .I(N__46106));
    Span4Mux_v I__11139 (
            .O(N__46106),
            .I(N__46102));
    InMux I__11138 (
            .O(N__46105),
            .I(N__46099));
    Sp12to4 I__11137 (
            .O(N__46102),
            .I(N__46094));
    LocalMux I__11136 (
            .O(N__46099),
            .I(N__46094));
    Odrv12 I__11135 (
            .O(N__46094),
            .I(\c0.n17665 ));
    CascadeMux I__11134 (
            .O(N__46091),
            .I(\c0.n12_adj_2482_cascade_ ));
    InMux I__11133 (
            .O(N__46088),
            .I(N__46083));
    InMux I__11132 (
            .O(N__46087),
            .I(N__46080));
    InMux I__11131 (
            .O(N__46086),
            .I(N__46076));
    LocalMux I__11130 (
            .O(N__46083),
            .I(N__46073));
    LocalMux I__11129 (
            .O(N__46080),
            .I(N__46070));
    InMux I__11128 (
            .O(N__46079),
            .I(N__46067));
    LocalMux I__11127 (
            .O(N__46076),
            .I(N__46064));
    Span4Mux_h I__11126 (
            .O(N__46073),
            .I(N__46057));
    Span4Mux_v I__11125 (
            .O(N__46070),
            .I(N__46057));
    LocalMux I__11124 (
            .O(N__46067),
            .I(N__46057));
    Span4Mux_h I__11123 (
            .O(N__46064),
            .I(N__46054));
    Odrv4 I__11122 (
            .O(N__46057),
            .I(\c0.data_out_7_3 ));
    Odrv4 I__11121 (
            .O(N__46054),
            .I(\c0.data_out_7_3 ));
    InMux I__11120 (
            .O(N__46049),
            .I(N__46042));
    InMux I__11119 (
            .O(N__46048),
            .I(N__46042));
    CEMux I__11118 (
            .O(N__46047),
            .I(N__46038));
    LocalMux I__11117 (
            .O(N__46042),
            .I(N__46026));
    InMux I__11116 (
            .O(N__46041),
            .I(N__46023));
    LocalMux I__11115 (
            .O(N__46038),
            .I(N__46019));
    CEMux I__11114 (
            .O(N__46037),
            .I(N__46016));
    CEMux I__11113 (
            .O(N__46036),
            .I(N__46012));
    CEMux I__11112 (
            .O(N__46035),
            .I(N__46009));
    CEMux I__11111 (
            .O(N__46034),
            .I(N__46005));
    InMux I__11110 (
            .O(N__46033),
            .I(N__46002));
    InMux I__11109 (
            .O(N__46032),
            .I(N__45995));
    InMux I__11108 (
            .O(N__46031),
            .I(N__45995));
    InMux I__11107 (
            .O(N__46030),
            .I(N__45995));
    CEMux I__11106 (
            .O(N__46029),
            .I(N__45992));
    Span4Mux_h I__11105 (
            .O(N__46026),
            .I(N__45987));
    LocalMux I__11104 (
            .O(N__46023),
            .I(N__45987));
    InMux I__11103 (
            .O(N__46022),
            .I(N__45984));
    Span4Mux_h I__11102 (
            .O(N__46019),
            .I(N__45981));
    LocalMux I__11101 (
            .O(N__46016),
            .I(N__45978));
    CEMux I__11100 (
            .O(N__46015),
            .I(N__45975));
    LocalMux I__11099 (
            .O(N__46012),
            .I(N__45970));
    LocalMux I__11098 (
            .O(N__46009),
            .I(N__45970));
    CEMux I__11097 (
            .O(N__46008),
            .I(N__45967));
    LocalMux I__11096 (
            .O(N__46005),
            .I(N__45964));
    LocalMux I__11095 (
            .O(N__46002),
            .I(N__45959));
    LocalMux I__11094 (
            .O(N__45995),
            .I(N__45959));
    LocalMux I__11093 (
            .O(N__45992),
            .I(N__45952));
    Span4Mux_h I__11092 (
            .O(N__45987),
            .I(N__45952));
    LocalMux I__11091 (
            .O(N__45984),
            .I(N__45952));
    Span4Mux_v I__11090 (
            .O(N__45981),
            .I(N__45949));
    Span4Mux_v I__11089 (
            .O(N__45978),
            .I(N__45942));
    LocalMux I__11088 (
            .O(N__45975),
            .I(N__45942));
    Span4Mux_v I__11087 (
            .O(N__45970),
            .I(N__45942));
    LocalMux I__11086 (
            .O(N__45967),
            .I(N__45939));
    Span4Mux_h I__11085 (
            .O(N__45964),
            .I(N__45934));
    Span4Mux_v I__11084 (
            .O(N__45959),
            .I(N__45934));
    Span4Mux_v I__11083 (
            .O(N__45952),
            .I(N__45931));
    Odrv4 I__11082 (
            .O(N__45949),
            .I(data_out_10__7__N_114));
    Odrv4 I__11081 (
            .O(N__45942),
            .I(data_out_10__7__N_114));
    Odrv12 I__11080 (
            .O(N__45939),
            .I(data_out_10__7__N_114));
    Odrv4 I__11079 (
            .O(N__45934),
            .I(data_out_10__7__N_114));
    Odrv4 I__11078 (
            .O(N__45931),
            .I(data_out_10__7__N_114));
    InMux I__11077 (
            .O(N__45920),
            .I(N__45917));
    LocalMux I__11076 (
            .O(N__45917),
            .I(\c0.data_out_9_7 ));
    InMux I__11075 (
            .O(N__45914),
            .I(N__45908));
    InMux I__11074 (
            .O(N__45913),
            .I(N__45905));
    InMux I__11073 (
            .O(N__45912),
            .I(N__45900));
    InMux I__11072 (
            .O(N__45911),
            .I(N__45900));
    LocalMux I__11071 (
            .O(N__45908),
            .I(N__45896));
    LocalMux I__11070 (
            .O(N__45905),
            .I(N__45891));
    LocalMux I__11069 (
            .O(N__45900),
            .I(N__45891));
    InMux I__11068 (
            .O(N__45899),
            .I(N__45888));
    Span4Mux_v I__11067 (
            .O(N__45896),
            .I(N__45883));
    Span4Mux_v I__11066 (
            .O(N__45891),
            .I(N__45883));
    LocalMux I__11065 (
            .O(N__45888),
            .I(N__45878));
    Span4Mux_h I__11064 (
            .O(N__45883),
            .I(N__45878));
    Odrv4 I__11063 (
            .O(N__45878),
            .I(data_out_8_7));
    InMux I__11062 (
            .O(N__45875),
            .I(N__45872));
    LocalMux I__11061 (
            .O(N__45872),
            .I(N__45869));
    Span12Mux_v I__11060 (
            .O(N__45869),
            .I(N__45866));
    Odrv12 I__11059 (
            .O(N__45866),
            .I(\c0.n8_adj_2538 ));
    InMux I__11058 (
            .O(N__45863),
            .I(N__45860));
    LocalMux I__11057 (
            .O(N__45860),
            .I(\c0.data_out_10_5 ));
    CascadeMux I__11056 (
            .O(N__45857),
            .I(N__45854));
    InMux I__11055 (
            .O(N__45854),
            .I(N__45851));
    LocalMux I__11054 (
            .O(N__45851),
            .I(N__45848));
    Odrv4 I__11053 (
            .O(N__45848),
            .I(\c0.n18064 ));
    InMux I__11052 (
            .O(N__45845),
            .I(N__45842));
    LocalMux I__11051 (
            .O(N__45842),
            .I(\c0.n17668 ));
    CascadeMux I__11050 (
            .O(N__45839),
            .I(N__45835));
    InMux I__11049 (
            .O(N__45838),
            .I(N__45831));
    InMux I__11048 (
            .O(N__45835),
            .I(N__45828));
    InMux I__11047 (
            .O(N__45834),
            .I(N__45825));
    LocalMux I__11046 (
            .O(N__45831),
            .I(N__45820));
    LocalMux I__11045 (
            .O(N__45828),
            .I(N__45820));
    LocalMux I__11044 (
            .O(N__45825),
            .I(N__45817));
    Span4Mux_v I__11043 (
            .O(N__45820),
            .I(N__45814));
    Span4Mux_v I__11042 (
            .O(N__45817),
            .I(N__45811));
    Span4Mux_h I__11041 (
            .O(N__45814),
            .I(N__45808));
    Odrv4 I__11040 (
            .O(N__45811),
            .I(\c0.n9087 ));
    Odrv4 I__11039 (
            .O(N__45808),
            .I(\c0.n9087 ));
    CascadeMux I__11038 (
            .O(N__45803),
            .I(\c0.n8_adj_2528_cascade_ ));
    InMux I__11037 (
            .O(N__45800),
            .I(N__45797));
    LocalMux I__11036 (
            .O(N__45797),
            .I(\c0.data_out_10_1 ));
    InMux I__11035 (
            .O(N__45794),
            .I(N__45791));
    LocalMux I__11034 (
            .O(N__45791),
            .I(N__45788));
    Span4Mux_v I__11033 (
            .O(N__45788),
            .I(N__45785));
    Span4Mux_h I__11032 (
            .O(N__45785),
            .I(N__45782));
    Odrv4 I__11031 (
            .O(N__45782),
            .I(\c0.n17556 ));
    InMux I__11030 (
            .O(N__45779),
            .I(N__45775));
    InMux I__11029 (
            .O(N__45778),
            .I(N__45772));
    LocalMux I__11028 (
            .O(N__45775),
            .I(N__45769));
    LocalMux I__11027 (
            .O(N__45772),
            .I(N__45766));
    Span4Mux_s2_v I__11026 (
            .O(N__45769),
            .I(N__45763));
    Odrv4 I__11025 (
            .O(N__45766),
            .I(\c0.data_out_6__7__N_675 ));
    Odrv4 I__11024 (
            .O(N__45763),
            .I(\c0.data_out_6__7__N_675 ));
    InMux I__11023 (
            .O(N__45758),
            .I(N__45755));
    LocalMux I__11022 (
            .O(N__45755),
            .I(N__45752));
    Odrv12 I__11021 (
            .O(N__45752),
            .I(\c0.data_out_10_7 ));
    InMux I__11020 (
            .O(N__45749),
            .I(N__45746));
    LocalMux I__11019 (
            .O(N__45746),
            .I(N__45742));
    InMux I__11018 (
            .O(N__45745),
            .I(N__45739));
    Span4Mux_v I__11017 (
            .O(N__45742),
            .I(N__45736));
    LocalMux I__11016 (
            .O(N__45739),
            .I(N__45733));
    Sp12to4 I__11015 (
            .O(N__45736),
            .I(N__45728));
    Span12Mux_s5_v I__11014 (
            .O(N__45733),
            .I(N__45728));
    Span12Mux_h I__11013 (
            .O(N__45728),
            .I(N__45725));
    Odrv12 I__11012 (
            .O(N__45725),
            .I(\c0.n8600 ));
    InMux I__11011 (
            .O(N__45722),
            .I(N__45718));
    InMux I__11010 (
            .O(N__45721),
            .I(N__45714));
    LocalMux I__11009 (
            .O(N__45718),
            .I(N__45710));
    InMux I__11008 (
            .O(N__45717),
            .I(N__45707));
    LocalMux I__11007 (
            .O(N__45714),
            .I(N__45704));
    InMux I__11006 (
            .O(N__45713),
            .I(N__45701));
    Span4Mux_v I__11005 (
            .O(N__45710),
            .I(N__45696));
    LocalMux I__11004 (
            .O(N__45707),
            .I(N__45696));
    Span4Mux_v I__11003 (
            .O(N__45704),
            .I(N__45691));
    LocalMux I__11002 (
            .O(N__45701),
            .I(N__45691));
    Span4Mux_h I__11001 (
            .O(N__45696),
            .I(N__45688));
    Span4Mux_h I__11000 (
            .O(N__45691),
            .I(N__45685));
    Odrv4 I__10999 (
            .O(N__45688),
            .I(\c0.data_out_5_3 ));
    Odrv4 I__10998 (
            .O(N__45685),
            .I(\c0.data_out_5_3 ));
    CascadeMux I__10997 (
            .O(N__45680),
            .I(\c0.n17635_cascade_ ));
    InMux I__10996 (
            .O(N__45677),
            .I(N__45674));
    LocalMux I__10995 (
            .O(N__45674),
            .I(N__45671));
    Span4Mux_s3_v I__10994 (
            .O(N__45671),
            .I(N__45668));
    Span4Mux_h I__10993 (
            .O(N__45668),
            .I(N__45665));
    Odrv4 I__10992 (
            .O(N__45665),
            .I(\c0.n17922 ));
    InMux I__10991 (
            .O(N__45662),
            .I(N__45659));
    LocalMux I__10990 (
            .O(N__45659),
            .I(N__45650));
    InMux I__10989 (
            .O(N__45658),
            .I(N__45647));
    InMux I__10988 (
            .O(N__45657),
            .I(N__45640));
    InMux I__10987 (
            .O(N__45656),
            .I(N__45640));
    InMux I__10986 (
            .O(N__45655),
            .I(N__45640));
    InMux I__10985 (
            .O(N__45654),
            .I(N__45635));
    InMux I__10984 (
            .O(N__45653),
            .I(N__45635));
    Span4Mux_h I__10983 (
            .O(N__45650),
            .I(N__45632));
    LocalMux I__10982 (
            .O(N__45647),
            .I(N__45629));
    LocalMux I__10981 (
            .O(N__45640),
            .I(N__45626));
    LocalMux I__10980 (
            .O(N__45635),
            .I(N__45622));
    Span4Mux_v I__10979 (
            .O(N__45632),
            .I(N__45619));
    Span4Mux_h I__10978 (
            .O(N__45629),
            .I(N__45614));
    Span4Mux_h I__10977 (
            .O(N__45626),
            .I(N__45614));
    InMux I__10976 (
            .O(N__45625),
            .I(N__45611));
    Span4Mux_h I__10975 (
            .O(N__45622),
            .I(N__45606));
    Span4Mux_v I__10974 (
            .O(N__45619),
            .I(N__45606));
    Odrv4 I__10973 (
            .O(N__45614),
            .I(\c0.data_out_7__7__N_519 ));
    LocalMux I__10972 (
            .O(N__45611),
            .I(\c0.data_out_7__7__N_519 ));
    Odrv4 I__10971 (
            .O(N__45606),
            .I(\c0.data_out_7__7__N_519 ));
    InMux I__10970 (
            .O(N__45599),
            .I(N__45591));
    InMux I__10969 (
            .O(N__45598),
            .I(N__45591));
    InMux I__10968 (
            .O(N__45597),
            .I(N__45587));
    InMux I__10967 (
            .O(N__45596),
            .I(N__45584));
    LocalMux I__10966 (
            .O(N__45591),
            .I(N__45581));
    InMux I__10965 (
            .O(N__45590),
            .I(N__45578));
    LocalMux I__10964 (
            .O(N__45587),
            .I(N__45575));
    LocalMux I__10963 (
            .O(N__45584),
            .I(N__45572));
    Span4Mux_v I__10962 (
            .O(N__45581),
            .I(N__45565));
    LocalMux I__10961 (
            .O(N__45578),
            .I(N__45565));
    Span4Mux_v I__10960 (
            .O(N__45575),
            .I(N__45565));
    Span4Mux_h I__10959 (
            .O(N__45572),
            .I(N__45562));
    Odrv4 I__10958 (
            .O(N__45565),
            .I(\c0.data_out_7_5 ));
    Odrv4 I__10957 (
            .O(N__45562),
            .I(\c0.data_out_7_5 ));
    InMux I__10956 (
            .O(N__45557),
            .I(N__45554));
    LocalMux I__10955 (
            .O(N__45554),
            .I(\c0.n17492 ));
    InMux I__10954 (
            .O(N__45551),
            .I(N__45548));
    LocalMux I__10953 (
            .O(N__45548),
            .I(\c0.n17635 ));
    CascadeMux I__10952 (
            .O(N__45545),
            .I(\c0.n17492_cascade_ ));
    InMux I__10951 (
            .O(N__45542),
            .I(N__45539));
    LocalMux I__10950 (
            .O(N__45539),
            .I(N__45536));
    Odrv4 I__10949 (
            .O(N__45536),
            .I(\c0.data_out_10_3 ));
    InMux I__10948 (
            .O(N__45533),
            .I(N__45530));
    LocalMux I__10947 (
            .O(N__45530),
            .I(\c0.n8_adj_2531 ));
    CascadeMux I__10946 (
            .O(N__45527),
            .I(\c0.n18069_cascade_ ));
    InMux I__10945 (
            .O(N__45524),
            .I(N__45521));
    LocalMux I__10944 (
            .O(N__45521),
            .I(N__45518));
    Span4Mux_h I__10943 (
            .O(N__45518),
            .I(N__45515));
    Odrv4 I__10942 (
            .O(N__45515),
            .I(\c0.n18070 ));
    InMux I__10941 (
            .O(N__45512),
            .I(N__45506));
    InMux I__10940 (
            .O(N__45511),
            .I(N__45506));
    LocalMux I__10939 (
            .O(N__45506),
            .I(N__45498));
    CascadeMux I__10938 (
            .O(N__45505),
            .I(N__45490));
    CascadeMux I__10937 (
            .O(N__45504),
            .I(N__45478));
    CascadeMux I__10936 (
            .O(N__45503),
            .I(N__45475));
    InMux I__10935 (
            .O(N__45502),
            .I(N__45469));
    InMux I__10934 (
            .O(N__45501),
            .I(N__45469));
    Span4Mux_v I__10933 (
            .O(N__45498),
            .I(N__45466));
    InMux I__10932 (
            .O(N__45497),
            .I(N__45461));
    InMux I__10931 (
            .O(N__45496),
            .I(N__45461));
    InMux I__10930 (
            .O(N__45495),
            .I(N__45457));
    CascadeMux I__10929 (
            .O(N__45494),
            .I(N__45448));
    InMux I__10928 (
            .O(N__45493),
            .I(N__45434));
    InMux I__10927 (
            .O(N__45490),
            .I(N__45434));
    InMux I__10926 (
            .O(N__45489),
            .I(N__45434));
    InMux I__10925 (
            .O(N__45488),
            .I(N__45434));
    InMux I__10924 (
            .O(N__45487),
            .I(N__45434));
    CascadeMux I__10923 (
            .O(N__45486),
            .I(N__45426));
    CascadeMux I__10922 (
            .O(N__45485),
            .I(N__45423));
    CascadeMux I__10921 (
            .O(N__45484),
            .I(N__45420));
    CascadeMux I__10920 (
            .O(N__45483),
            .I(N__45412));
    InMux I__10919 (
            .O(N__45482),
            .I(N__45406));
    InMux I__10918 (
            .O(N__45481),
            .I(N__45403));
    InMux I__10917 (
            .O(N__45478),
            .I(N__45396));
    InMux I__10916 (
            .O(N__45475),
            .I(N__45396));
    InMux I__10915 (
            .O(N__45474),
            .I(N__45396));
    LocalMux I__10914 (
            .O(N__45469),
            .I(N__45389));
    Span4Mux_h I__10913 (
            .O(N__45466),
            .I(N__45389));
    LocalMux I__10912 (
            .O(N__45461),
            .I(N__45389));
    InMux I__10911 (
            .O(N__45460),
            .I(N__45386));
    LocalMux I__10910 (
            .O(N__45457),
            .I(N__45382));
    InMux I__10909 (
            .O(N__45456),
            .I(N__45375));
    InMux I__10908 (
            .O(N__45455),
            .I(N__45375));
    InMux I__10907 (
            .O(N__45454),
            .I(N__45375));
    InMux I__10906 (
            .O(N__45453),
            .I(N__45360));
    InMux I__10905 (
            .O(N__45452),
            .I(N__45360));
    InMux I__10904 (
            .O(N__45451),
            .I(N__45360));
    InMux I__10903 (
            .O(N__45448),
            .I(N__45360));
    InMux I__10902 (
            .O(N__45447),
            .I(N__45360));
    InMux I__10901 (
            .O(N__45446),
            .I(N__45360));
    InMux I__10900 (
            .O(N__45445),
            .I(N__45360));
    LocalMux I__10899 (
            .O(N__45434),
            .I(N__45357));
    InMux I__10898 (
            .O(N__45433),
            .I(N__45354));
    InMux I__10897 (
            .O(N__45432),
            .I(N__45331));
    InMux I__10896 (
            .O(N__45431),
            .I(N__45331));
    InMux I__10895 (
            .O(N__45430),
            .I(N__45331));
    InMux I__10894 (
            .O(N__45429),
            .I(N__45331));
    InMux I__10893 (
            .O(N__45426),
            .I(N__45324));
    InMux I__10892 (
            .O(N__45423),
            .I(N__45324));
    InMux I__10891 (
            .O(N__45420),
            .I(N__45317));
    InMux I__10890 (
            .O(N__45419),
            .I(N__45317));
    InMux I__10889 (
            .O(N__45418),
            .I(N__45317));
    InMux I__10888 (
            .O(N__45417),
            .I(N__45302));
    InMux I__10887 (
            .O(N__45416),
            .I(N__45302));
    InMux I__10886 (
            .O(N__45415),
            .I(N__45302));
    InMux I__10885 (
            .O(N__45412),
            .I(N__45302));
    InMux I__10884 (
            .O(N__45411),
            .I(N__45302));
    InMux I__10883 (
            .O(N__45410),
            .I(N__45302));
    InMux I__10882 (
            .O(N__45409),
            .I(N__45302));
    LocalMux I__10881 (
            .O(N__45406),
            .I(N__45299));
    LocalMux I__10880 (
            .O(N__45403),
            .I(N__45296));
    LocalMux I__10879 (
            .O(N__45396),
            .I(N__45284));
    Span4Mux_h I__10878 (
            .O(N__45389),
            .I(N__45284));
    LocalMux I__10877 (
            .O(N__45386),
            .I(N__45284));
    InMux I__10876 (
            .O(N__45385),
            .I(N__45281));
    Span4Mux_v I__10875 (
            .O(N__45382),
            .I(N__45277));
    LocalMux I__10874 (
            .O(N__45375),
            .I(N__45270));
    LocalMux I__10873 (
            .O(N__45360),
            .I(N__45270));
    Span4Mux_v I__10872 (
            .O(N__45357),
            .I(N__45270));
    LocalMux I__10871 (
            .O(N__45354),
            .I(N__45267));
    InMux I__10870 (
            .O(N__45353),
            .I(N__45264));
    InMux I__10869 (
            .O(N__45352),
            .I(N__45255));
    InMux I__10868 (
            .O(N__45351),
            .I(N__45255));
    InMux I__10867 (
            .O(N__45350),
            .I(N__45255));
    InMux I__10866 (
            .O(N__45349),
            .I(N__45255));
    CascadeMux I__10865 (
            .O(N__45348),
            .I(N__45242));
    CascadeMux I__10864 (
            .O(N__45347),
            .I(N__45239));
    InMux I__10863 (
            .O(N__45346),
            .I(N__45235));
    CascadeMux I__10862 (
            .O(N__45345),
            .I(N__45228));
    InMux I__10861 (
            .O(N__45344),
            .I(N__45223));
    CascadeMux I__10860 (
            .O(N__45343),
            .I(N__45220));
    CascadeMux I__10859 (
            .O(N__45342),
            .I(N__45217));
    CascadeMux I__10858 (
            .O(N__45341),
            .I(N__45214));
    InMux I__10857 (
            .O(N__45340),
            .I(N__45193));
    LocalMux I__10856 (
            .O(N__45331),
            .I(N__45190));
    InMux I__10855 (
            .O(N__45330),
            .I(N__45185));
    InMux I__10854 (
            .O(N__45329),
            .I(N__45185));
    LocalMux I__10853 (
            .O(N__45324),
            .I(N__45178));
    LocalMux I__10852 (
            .O(N__45317),
            .I(N__45178));
    LocalMux I__10851 (
            .O(N__45302),
            .I(N__45178));
    Span4Mux_v I__10850 (
            .O(N__45299),
            .I(N__45173));
    Span4Mux_s2_h I__10849 (
            .O(N__45296),
            .I(N__45173));
    InMux I__10848 (
            .O(N__45295),
            .I(N__45168));
    InMux I__10847 (
            .O(N__45294),
            .I(N__45168));
    InMux I__10846 (
            .O(N__45293),
            .I(N__45165));
    InMux I__10845 (
            .O(N__45292),
            .I(N__45149));
    InMux I__10844 (
            .O(N__45291),
            .I(N__45146));
    Span4Mux_v I__10843 (
            .O(N__45284),
            .I(N__45143));
    LocalMux I__10842 (
            .O(N__45281),
            .I(N__45137));
    InMux I__10841 (
            .O(N__45280),
            .I(N__45134));
    Span4Mux_h I__10840 (
            .O(N__45277),
            .I(N__45123));
    Span4Mux_h I__10839 (
            .O(N__45270),
            .I(N__45123));
    Span4Mux_v I__10838 (
            .O(N__45267),
            .I(N__45123));
    LocalMux I__10837 (
            .O(N__45264),
            .I(N__45123));
    LocalMux I__10836 (
            .O(N__45255),
            .I(N__45123));
    InMux I__10835 (
            .O(N__45254),
            .I(N__45118));
    InMux I__10834 (
            .O(N__45253),
            .I(N__45118));
    CascadeMux I__10833 (
            .O(N__45252),
            .I(N__45107));
    InMux I__10832 (
            .O(N__45251),
            .I(N__45100));
    InMux I__10831 (
            .O(N__45250),
            .I(N__45100));
    InMux I__10830 (
            .O(N__45249),
            .I(N__45093));
    InMux I__10829 (
            .O(N__45248),
            .I(N__45093));
    InMux I__10828 (
            .O(N__45247),
            .I(N__45093));
    InMux I__10827 (
            .O(N__45246),
            .I(N__45088));
    InMux I__10826 (
            .O(N__45245),
            .I(N__45088));
    InMux I__10825 (
            .O(N__45242),
            .I(N__45081));
    InMux I__10824 (
            .O(N__45239),
            .I(N__45081));
    InMux I__10823 (
            .O(N__45238),
            .I(N__45081));
    LocalMux I__10822 (
            .O(N__45235),
            .I(N__45078));
    InMux I__10821 (
            .O(N__45234),
            .I(N__45072));
    InMux I__10820 (
            .O(N__45233),
            .I(N__45072));
    InMux I__10819 (
            .O(N__45232),
            .I(N__45069));
    InMux I__10818 (
            .O(N__45231),
            .I(N__45057));
    InMux I__10817 (
            .O(N__45228),
            .I(N__45057));
    InMux I__10816 (
            .O(N__45227),
            .I(N__45057));
    InMux I__10815 (
            .O(N__45226),
            .I(N__45057));
    LocalMux I__10814 (
            .O(N__45223),
            .I(N__45047));
    InMux I__10813 (
            .O(N__45220),
            .I(N__45032));
    InMux I__10812 (
            .O(N__45217),
            .I(N__45032));
    InMux I__10811 (
            .O(N__45214),
            .I(N__45032));
    InMux I__10810 (
            .O(N__45213),
            .I(N__45032));
    InMux I__10809 (
            .O(N__45212),
            .I(N__45032));
    InMux I__10808 (
            .O(N__45211),
            .I(N__45032));
    InMux I__10807 (
            .O(N__45210),
            .I(N__45032));
    InMux I__10806 (
            .O(N__45209),
            .I(N__45029));
    InMux I__10805 (
            .O(N__45208),
            .I(N__45020));
    InMux I__10804 (
            .O(N__45207),
            .I(N__45020));
    InMux I__10803 (
            .O(N__45206),
            .I(N__45020));
    InMux I__10802 (
            .O(N__45205),
            .I(N__45020));
    InMux I__10801 (
            .O(N__45204),
            .I(N__45017));
    InMux I__10800 (
            .O(N__45203),
            .I(N__45014));
    InMux I__10799 (
            .O(N__45202),
            .I(N__45007));
    InMux I__10798 (
            .O(N__45201),
            .I(N__45007));
    InMux I__10797 (
            .O(N__45200),
            .I(N__45007));
    InMux I__10796 (
            .O(N__45199),
            .I(N__45000));
    InMux I__10795 (
            .O(N__45198),
            .I(N__45000));
    InMux I__10794 (
            .O(N__45197),
            .I(N__45000));
    InMux I__10793 (
            .O(N__45196),
            .I(N__44997));
    LocalMux I__10792 (
            .O(N__45193),
            .I(N__44984));
    Span4Mux_v I__10791 (
            .O(N__45190),
            .I(N__44984));
    LocalMux I__10790 (
            .O(N__45185),
            .I(N__44984));
    Span4Mux_v I__10789 (
            .O(N__45178),
            .I(N__44984));
    Span4Mux_h I__10788 (
            .O(N__45173),
            .I(N__44984));
    LocalMux I__10787 (
            .O(N__45168),
            .I(N__44984));
    LocalMux I__10786 (
            .O(N__45165),
            .I(N__44981));
    InMux I__10785 (
            .O(N__45164),
            .I(N__44978));
    InMux I__10784 (
            .O(N__45163),
            .I(N__44969));
    InMux I__10783 (
            .O(N__45162),
            .I(N__44969));
    InMux I__10782 (
            .O(N__45161),
            .I(N__44969));
    InMux I__10781 (
            .O(N__45160),
            .I(N__44969));
    InMux I__10780 (
            .O(N__45159),
            .I(N__44963));
    InMux I__10779 (
            .O(N__45158),
            .I(N__44963));
    InMux I__10778 (
            .O(N__45157),
            .I(N__44960));
    InMux I__10777 (
            .O(N__45156),
            .I(N__44953));
    InMux I__10776 (
            .O(N__45155),
            .I(N__44953));
    InMux I__10775 (
            .O(N__45154),
            .I(N__44953));
    CascadeMux I__10774 (
            .O(N__45153),
            .I(N__44941));
    CascadeMux I__10773 (
            .O(N__45152),
            .I(N__44938));
    LocalMux I__10772 (
            .O(N__45149),
            .I(N__44929));
    LocalMux I__10771 (
            .O(N__45146),
            .I(N__44929));
    Span4Mux_v I__10770 (
            .O(N__45143),
            .I(N__44926));
    InMux I__10769 (
            .O(N__45142),
            .I(N__44923));
    InMux I__10768 (
            .O(N__45141),
            .I(N__44918));
    InMux I__10767 (
            .O(N__45140),
            .I(N__44918));
    Span4Mux_h I__10766 (
            .O(N__45137),
            .I(N__44913));
    LocalMux I__10765 (
            .O(N__45134),
            .I(N__44913));
    Span4Mux_h I__10764 (
            .O(N__45123),
            .I(N__44908));
    LocalMux I__10763 (
            .O(N__45118),
            .I(N__44908));
    InMux I__10762 (
            .O(N__45117),
            .I(N__44903));
    InMux I__10761 (
            .O(N__45116),
            .I(N__44903));
    InMux I__10760 (
            .O(N__45115),
            .I(N__44899));
    InMux I__10759 (
            .O(N__45114),
            .I(N__44894));
    InMux I__10758 (
            .O(N__45113),
            .I(N__44894));
    CascadeMux I__10757 (
            .O(N__45112),
            .I(N__44891));
    InMux I__10756 (
            .O(N__45111),
            .I(N__44885));
    InMux I__10755 (
            .O(N__45110),
            .I(N__44876));
    InMux I__10754 (
            .O(N__45107),
            .I(N__44876));
    InMux I__10753 (
            .O(N__45106),
            .I(N__44876));
    InMux I__10752 (
            .O(N__45105),
            .I(N__44876));
    LocalMux I__10751 (
            .O(N__45100),
            .I(N__44867));
    LocalMux I__10750 (
            .O(N__45093),
            .I(N__44867));
    LocalMux I__10749 (
            .O(N__45088),
            .I(N__44867));
    LocalMux I__10748 (
            .O(N__45081),
            .I(N__44867));
    Span4Mux_v I__10747 (
            .O(N__45078),
            .I(N__44862));
    InMux I__10746 (
            .O(N__45077),
            .I(N__44859));
    LocalMux I__10745 (
            .O(N__45072),
            .I(N__44854));
    LocalMux I__10744 (
            .O(N__45069),
            .I(N__44854));
    InMux I__10743 (
            .O(N__45068),
            .I(N__44847));
    InMux I__10742 (
            .O(N__45067),
            .I(N__44847));
    InMux I__10741 (
            .O(N__45066),
            .I(N__44847));
    LocalMux I__10740 (
            .O(N__45057),
            .I(N__44844));
    InMux I__10739 (
            .O(N__45056),
            .I(N__44839));
    InMux I__10738 (
            .O(N__45055),
            .I(N__44839));
    InMux I__10737 (
            .O(N__45054),
            .I(N__44836));
    InMux I__10736 (
            .O(N__45053),
            .I(N__44827));
    InMux I__10735 (
            .O(N__45052),
            .I(N__44827));
    InMux I__10734 (
            .O(N__45051),
            .I(N__44827));
    InMux I__10733 (
            .O(N__45050),
            .I(N__44827));
    Span4Mux_h I__10732 (
            .O(N__45047),
            .I(N__44824));
    LocalMux I__10731 (
            .O(N__45032),
            .I(N__44817));
    LocalMux I__10730 (
            .O(N__45029),
            .I(N__44817));
    LocalMux I__10729 (
            .O(N__45020),
            .I(N__44817));
    LocalMux I__10728 (
            .O(N__45017),
            .I(N__44812));
    LocalMux I__10727 (
            .O(N__45014),
            .I(N__44812));
    LocalMux I__10726 (
            .O(N__45007),
            .I(N__44801));
    LocalMux I__10725 (
            .O(N__45000),
            .I(N__44801));
    LocalMux I__10724 (
            .O(N__44997),
            .I(N__44801));
    Span4Mux_h I__10723 (
            .O(N__44984),
            .I(N__44801));
    Span4Mux_h I__10722 (
            .O(N__44981),
            .I(N__44801));
    LocalMux I__10721 (
            .O(N__44978),
            .I(N__44796));
    LocalMux I__10720 (
            .O(N__44969),
            .I(N__44796));
    CascadeMux I__10719 (
            .O(N__44968),
            .I(N__44793));
    LocalMux I__10718 (
            .O(N__44963),
            .I(N__44786));
    LocalMux I__10717 (
            .O(N__44960),
            .I(N__44786));
    LocalMux I__10716 (
            .O(N__44953),
            .I(N__44783));
    InMux I__10715 (
            .O(N__44952),
            .I(N__44776));
    InMux I__10714 (
            .O(N__44951),
            .I(N__44776));
    InMux I__10713 (
            .O(N__44950),
            .I(N__44776));
    InMux I__10712 (
            .O(N__44949),
            .I(N__44769));
    InMux I__10711 (
            .O(N__44948),
            .I(N__44769));
    InMux I__10710 (
            .O(N__44947),
            .I(N__44769));
    InMux I__10709 (
            .O(N__44946),
            .I(N__44762));
    InMux I__10708 (
            .O(N__44945),
            .I(N__44762));
    InMux I__10707 (
            .O(N__44944),
            .I(N__44759));
    InMux I__10706 (
            .O(N__44941),
            .I(N__44746));
    InMux I__10705 (
            .O(N__44938),
            .I(N__44746));
    InMux I__10704 (
            .O(N__44937),
            .I(N__44746));
    InMux I__10703 (
            .O(N__44936),
            .I(N__44746));
    InMux I__10702 (
            .O(N__44935),
            .I(N__44746));
    InMux I__10701 (
            .O(N__44934),
            .I(N__44746));
    Span4Mux_h I__10700 (
            .O(N__44929),
            .I(N__44741));
    Span4Mux_v I__10699 (
            .O(N__44926),
            .I(N__44741));
    LocalMux I__10698 (
            .O(N__44923),
            .I(N__44730));
    LocalMux I__10697 (
            .O(N__44918),
            .I(N__44730));
    Span4Mux_h I__10696 (
            .O(N__44913),
            .I(N__44730));
    Span4Mux_v I__10695 (
            .O(N__44908),
            .I(N__44730));
    LocalMux I__10694 (
            .O(N__44903),
            .I(N__44730));
    InMux I__10693 (
            .O(N__44902),
            .I(N__44727));
    LocalMux I__10692 (
            .O(N__44899),
            .I(N__44722));
    LocalMux I__10691 (
            .O(N__44894),
            .I(N__44722));
    InMux I__10690 (
            .O(N__44891),
            .I(N__44713));
    InMux I__10689 (
            .O(N__44890),
            .I(N__44713));
    InMux I__10688 (
            .O(N__44889),
            .I(N__44713));
    InMux I__10687 (
            .O(N__44888),
            .I(N__44713));
    LocalMux I__10686 (
            .O(N__44885),
            .I(N__44710));
    LocalMux I__10685 (
            .O(N__44876),
            .I(N__44705));
    Span4Mux_v I__10684 (
            .O(N__44867),
            .I(N__44705));
    InMux I__10683 (
            .O(N__44866),
            .I(N__44700));
    InMux I__10682 (
            .O(N__44865),
            .I(N__44700));
    Span4Mux_v I__10681 (
            .O(N__44862),
            .I(N__44689));
    LocalMux I__10680 (
            .O(N__44859),
            .I(N__44689));
    Span4Mux_v I__10679 (
            .O(N__44854),
            .I(N__44689));
    LocalMux I__10678 (
            .O(N__44847),
            .I(N__44689));
    Span4Mux_h I__10677 (
            .O(N__44844),
            .I(N__44689));
    LocalMux I__10676 (
            .O(N__44839),
            .I(N__44672));
    LocalMux I__10675 (
            .O(N__44836),
            .I(N__44672));
    LocalMux I__10674 (
            .O(N__44827),
            .I(N__44672));
    Span4Mux_h I__10673 (
            .O(N__44824),
            .I(N__44672));
    Span4Mux_v I__10672 (
            .O(N__44817),
            .I(N__44672));
    Span4Mux_h I__10671 (
            .O(N__44812),
            .I(N__44672));
    Span4Mux_v I__10670 (
            .O(N__44801),
            .I(N__44672));
    Span4Mux_h I__10669 (
            .O(N__44796),
            .I(N__44672));
    InMux I__10668 (
            .O(N__44793),
            .I(N__44665));
    InMux I__10667 (
            .O(N__44792),
            .I(N__44665));
    InMux I__10666 (
            .O(N__44791),
            .I(N__44665));
    Span4Mux_h I__10665 (
            .O(N__44786),
            .I(N__44656));
    Span4Mux_h I__10664 (
            .O(N__44783),
            .I(N__44656));
    LocalMux I__10663 (
            .O(N__44776),
            .I(N__44656));
    LocalMux I__10662 (
            .O(N__44769),
            .I(N__44656));
    CascadeMux I__10661 (
            .O(N__44768),
            .I(N__44653));
    InMux I__10660 (
            .O(N__44767),
            .I(N__44645));
    LocalMux I__10659 (
            .O(N__44762),
            .I(N__44640));
    LocalMux I__10658 (
            .O(N__44759),
            .I(N__44640));
    LocalMux I__10657 (
            .O(N__44746),
            .I(N__44637));
    Span4Mux_h I__10656 (
            .O(N__44741),
            .I(N__44632));
    Span4Mux_v I__10655 (
            .O(N__44730),
            .I(N__44632));
    LocalMux I__10654 (
            .O(N__44727),
            .I(N__44625));
    Span4Mux_v I__10653 (
            .O(N__44722),
            .I(N__44625));
    LocalMux I__10652 (
            .O(N__44713),
            .I(N__44625));
    Span4Mux_v I__10651 (
            .O(N__44710),
            .I(N__44614));
    Span4Mux_h I__10650 (
            .O(N__44705),
            .I(N__44614));
    LocalMux I__10649 (
            .O(N__44700),
            .I(N__44614));
    Span4Mux_h I__10648 (
            .O(N__44689),
            .I(N__44614));
    Span4Mux_v I__10647 (
            .O(N__44672),
            .I(N__44614));
    LocalMux I__10646 (
            .O(N__44665),
            .I(N__44609));
    Span4Mux_v I__10645 (
            .O(N__44656),
            .I(N__44609));
    InMux I__10644 (
            .O(N__44653),
            .I(N__44606));
    InMux I__10643 (
            .O(N__44652),
            .I(N__44601));
    InMux I__10642 (
            .O(N__44651),
            .I(N__44601));
    InMux I__10641 (
            .O(N__44650),
            .I(N__44594));
    InMux I__10640 (
            .O(N__44649),
            .I(N__44594));
    InMux I__10639 (
            .O(N__44648),
            .I(N__44594));
    LocalMux I__10638 (
            .O(N__44645),
            .I(N__44589));
    Span12Mux_h I__10637 (
            .O(N__44640),
            .I(N__44589));
    Span4Mux_h I__10636 (
            .O(N__44637),
            .I(N__44584));
    Span4Mux_v I__10635 (
            .O(N__44632),
            .I(N__44584));
    Span4Mux_v I__10634 (
            .O(N__44625),
            .I(N__44579));
    Span4Mux_v I__10633 (
            .O(N__44614),
            .I(N__44579));
    Span4Mux_v I__10632 (
            .O(N__44609),
            .I(N__44576));
    LocalMux I__10631 (
            .O(N__44606),
            .I(rx_data_ready));
    LocalMux I__10630 (
            .O(N__44601),
            .I(rx_data_ready));
    LocalMux I__10629 (
            .O(N__44594),
            .I(rx_data_ready));
    Odrv12 I__10628 (
            .O(N__44589),
            .I(rx_data_ready));
    Odrv4 I__10627 (
            .O(N__44584),
            .I(rx_data_ready));
    Odrv4 I__10626 (
            .O(N__44579),
            .I(rx_data_ready));
    Odrv4 I__10625 (
            .O(N__44576),
            .I(rx_data_ready));
    InMux I__10624 (
            .O(N__44561),
            .I(N__44558));
    LocalMux I__10623 (
            .O(N__44558),
            .I(N__44555));
    Span4Mux_h I__10622 (
            .O(N__44555),
            .I(N__44552));
    Span4Mux_h I__10621 (
            .O(N__44552),
            .I(N__44548));
    InMux I__10620 (
            .O(N__44551),
            .I(N__44545));
    Odrv4 I__10619 (
            .O(N__44548),
            .I(data_in_14_6));
    LocalMux I__10618 (
            .O(N__44545),
            .I(data_in_14_6));
    InMux I__10617 (
            .O(N__44540),
            .I(N__44537));
    LocalMux I__10616 (
            .O(N__44537),
            .I(N__44534));
    Span4Mux_h I__10615 (
            .O(N__44534),
            .I(N__44530));
    InMux I__10614 (
            .O(N__44533),
            .I(N__44527));
    Odrv4 I__10613 (
            .O(N__44530),
            .I(data_in_13_6));
    LocalMux I__10612 (
            .O(N__44527),
            .I(data_in_13_6));
    InMux I__10611 (
            .O(N__44522),
            .I(N__44519));
    LocalMux I__10610 (
            .O(N__44519),
            .I(N__44516));
    Odrv12 I__10609 (
            .O(N__44516),
            .I(\c0.n17445 ));
    InMux I__10608 (
            .O(N__44513),
            .I(N__44509));
    InMux I__10607 (
            .O(N__44512),
            .I(N__44506));
    LocalMux I__10606 (
            .O(N__44509),
            .I(N__44503));
    LocalMux I__10605 (
            .O(N__44506),
            .I(N__44500));
    Odrv4 I__10604 (
            .O(N__44503),
            .I(\c0.n17510 ));
    Odrv4 I__10603 (
            .O(N__44500),
            .I(\c0.n17510 ));
    InMux I__10602 (
            .O(N__44495),
            .I(N__44492));
    LocalMux I__10601 (
            .O(N__44492),
            .I(\c0.data_out_9_1 ));
    InMux I__10600 (
            .O(N__44489),
            .I(N__44485));
    InMux I__10599 (
            .O(N__44488),
            .I(N__44482));
    LocalMux I__10598 (
            .O(N__44485),
            .I(N__44478));
    LocalMux I__10597 (
            .O(N__44482),
            .I(N__44475));
    InMux I__10596 (
            .O(N__44481),
            .I(N__44471));
    Span4Mux_h I__10595 (
            .O(N__44478),
            .I(N__44468));
    Span4Mux_v I__10594 (
            .O(N__44475),
            .I(N__44465));
    InMux I__10593 (
            .O(N__44474),
            .I(N__44462));
    LocalMux I__10592 (
            .O(N__44471),
            .I(data_out_8_1));
    Odrv4 I__10591 (
            .O(N__44468),
            .I(data_out_8_1));
    Odrv4 I__10590 (
            .O(N__44465),
            .I(data_out_8_1));
    LocalMux I__10589 (
            .O(N__44462),
            .I(data_out_8_1));
    InMux I__10588 (
            .O(N__44453),
            .I(N__44450));
    LocalMux I__10587 (
            .O(N__44450),
            .I(\c0.n8_adj_2519 ));
    InMux I__10586 (
            .O(N__44447),
            .I(N__44444));
    LocalMux I__10585 (
            .O(N__44444),
            .I(N__44441));
    Span4Mux_h I__10584 (
            .O(N__44441),
            .I(N__44438));
    Odrv4 I__10583 (
            .O(N__44438),
            .I(\c0.n8_adj_2535 ));
    InMux I__10582 (
            .O(N__44435),
            .I(N__44432));
    LocalMux I__10581 (
            .O(N__44432),
            .I(N__44429));
    Span4Mux_h I__10580 (
            .O(N__44429),
            .I(N__44426));
    Odrv4 I__10579 (
            .O(N__44426),
            .I(\c0.n17398 ));
    CascadeMux I__10578 (
            .O(N__44423),
            .I(N__44420));
    InMux I__10577 (
            .O(N__44420),
            .I(N__44416));
    InMux I__10576 (
            .O(N__44419),
            .I(N__44413));
    LocalMux I__10575 (
            .O(N__44416),
            .I(N__44410));
    LocalMux I__10574 (
            .O(N__44413),
            .I(N__44407));
    Odrv4 I__10573 (
            .O(N__44410),
            .I(\c0.n9091 ));
    Odrv12 I__10572 (
            .O(N__44407),
            .I(\c0.n9091 ));
    InMux I__10571 (
            .O(N__44402),
            .I(N__44399));
    LocalMux I__10570 (
            .O(N__44399),
            .I(\c0.data_out_9_4 ));
    InMux I__10569 (
            .O(N__44396),
            .I(N__44392));
    InMux I__10568 (
            .O(N__44395),
            .I(N__44389));
    LocalMux I__10567 (
            .O(N__44392),
            .I(N__44383));
    LocalMux I__10566 (
            .O(N__44389),
            .I(N__44383));
    InMux I__10565 (
            .O(N__44388),
            .I(N__44380));
    Odrv4 I__10564 (
            .O(N__44383),
            .I(\c0.data_out_6_1 ));
    LocalMux I__10563 (
            .O(N__44380),
            .I(\c0.data_out_6_1 ));
    CascadeMux I__10562 (
            .O(N__44375),
            .I(N__44372));
    InMux I__10561 (
            .O(N__44372),
            .I(N__44369));
    LocalMux I__10560 (
            .O(N__44369),
            .I(N__44365));
    InMux I__10559 (
            .O(N__44368),
            .I(N__44362));
    Span4Mux_h I__10558 (
            .O(N__44365),
            .I(N__44359));
    LocalMux I__10557 (
            .O(N__44362),
            .I(\c0.n17499 ));
    Odrv4 I__10556 (
            .O(N__44359),
            .I(\c0.n17499 ));
    InMux I__10555 (
            .O(N__44354),
            .I(N__44351));
    LocalMux I__10554 (
            .O(N__44351),
            .I(N__44348));
    Span4Mux_h I__10553 (
            .O(N__44348),
            .I(N__44345));
    Odrv4 I__10552 (
            .O(N__44345),
            .I(\c0.n6_adj_2451 ));
    CascadeMux I__10551 (
            .O(N__44342),
            .I(\c0.n18065_cascade_ ));
    InMux I__10550 (
            .O(N__44339),
            .I(N__44336));
    LocalMux I__10549 (
            .O(N__44336),
            .I(N__44333));
    Odrv4 I__10548 (
            .O(N__44333),
            .I(tx_data_5_N_keep));
    CascadeMux I__10547 (
            .O(N__44330),
            .I(N__44327));
    InMux I__10546 (
            .O(N__44327),
            .I(N__44324));
    LocalMux I__10545 (
            .O(N__44324),
            .I(N__44321));
    Odrv4 I__10544 (
            .O(N__44321),
            .I(\c0.n18014 ));
    InMux I__10543 (
            .O(N__44318),
            .I(N__44315));
    LocalMux I__10542 (
            .O(N__44315),
            .I(tx_data_1_N_keep));
    InMux I__10541 (
            .O(N__44312),
            .I(N__44309));
    LocalMux I__10540 (
            .O(N__44309),
            .I(N__44306));
    Odrv4 I__10539 (
            .O(N__44306),
            .I(\c0.n17943 ));
    CascadeMux I__10538 (
            .O(N__44303),
            .I(\c0.n5_adj_2481_cascade_ ));
    InMux I__10537 (
            .O(N__44300),
            .I(N__44297));
    LocalMux I__10536 (
            .O(N__44297),
            .I(\c0.n18091 ));
    CascadeMux I__10535 (
            .O(N__44294),
            .I(\c0.n18402_cascade_ ));
    InMux I__10534 (
            .O(N__44291),
            .I(N__44288));
    LocalMux I__10533 (
            .O(N__44288),
            .I(N__44285));
    Span4Mux_h I__10532 (
            .O(N__44285),
            .I(N__44282));
    Odrv4 I__10531 (
            .O(N__44282),
            .I(\c0.n2_adj_2476 ));
    InMux I__10530 (
            .O(N__44279),
            .I(N__44276));
    LocalMux I__10529 (
            .O(N__44276),
            .I(\c0.n18405 ));
    InMux I__10528 (
            .O(N__44273),
            .I(N__44269));
    CascadeMux I__10527 (
            .O(N__44272),
            .I(N__44265));
    LocalMux I__10526 (
            .O(N__44269),
            .I(N__44261));
    InMux I__10525 (
            .O(N__44268),
            .I(N__44258));
    InMux I__10524 (
            .O(N__44265),
            .I(N__44255));
    InMux I__10523 (
            .O(N__44264),
            .I(N__44252));
    Span4Mux_v I__10522 (
            .O(N__44261),
            .I(N__44247));
    LocalMux I__10521 (
            .O(N__44258),
            .I(N__44247));
    LocalMux I__10520 (
            .O(N__44255),
            .I(\c0.data_out_5_1 ));
    LocalMux I__10519 (
            .O(N__44252),
            .I(\c0.data_out_5_1 ));
    Odrv4 I__10518 (
            .O(N__44247),
            .I(\c0.data_out_5_1 ));
    CascadeMux I__10517 (
            .O(N__44240),
            .I(\c0.n45_adj_2518_cascade_ ));
    InMux I__10516 (
            .O(N__44237),
            .I(N__44234));
    LocalMux I__10515 (
            .O(N__44234),
            .I(N__44231));
    Odrv4 I__10514 (
            .O(N__44231),
            .I(\c0.n1_adj_2522 ));
    CascadeMux I__10513 (
            .O(N__44228),
            .I(\c0.n46_cascade_ ));
    InMux I__10512 (
            .O(N__44225),
            .I(N__44222));
    LocalMux I__10511 (
            .O(N__44222),
            .I(\c0.n44_adj_2524 ));
    CascadeMux I__10510 (
            .O(N__44219),
            .I(N__44216));
    InMux I__10509 (
            .O(N__44216),
            .I(N__44213));
    LocalMux I__10508 (
            .O(N__44213),
            .I(N__44210));
    Span4Mux_v I__10507 (
            .O(N__44210),
            .I(N__44206));
    CascadeMux I__10506 (
            .O(N__44209),
            .I(N__44203));
    Span4Mux_h I__10505 (
            .O(N__44206),
            .I(N__44200));
    InMux I__10504 (
            .O(N__44203),
            .I(N__44197));
    Odrv4 I__10503 (
            .O(N__44200),
            .I(rand_setpoint_9));
    LocalMux I__10502 (
            .O(N__44197),
            .I(rand_setpoint_9));
    CEMux I__10501 (
            .O(N__44192),
            .I(N__44189));
    LocalMux I__10500 (
            .O(N__44189),
            .I(N__44183));
    CEMux I__10499 (
            .O(N__44188),
            .I(N__44180));
    CEMux I__10498 (
            .O(N__44187),
            .I(N__44177));
    CEMux I__10497 (
            .O(N__44186),
            .I(N__44174));
    Span4Mux_h I__10496 (
            .O(N__44183),
            .I(N__44168));
    LocalMux I__10495 (
            .O(N__44180),
            .I(N__44168));
    LocalMux I__10494 (
            .O(N__44177),
            .I(N__44165));
    LocalMux I__10493 (
            .O(N__44174),
            .I(N__44162));
    CEMux I__10492 (
            .O(N__44173),
            .I(N__44159));
    Span4Mux_h I__10491 (
            .O(N__44168),
            .I(N__44156));
    Sp12to4 I__10490 (
            .O(N__44165),
            .I(N__44153));
    Span4Mux_h I__10489 (
            .O(N__44162),
            .I(N__44148));
    LocalMux I__10488 (
            .O(N__44159),
            .I(N__44148));
    Odrv4 I__10487 (
            .O(N__44156),
            .I(\c0.n9518 ));
    Odrv12 I__10486 (
            .O(N__44153),
            .I(\c0.n9518 ));
    Odrv4 I__10485 (
            .O(N__44148),
            .I(\c0.n9518 ));
    InMux I__10484 (
            .O(N__44141),
            .I(N__44135));
    InMux I__10483 (
            .O(N__44140),
            .I(N__44132));
    InMux I__10482 (
            .O(N__44139),
            .I(N__44129));
    InMux I__10481 (
            .O(N__44138),
            .I(N__44125));
    LocalMux I__10480 (
            .O(N__44135),
            .I(N__44120));
    LocalMux I__10479 (
            .O(N__44132),
            .I(N__44115));
    LocalMux I__10478 (
            .O(N__44129),
            .I(N__44115));
    InMux I__10477 (
            .O(N__44128),
            .I(N__44112));
    LocalMux I__10476 (
            .O(N__44125),
            .I(N__44109));
    InMux I__10475 (
            .O(N__44124),
            .I(N__44106));
    InMux I__10474 (
            .O(N__44123),
            .I(N__44103));
    Span4Mux_h I__10473 (
            .O(N__44120),
            .I(N__44100));
    Span4Mux_v I__10472 (
            .O(N__44115),
            .I(N__44095));
    LocalMux I__10471 (
            .O(N__44112),
            .I(N__44095));
    Odrv12 I__10470 (
            .O(N__44109),
            .I(data_out_6__2__N_804));
    LocalMux I__10469 (
            .O(N__44106),
            .I(data_out_6__2__N_804));
    LocalMux I__10468 (
            .O(N__44103),
            .I(data_out_6__2__N_804));
    Odrv4 I__10467 (
            .O(N__44100),
            .I(data_out_6__2__N_804));
    Odrv4 I__10466 (
            .O(N__44095),
            .I(data_out_6__2__N_804));
    InMux I__10465 (
            .O(N__44084),
            .I(N__44081));
    LocalMux I__10464 (
            .O(N__44081),
            .I(N__44077));
    InMux I__10463 (
            .O(N__44080),
            .I(N__44074));
    Odrv4 I__10462 (
            .O(N__44077),
            .I(\c0.n17457 ));
    LocalMux I__10461 (
            .O(N__44074),
            .I(\c0.n17457 ));
    InMux I__10460 (
            .O(N__44069),
            .I(N__44066));
    LocalMux I__10459 (
            .O(N__44066),
            .I(\c0.n17654 ));
    InMux I__10458 (
            .O(N__44063),
            .I(N__44060));
    LocalMux I__10457 (
            .O(N__44060),
            .I(N__44057));
    Span4Mux_h I__10456 (
            .O(N__44057),
            .I(N__44054));
    Odrv4 I__10455 (
            .O(N__44054),
            .I(\c0.n18061 ));
    InMux I__10454 (
            .O(N__44051),
            .I(N__44047));
    InMux I__10453 (
            .O(N__44050),
            .I(N__44043));
    LocalMux I__10452 (
            .O(N__44047),
            .I(N__44040));
    InMux I__10451 (
            .O(N__44046),
            .I(N__44037));
    LocalMux I__10450 (
            .O(N__44043),
            .I(N__44034));
    Span4Mux_s3_v I__10449 (
            .O(N__44040),
            .I(N__44029));
    LocalMux I__10448 (
            .O(N__44037),
            .I(N__44029));
    Span4Mux_v I__10447 (
            .O(N__44034),
            .I(N__44026));
    Span4Mux_h I__10446 (
            .O(N__44029),
            .I(N__44023));
    Span4Mux_h I__10445 (
            .O(N__44026),
            .I(N__44020));
    Odrv4 I__10444 (
            .O(N__44023),
            .I(\c0.data_out_7__5__N_543 ));
    Odrv4 I__10443 (
            .O(N__44020),
            .I(\c0.data_out_7__5__N_543 ));
    InMux I__10442 (
            .O(N__44015),
            .I(N__44010));
    InMux I__10441 (
            .O(N__44014),
            .I(N__44005));
    InMux I__10440 (
            .O(N__44013),
            .I(N__44005));
    LocalMux I__10439 (
            .O(N__44010),
            .I(N__44002));
    LocalMux I__10438 (
            .O(N__44005),
            .I(N__43995));
    Span4Mux_v I__10437 (
            .O(N__44002),
            .I(N__43995));
    CascadeMux I__10436 (
            .O(N__44001),
            .I(N__43991));
    InMux I__10435 (
            .O(N__44000),
            .I(N__43988));
    Span4Mux_h I__10434 (
            .O(N__43995),
            .I(N__43985));
    InMux I__10433 (
            .O(N__43994),
            .I(N__43980));
    InMux I__10432 (
            .O(N__43991),
            .I(N__43980));
    LocalMux I__10431 (
            .O(N__43988),
            .I(data_out_6__1__N_850));
    Odrv4 I__10430 (
            .O(N__43985),
            .I(data_out_6__1__N_850));
    LocalMux I__10429 (
            .O(N__43980),
            .I(data_out_6__1__N_850));
    InMux I__10428 (
            .O(N__43973),
            .I(N__43970));
    LocalMux I__10427 (
            .O(N__43970),
            .I(N__43967));
    Span4Mux_v I__10426 (
            .O(N__43967),
            .I(N__43964));
    Odrv4 I__10425 (
            .O(N__43964),
            .I(\c0.n2 ));
    CascadeMux I__10424 (
            .O(N__43961),
            .I(N__43958));
    InMux I__10423 (
            .O(N__43958),
            .I(N__43955));
    LocalMux I__10422 (
            .O(N__43955),
            .I(N__43952));
    Odrv12 I__10421 (
            .O(N__43952),
            .I(\c0.n18060 ));
    InMux I__10420 (
            .O(N__43949),
            .I(N__43941));
    InMux I__10419 (
            .O(N__43948),
            .I(N__43937));
    InMux I__10418 (
            .O(N__43947),
            .I(N__43934));
    CascadeMux I__10417 (
            .O(N__43946),
            .I(N__43931));
    InMux I__10416 (
            .O(N__43945),
            .I(N__43926));
    InMux I__10415 (
            .O(N__43944),
            .I(N__43926));
    LocalMux I__10414 (
            .O(N__43941),
            .I(N__43923));
    InMux I__10413 (
            .O(N__43940),
            .I(N__43920));
    LocalMux I__10412 (
            .O(N__43937),
            .I(N__43917));
    LocalMux I__10411 (
            .O(N__43934),
            .I(N__43914));
    InMux I__10410 (
            .O(N__43931),
            .I(N__43911));
    LocalMux I__10409 (
            .O(N__43926),
            .I(N__43906));
    Span4Mux_h I__10408 (
            .O(N__43923),
            .I(N__43906));
    LocalMux I__10407 (
            .O(N__43920),
            .I(N__43901));
    Span12Mux_h I__10406 (
            .O(N__43917),
            .I(N__43901));
    Span4Mux_h I__10405 (
            .O(N__43914),
            .I(N__43898));
    LocalMux I__10404 (
            .O(N__43911),
            .I(data_out_0_5));
    Odrv4 I__10403 (
            .O(N__43906),
            .I(data_out_0_5));
    Odrv12 I__10402 (
            .O(N__43901),
            .I(data_out_0_5));
    Odrv4 I__10401 (
            .O(N__43898),
            .I(data_out_0_5));
    InMux I__10400 (
            .O(N__43889),
            .I(N__43886));
    LocalMux I__10399 (
            .O(N__43886),
            .I(N__43883));
    Span4Mux_h I__10398 (
            .O(N__43883),
            .I(N__43880));
    Span4Mux_h I__10397 (
            .O(N__43880),
            .I(N__43876));
    InMux I__10396 (
            .O(N__43879),
            .I(N__43873));
    Odrv4 I__10395 (
            .O(N__43876),
            .I(rand_setpoint_21));
    LocalMux I__10394 (
            .O(N__43873),
            .I(rand_setpoint_21));
    CascadeMux I__10393 (
            .O(N__43868),
            .I(\c0.n9656_cascade_ ));
    InMux I__10392 (
            .O(N__43865),
            .I(N__43862));
    LocalMux I__10391 (
            .O(N__43862),
            .I(N__43859));
    Span4Mux_s3_v I__10390 (
            .O(N__43859),
            .I(N__43855));
    CascadeMux I__10389 (
            .O(N__43858),
            .I(N__43852));
    Span4Mux_h I__10388 (
            .O(N__43855),
            .I(N__43849));
    InMux I__10387 (
            .O(N__43852),
            .I(N__43846));
    Odrv4 I__10386 (
            .O(N__43849),
            .I(rand_setpoint_17));
    LocalMux I__10385 (
            .O(N__43846),
            .I(rand_setpoint_17));
    CascadeMux I__10384 (
            .O(N__43841),
            .I(\c0.n2251_cascade_ ));
    InMux I__10383 (
            .O(N__43838),
            .I(N__43835));
    LocalMux I__10382 (
            .O(N__43835),
            .I(N__43832));
    Odrv12 I__10381 (
            .O(N__43832),
            .I(\c0.n17962 ));
    CascadeMux I__10380 (
            .O(N__43829),
            .I(N__43826));
    InMux I__10379 (
            .O(N__43826),
            .I(N__43820));
    InMux I__10378 (
            .O(N__43825),
            .I(N__43820));
    LocalMux I__10377 (
            .O(N__43820),
            .I(N__43817));
    Span4Mux_h I__10376 (
            .O(N__43817),
            .I(N__43814));
    Odrv4 I__10375 (
            .O(N__43814),
            .I(\c0.data_out_6__1__N_849 ));
    InMux I__10374 (
            .O(N__43811),
            .I(N__43807));
    InMux I__10373 (
            .O(N__43810),
            .I(N__43804));
    LocalMux I__10372 (
            .O(N__43807),
            .I(N__43798));
    LocalMux I__10371 (
            .O(N__43804),
            .I(N__43798));
    InMux I__10370 (
            .O(N__43803),
            .I(N__43793));
    Span4Mux_v I__10369 (
            .O(N__43798),
            .I(N__43790));
    InMux I__10368 (
            .O(N__43797),
            .I(N__43787));
    InMux I__10367 (
            .O(N__43796),
            .I(N__43784));
    LocalMux I__10366 (
            .O(N__43793),
            .I(N__43777));
    Span4Mux_v I__10365 (
            .O(N__43790),
            .I(N__43777));
    LocalMux I__10364 (
            .O(N__43787),
            .I(N__43777));
    LocalMux I__10363 (
            .O(N__43784),
            .I(\c0.data_out_1_1 ));
    Odrv4 I__10362 (
            .O(N__43777),
            .I(\c0.data_out_1_1 ));
    InMux I__10361 (
            .O(N__43772),
            .I(N__43766));
    CascadeMux I__10360 (
            .O(N__43771),
            .I(N__43763));
    CascadeMux I__10359 (
            .O(N__43770),
            .I(N__43760));
    InMux I__10358 (
            .O(N__43769),
            .I(N__43757));
    LocalMux I__10357 (
            .O(N__43766),
            .I(N__43754));
    InMux I__10356 (
            .O(N__43763),
            .I(N__43751));
    InMux I__10355 (
            .O(N__43760),
            .I(N__43746));
    LocalMux I__10354 (
            .O(N__43757),
            .I(N__43743));
    Span4Mux_h I__10353 (
            .O(N__43754),
            .I(N__43738));
    LocalMux I__10352 (
            .O(N__43751),
            .I(N__43738));
    InMux I__10351 (
            .O(N__43750),
            .I(N__43733));
    InMux I__10350 (
            .O(N__43749),
            .I(N__43733));
    LocalMux I__10349 (
            .O(N__43746),
            .I(N__43726));
    Span4Mux_v I__10348 (
            .O(N__43743),
            .I(N__43726));
    Span4Mux_v I__10347 (
            .O(N__43738),
            .I(N__43726));
    LocalMux I__10346 (
            .O(N__43733),
            .I(data_out_1_2));
    Odrv4 I__10345 (
            .O(N__43726),
            .I(data_out_1_2));
    CascadeMux I__10344 (
            .O(N__43721),
            .I(\c0.n8767_cascade_ ));
    InMux I__10343 (
            .O(N__43718),
            .I(N__43715));
    LocalMux I__10342 (
            .O(N__43715),
            .I(N__43712));
    Odrv4 I__10341 (
            .O(N__43712),
            .I(\c0.n17525 ));
    InMux I__10340 (
            .O(N__43709),
            .I(N__43705));
    InMux I__10339 (
            .O(N__43708),
            .I(N__43702));
    LocalMux I__10338 (
            .O(N__43705),
            .I(N__43699));
    LocalMux I__10337 (
            .O(N__43702),
            .I(N__43696));
    Span4Mux_v I__10336 (
            .O(N__43699),
            .I(N__43693));
    Span4Mux_h I__10335 (
            .O(N__43696),
            .I(N__43690));
    Sp12to4 I__10334 (
            .O(N__43693),
            .I(N__43687));
    Odrv4 I__10333 (
            .O(N__43690),
            .I(\c0.n17641 ));
    Odrv12 I__10332 (
            .O(N__43687),
            .I(\c0.n17641 ));
    CascadeMux I__10331 (
            .O(N__43682),
            .I(\c0.n17457_cascade_ ));
    InMux I__10330 (
            .O(N__43679),
            .I(N__43676));
    LocalMux I__10329 (
            .O(N__43676),
            .I(N__43673));
    Span4Mux_h I__10328 (
            .O(N__43673),
            .I(N__43669));
    InMux I__10327 (
            .O(N__43672),
            .I(N__43666));
    Odrv4 I__10326 (
            .O(N__43669),
            .I(\c0.n8964 ));
    LocalMux I__10325 (
            .O(N__43666),
            .I(\c0.n8964 ));
    InMux I__10324 (
            .O(N__43661),
            .I(N__43658));
    LocalMux I__10323 (
            .O(N__43658),
            .I(\c0.n17415 ));
    InMux I__10322 (
            .O(N__43655),
            .I(N__43652));
    LocalMux I__10321 (
            .O(N__43652),
            .I(N__43643));
    InMux I__10320 (
            .O(N__43651),
            .I(N__43640));
    InMux I__10319 (
            .O(N__43650),
            .I(N__43637));
    InMux I__10318 (
            .O(N__43649),
            .I(N__43634));
    InMux I__10317 (
            .O(N__43648),
            .I(N__43631));
    InMux I__10316 (
            .O(N__43647),
            .I(N__43628));
    InMux I__10315 (
            .O(N__43646),
            .I(N__43625));
    Span4Mux_h I__10314 (
            .O(N__43643),
            .I(N__43620));
    LocalMux I__10313 (
            .O(N__43640),
            .I(N__43620));
    LocalMux I__10312 (
            .O(N__43637),
            .I(N__43617));
    LocalMux I__10311 (
            .O(N__43634),
            .I(N__43614));
    LocalMux I__10310 (
            .O(N__43631),
            .I(N__43607));
    LocalMux I__10309 (
            .O(N__43628),
            .I(N__43607));
    LocalMux I__10308 (
            .O(N__43625),
            .I(N__43607));
    Span4Mux_h I__10307 (
            .O(N__43620),
            .I(N__43604));
    Span4Mux_h I__10306 (
            .O(N__43617),
            .I(N__43601));
    Odrv12 I__10305 (
            .O(N__43614),
            .I(\c0.data_out_6__3__N_788 ));
    Odrv12 I__10304 (
            .O(N__43607),
            .I(\c0.data_out_6__3__N_788 ));
    Odrv4 I__10303 (
            .O(N__43604),
            .I(\c0.data_out_6__3__N_788 ));
    Odrv4 I__10302 (
            .O(N__43601),
            .I(\c0.data_out_6__3__N_788 ));
    CascadeMux I__10301 (
            .O(N__43592),
            .I(\c0.n17415_cascade_ ));
    InMux I__10300 (
            .O(N__43589),
            .I(N__43585));
    InMux I__10299 (
            .O(N__43588),
            .I(N__43581));
    LocalMux I__10298 (
            .O(N__43585),
            .I(N__43577));
    InMux I__10297 (
            .O(N__43584),
            .I(N__43574));
    LocalMux I__10296 (
            .O(N__43581),
            .I(N__43571));
    InMux I__10295 (
            .O(N__43580),
            .I(N__43568));
    Span4Mux_v I__10294 (
            .O(N__43577),
            .I(N__43563));
    LocalMux I__10293 (
            .O(N__43574),
            .I(N__43563));
    Span4Mux_h I__10292 (
            .O(N__43571),
            .I(N__43558));
    LocalMux I__10291 (
            .O(N__43568),
            .I(N__43555));
    Span4Mux_h I__10290 (
            .O(N__43563),
            .I(N__43552));
    InMux I__10289 (
            .O(N__43562),
            .I(N__43549));
    InMux I__10288 (
            .O(N__43561),
            .I(N__43546));
    Span4Mux_v I__10287 (
            .O(N__43558),
            .I(N__43543));
    Odrv4 I__10286 (
            .O(N__43555),
            .I(\c0.data_out_5_2 ));
    Odrv4 I__10285 (
            .O(N__43552),
            .I(\c0.data_out_5_2 ));
    LocalMux I__10284 (
            .O(N__43549),
            .I(\c0.data_out_5_2 ));
    LocalMux I__10283 (
            .O(N__43546),
            .I(\c0.data_out_5_2 ));
    Odrv4 I__10282 (
            .O(N__43543),
            .I(\c0.data_out_5_2 ));
    InMux I__10281 (
            .O(N__43532),
            .I(N__43529));
    LocalMux I__10280 (
            .O(N__43529),
            .I(N__43524));
    InMux I__10279 (
            .O(N__43528),
            .I(N__43521));
    InMux I__10278 (
            .O(N__43527),
            .I(N__43518));
    Span4Mux_h I__10277 (
            .O(N__43524),
            .I(N__43515));
    LocalMux I__10276 (
            .O(N__43521),
            .I(N__43512));
    LocalMux I__10275 (
            .O(N__43518),
            .I(N__43509));
    Span4Mux_v I__10274 (
            .O(N__43515),
            .I(N__43502));
    Span4Mux_h I__10273 (
            .O(N__43512),
            .I(N__43502));
    Span4Mux_h I__10272 (
            .O(N__43509),
            .I(N__43502));
    Odrv4 I__10271 (
            .O(N__43502),
            .I(\c0.data_out_6_7 ));
    InMux I__10270 (
            .O(N__43499),
            .I(N__43496));
    LocalMux I__10269 (
            .O(N__43496),
            .I(\c0.n9195 ));
    CascadeMux I__10268 (
            .O(N__43493),
            .I(\c0.n17668_cascade_ ));
    InMux I__10267 (
            .O(N__43490),
            .I(N__43487));
    LocalMux I__10266 (
            .O(N__43487),
            .I(N__43483));
    InMux I__10265 (
            .O(N__43486),
            .I(N__43480));
    Odrv4 I__10264 (
            .O(N__43483),
            .I(\c0.n8812 ));
    LocalMux I__10263 (
            .O(N__43480),
            .I(\c0.n8812 ));
    CascadeMux I__10262 (
            .O(N__43475),
            .I(\c0.n8_adj_2511_cascade_ ));
    InMux I__10261 (
            .O(N__43472),
            .I(N__43469));
    LocalMux I__10260 (
            .O(N__43469),
            .I(\c0.n17623 ));
    InMux I__10259 (
            .O(N__43466),
            .I(N__43462));
    InMux I__10258 (
            .O(N__43465),
            .I(N__43458));
    LocalMux I__10257 (
            .O(N__43462),
            .I(N__43455));
    InMux I__10256 (
            .O(N__43461),
            .I(N__43452));
    LocalMux I__10255 (
            .O(N__43458),
            .I(N__43449));
    Span4Mux_h I__10254 (
            .O(N__43455),
            .I(N__43446));
    LocalMux I__10253 (
            .O(N__43452),
            .I(\c0.n8950 ));
    Odrv4 I__10252 (
            .O(N__43449),
            .I(\c0.n8950 ));
    Odrv4 I__10251 (
            .O(N__43446),
            .I(\c0.n8950 ));
    InMux I__10250 (
            .O(N__43439),
            .I(N__43436));
    LocalMux I__10249 (
            .O(N__43436),
            .I(\c0.data_out_9_0 ));
    InMux I__10248 (
            .O(N__43433),
            .I(N__43430));
    LocalMux I__10247 (
            .O(N__43430),
            .I(\c0.data_out_10_0 ));
    InMux I__10246 (
            .O(N__43427),
            .I(N__43424));
    LocalMux I__10245 (
            .O(N__43424),
            .I(\c0.n18016 ));
    CascadeMux I__10244 (
            .O(N__43421),
            .I(N__43417));
    InMux I__10243 (
            .O(N__43420),
            .I(N__43414));
    InMux I__10242 (
            .O(N__43417),
            .I(N__43410));
    LocalMux I__10241 (
            .O(N__43414),
            .I(N__43404));
    InMux I__10240 (
            .O(N__43413),
            .I(N__43401));
    LocalMux I__10239 (
            .O(N__43410),
            .I(N__43398));
    CascadeMux I__10238 (
            .O(N__43409),
            .I(N__43395));
    InMux I__10237 (
            .O(N__43408),
            .I(N__43391));
    InMux I__10236 (
            .O(N__43407),
            .I(N__43388));
    Span4Mux_v I__10235 (
            .O(N__43404),
            .I(N__43385));
    LocalMux I__10234 (
            .O(N__43401),
            .I(N__43380));
    Span4Mux_h I__10233 (
            .O(N__43398),
            .I(N__43380));
    InMux I__10232 (
            .O(N__43395),
            .I(N__43375));
    InMux I__10231 (
            .O(N__43394),
            .I(N__43375));
    LocalMux I__10230 (
            .O(N__43391),
            .I(N__43370));
    LocalMux I__10229 (
            .O(N__43388),
            .I(N__43370));
    Odrv4 I__10228 (
            .O(N__43385),
            .I(\c0.data_out_2_3 ));
    Odrv4 I__10227 (
            .O(N__43380),
            .I(\c0.data_out_2_3 ));
    LocalMux I__10226 (
            .O(N__43375),
            .I(\c0.data_out_2_3 ));
    Odrv12 I__10225 (
            .O(N__43370),
            .I(\c0.data_out_2_3 ));
    CascadeMux I__10224 (
            .O(N__43361),
            .I(\c0.n4_adj_2543_cascade_ ));
    CascadeMux I__10223 (
            .O(N__43358),
            .I(\c0.n18073_cascade_ ));
    InMux I__10222 (
            .O(N__43355),
            .I(N__43352));
    LocalMux I__10221 (
            .O(N__43352),
            .I(N__43348));
    CascadeMux I__10220 (
            .O(N__43351),
            .I(N__43345));
    Span12Mux_h I__10219 (
            .O(N__43348),
            .I(N__43342));
    InMux I__10218 (
            .O(N__43345),
            .I(N__43339));
    Odrv12 I__10217 (
            .O(N__43342),
            .I(rand_setpoint_3));
    LocalMux I__10216 (
            .O(N__43339),
            .I(rand_setpoint_3));
    InMux I__10215 (
            .O(N__43334),
            .I(N__43329));
    InMux I__10214 (
            .O(N__43333),
            .I(N__43325));
    InMux I__10213 (
            .O(N__43332),
            .I(N__43322));
    LocalMux I__10212 (
            .O(N__43329),
            .I(N__43319));
    InMux I__10211 (
            .O(N__43328),
            .I(N__43316));
    LocalMux I__10210 (
            .O(N__43325),
            .I(N__43313));
    LocalMux I__10209 (
            .O(N__43322),
            .I(N__43308));
    Span4Mux_h I__10208 (
            .O(N__43319),
            .I(N__43308));
    LocalMux I__10207 (
            .O(N__43316),
            .I(data_out_8_2));
    Odrv12 I__10206 (
            .O(N__43313),
            .I(data_out_8_2));
    Odrv4 I__10205 (
            .O(N__43308),
            .I(data_out_8_2));
    InMux I__10204 (
            .O(N__43301),
            .I(N__43297));
    InMux I__10203 (
            .O(N__43300),
            .I(N__43294));
    LocalMux I__10202 (
            .O(N__43297),
            .I(N__43291));
    LocalMux I__10201 (
            .O(N__43294),
            .I(N__43288));
    Span4Mux_h I__10200 (
            .O(N__43291),
            .I(N__43285));
    Odrv12 I__10199 (
            .O(N__43288),
            .I(\c0.data_out_6_4 ));
    Odrv4 I__10198 (
            .O(N__43285),
            .I(\c0.data_out_6_4 ));
    CascadeMux I__10197 (
            .O(N__43280),
            .I(\c0.n9091_cascade_ ));
    CascadeMux I__10196 (
            .O(N__43277),
            .I(\c0.n17566_cascade_ ));
    InMux I__10195 (
            .O(N__43274),
            .I(N__43271));
    LocalMux I__10194 (
            .O(N__43271),
            .I(N__43266));
    InMux I__10193 (
            .O(N__43270),
            .I(N__43263));
    InMux I__10192 (
            .O(N__43269),
            .I(N__43260));
    Span4Mux_h I__10191 (
            .O(N__43266),
            .I(N__43257));
    LocalMux I__10190 (
            .O(N__43263),
            .I(N__43254));
    LocalMux I__10189 (
            .O(N__43260),
            .I(N__43251));
    Span4Mux_v I__10188 (
            .O(N__43257),
            .I(N__43248));
    Span4Mux_h I__10187 (
            .O(N__43254),
            .I(N__43245));
    Span4Mux_v I__10186 (
            .O(N__43251),
            .I(N__43242));
    Odrv4 I__10185 (
            .O(N__43248),
            .I(\c0.data_out_6_3 ));
    Odrv4 I__10184 (
            .O(N__43245),
            .I(\c0.data_out_6_3 ));
    Odrv4 I__10183 (
            .O(N__43242),
            .I(\c0.data_out_6_3 ));
    CascadeMux I__10182 (
            .O(N__43235),
            .I(\c0.n9195_cascade_ ));
    InMux I__10181 (
            .O(N__43232),
            .I(N__43227));
    InMux I__10180 (
            .O(N__43231),
            .I(N__43223));
    InMux I__10179 (
            .O(N__43230),
            .I(N__43220));
    LocalMux I__10178 (
            .O(N__43227),
            .I(N__43217));
    InMux I__10177 (
            .O(N__43226),
            .I(N__43214));
    LocalMux I__10176 (
            .O(N__43223),
            .I(N__43211));
    LocalMux I__10175 (
            .O(N__43220),
            .I(\c0.data_out_7__4__N_556 ));
    Odrv4 I__10174 (
            .O(N__43217),
            .I(\c0.data_out_7__4__N_556 ));
    LocalMux I__10173 (
            .O(N__43214),
            .I(\c0.data_out_7__4__N_556 ));
    Odrv12 I__10172 (
            .O(N__43211),
            .I(\c0.data_out_7__4__N_556 ));
    InMux I__10171 (
            .O(N__43202),
            .I(N__43199));
    LocalMux I__10170 (
            .O(N__43199),
            .I(N__43196));
    Span4Mux_h I__10169 (
            .O(N__43196),
            .I(N__43193));
    Odrv4 I__10168 (
            .O(N__43193),
            .I(\c0.n18015 ));
    CascadeMux I__10167 (
            .O(N__43190),
            .I(N__43187));
    InMux I__10166 (
            .O(N__43187),
            .I(N__43184));
    LocalMux I__10165 (
            .O(N__43184),
            .I(\c0.n8_adj_2516 ));
    InMux I__10164 (
            .O(N__43181),
            .I(N__43177));
    InMux I__10163 (
            .O(N__43180),
            .I(N__43174));
    LocalMux I__10162 (
            .O(N__43177),
            .I(N__43171));
    LocalMux I__10161 (
            .O(N__43174),
            .I(r_Tx_Data_1));
    Odrv12 I__10160 (
            .O(N__43171),
            .I(r_Tx_Data_1));
    InMux I__10159 (
            .O(N__43166),
            .I(N__43163));
    LocalMux I__10158 (
            .O(N__43163),
            .I(\c0.n18071 ));
    CascadeMux I__10157 (
            .O(N__43160),
            .I(\c0.n8_adj_2526_cascade_ ));
    InMux I__10156 (
            .O(N__43157),
            .I(N__43154));
    LocalMux I__10155 (
            .O(N__43154),
            .I(N__43151));
    Span4Mux_h I__10154 (
            .O(N__43151),
            .I(N__43148));
    Odrv4 I__10153 (
            .O(N__43148),
            .I(\c0.n18072 ));
    CascadeMux I__10152 (
            .O(N__43145),
            .I(N__43142));
    InMux I__10151 (
            .O(N__43142),
            .I(N__43139));
    LocalMux I__10150 (
            .O(N__43139),
            .I(N__43136));
    Span4Mux_v I__10149 (
            .O(N__43136),
            .I(N__43133));
    Span4Mux_h I__10148 (
            .O(N__43133),
            .I(N__43129));
    InMux I__10147 (
            .O(N__43132),
            .I(N__43126));
    Odrv4 I__10146 (
            .O(N__43129),
            .I(\c0.n17644 ));
    LocalMux I__10145 (
            .O(N__43126),
            .I(\c0.n17644 ));
    InMux I__10144 (
            .O(N__43121),
            .I(N__43118));
    LocalMux I__10143 (
            .O(N__43118),
            .I(N__43115));
    Span4Mux_v I__10142 (
            .O(N__43115),
            .I(N__43112));
    Odrv4 I__10141 (
            .O(N__43112),
            .I(\c0.data_out_7__2__N_574 ));
    CascadeMux I__10140 (
            .O(N__43109),
            .I(\c0.data_out_7__2__N_574_cascade_ ));
    InMux I__10139 (
            .O(N__43106),
            .I(N__43103));
    LocalMux I__10138 (
            .O(N__43103),
            .I(\c0.data_out_10_2 ));
    InMux I__10137 (
            .O(N__43100),
            .I(N__43097));
    LocalMux I__10136 (
            .O(N__43097),
            .I(\c0.data_out_9_2 ));
    InMux I__10135 (
            .O(N__43094),
            .I(N__43091));
    LocalMux I__10134 (
            .O(N__43091),
            .I(N__43088));
    Span4Mux_h I__10133 (
            .O(N__43088),
            .I(N__43085));
    Span4Mux_h I__10132 (
            .O(N__43085),
            .I(N__43082));
    Odrv4 I__10131 (
            .O(N__43082),
            .I(\c0.data_out_9_3 ));
    InMux I__10130 (
            .O(N__43079),
            .I(N__43076));
    LocalMux I__10129 (
            .O(N__43076),
            .I(\c0.n2650 ));
    InMux I__10128 (
            .O(N__43073),
            .I(N__43070));
    LocalMux I__10127 (
            .O(N__43070),
            .I(N__43065));
    InMux I__10126 (
            .O(N__43069),
            .I(N__43062));
    InMux I__10125 (
            .O(N__43068),
            .I(N__43059));
    Odrv4 I__10124 (
            .O(N__43065),
            .I(\c0.tx_transmit_N_2239_0 ));
    LocalMux I__10123 (
            .O(N__43062),
            .I(\c0.tx_transmit_N_2239_0 ));
    LocalMux I__10122 (
            .O(N__43059),
            .I(\c0.tx_transmit_N_2239_0 ));
    InMux I__10121 (
            .O(N__43052),
            .I(N__43047));
    InMux I__10120 (
            .O(N__43051),
            .I(N__43044));
    InMux I__10119 (
            .O(N__43050),
            .I(N__43041));
    LocalMux I__10118 (
            .O(N__43047),
            .I(\c0.tx_transmit_N_2239_1 ));
    LocalMux I__10117 (
            .O(N__43044),
            .I(\c0.tx_transmit_N_2239_1 ));
    LocalMux I__10116 (
            .O(N__43041),
            .I(\c0.tx_transmit_N_2239_1 ));
    InMux I__10115 (
            .O(N__43034),
            .I(N__43031));
    LocalMux I__10114 (
            .O(N__43031),
            .I(N__43028));
    Span4Mux_h I__10113 (
            .O(N__43028),
            .I(N__43023));
    InMux I__10112 (
            .O(N__43027),
            .I(N__43020));
    InMux I__10111 (
            .O(N__43026),
            .I(N__43017));
    Odrv4 I__10110 (
            .O(N__43023),
            .I(tx_transmit_N_2239_2));
    LocalMux I__10109 (
            .O(N__43020),
            .I(tx_transmit_N_2239_2));
    LocalMux I__10108 (
            .O(N__43017),
            .I(tx_transmit_N_2239_2));
    InMux I__10107 (
            .O(N__43010),
            .I(N__43007));
    LocalMux I__10106 (
            .O(N__43007),
            .I(N__43003));
    InMux I__10105 (
            .O(N__43006),
            .I(N__42999));
    Span4Mux_v I__10104 (
            .O(N__43003),
            .I(N__42996));
    InMux I__10103 (
            .O(N__43002),
            .I(N__42993));
    LocalMux I__10102 (
            .O(N__42999),
            .I(\c0.n97 ));
    Odrv4 I__10101 (
            .O(N__42996),
            .I(\c0.n97 ));
    LocalMux I__10100 (
            .O(N__42993),
            .I(\c0.n97 ));
    CascadeMux I__10099 (
            .O(N__42986),
            .I(N__42980));
    CascadeMux I__10098 (
            .O(N__42985),
            .I(N__42976));
    InMux I__10097 (
            .O(N__42984),
            .I(N__42971));
    InMux I__10096 (
            .O(N__42983),
            .I(N__42971));
    InMux I__10095 (
            .O(N__42980),
            .I(N__42968));
    InMux I__10094 (
            .O(N__42979),
            .I(N__42965));
    InMux I__10093 (
            .O(N__42976),
            .I(N__42962));
    LocalMux I__10092 (
            .O(N__42971),
            .I(N__42959));
    LocalMux I__10091 (
            .O(N__42968),
            .I(N__42956));
    LocalMux I__10090 (
            .O(N__42965),
            .I(N__42951));
    LocalMux I__10089 (
            .O(N__42962),
            .I(N__42951));
    Span4Mux_v I__10088 (
            .O(N__42959),
            .I(N__42947));
    Span12Mux_h I__10087 (
            .O(N__42956),
            .I(N__42942));
    Span12Mux_h I__10086 (
            .O(N__42951),
            .I(N__42942));
    InMux I__10085 (
            .O(N__42950),
            .I(N__42939));
    Odrv4 I__10084 (
            .O(N__42947),
            .I(\c0.tx_transmit ));
    Odrv12 I__10083 (
            .O(N__42942),
            .I(\c0.tx_transmit ));
    LocalMux I__10082 (
            .O(N__42939),
            .I(\c0.tx_transmit ));
    InMux I__10081 (
            .O(N__42932),
            .I(N__42927));
    InMux I__10080 (
            .O(N__42931),
            .I(N__42924));
    InMux I__10079 (
            .O(N__42930),
            .I(N__42921));
    LocalMux I__10078 (
            .O(N__42927),
            .I(N__42916));
    LocalMux I__10077 (
            .O(N__42924),
            .I(N__42916));
    LocalMux I__10076 (
            .O(N__42921),
            .I(N__42910));
    Span4Mux_v I__10075 (
            .O(N__42916),
            .I(N__42907));
    InMux I__10074 (
            .O(N__42915),
            .I(N__42900));
    InMux I__10073 (
            .O(N__42914),
            .I(N__42900));
    InMux I__10072 (
            .O(N__42913),
            .I(N__42900));
    Odrv4 I__10071 (
            .O(N__42910),
            .I(tx_active));
    Odrv4 I__10070 (
            .O(N__42907),
            .I(tx_active));
    LocalMux I__10069 (
            .O(N__42900),
            .I(tx_active));
    CascadeMux I__10068 (
            .O(N__42893),
            .I(N__42889));
    CascadeMux I__10067 (
            .O(N__42892),
            .I(N__42885));
    InMux I__10066 (
            .O(N__42889),
            .I(N__42881));
    InMux I__10065 (
            .O(N__42888),
            .I(N__42878));
    InMux I__10064 (
            .O(N__42885),
            .I(N__42875));
    InMux I__10063 (
            .O(N__42884),
            .I(N__42871));
    LocalMux I__10062 (
            .O(N__42881),
            .I(N__42867));
    LocalMux I__10061 (
            .O(N__42878),
            .I(N__42862));
    LocalMux I__10060 (
            .O(N__42875),
            .I(N__42862));
    InMux I__10059 (
            .O(N__42874),
            .I(N__42859));
    LocalMux I__10058 (
            .O(N__42871),
            .I(N__42856));
    InMux I__10057 (
            .O(N__42870),
            .I(N__42853));
    Span4Mux_v I__10056 (
            .O(N__42867),
            .I(N__42848));
    Span4Mux_v I__10055 (
            .O(N__42862),
            .I(N__42848));
    LocalMux I__10054 (
            .O(N__42859),
            .I(n13415));
    Odrv4 I__10053 (
            .O(N__42856),
            .I(n13415));
    LocalMux I__10052 (
            .O(N__42853),
            .I(n13415));
    Odrv4 I__10051 (
            .O(N__42848),
            .I(n13415));
    InMux I__10050 (
            .O(N__42839),
            .I(N__42833));
    InMux I__10049 (
            .O(N__42838),
            .I(N__42830));
    InMux I__10048 (
            .O(N__42837),
            .I(N__42824));
    InMux I__10047 (
            .O(N__42836),
            .I(N__42821));
    LocalMux I__10046 (
            .O(N__42833),
            .I(N__42818));
    LocalMux I__10045 (
            .O(N__42830),
            .I(N__42815));
    InMux I__10044 (
            .O(N__42829),
            .I(N__42808));
    InMux I__10043 (
            .O(N__42828),
            .I(N__42808));
    InMux I__10042 (
            .O(N__42827),
            .I(N__42808));
    LocalMux I__10041 (
            .O(N__42824),
            .I(tx_transmit_N_2239_3));
    LocalMux I__10040 (
            .O(N__42821),
            .I(tx_transmit_N_2239_3));
    Odrv12 I__10039 (
            .O(N__42818),
            .I(tx_transmit_N_2239_3));
    Odrv4 I__10038 (
            .O(N__42815),
            .I(tx_transmit_N_2239_3));
    LocalMux I__10037 (
            .O(N__42808),
            .I(tx_transmit_N_2239_3));
    CascadeMux I__10036 (
            .O(N__42797),
            .I(N__42794));
    InMux I__10035 (
            .O(N__42794),
            .I(N__42790));
    InMux I__10034 (
            .O(N__42793),
            .I(N__42787));
    LocalMux I__10033 (
            .O(N__42790),
            .I(N__42784));
    LocalMux I__10032 (
            .O(N__42787),
            .I(r_Tx_Data_5));
    Odrv12 I__10031 (
            .O(N__42784),
            .I(r_Tx_Data_5));
    InMux I__10030 (
            .O(N__42779),
            .I(N__42775));
    InMux I__10029 (
            .O(N__42778),
            .I(N__42772));
    LocalMux I__10028 (
            .O(N__42775),
            .I(N__42769));
    LocalMux I__10027 (
            .O(N__42772),
            .I(n16485));
    Odrv4 I__10026 (
            .O(N__42769),
            .I(n16485));
    CascadeMux I__10025 (
            .O(N__42764),
            .I(N__42761));
    InMux I__10024 (
            .O(N__42761),
            .I(N__42758));
    LocalMux I__10023 (
            .O(N__42758),
            .I(N__42755));
    Span4Mux_h I__10022 (
            .O(N__42755),
            .I(N__42752));
    Odrv4 I__10021 (
            .O(N__42752),
            .I(\c0.n7428 ));
    InMux I__10020 (
            .O(N__42749),
            .I(N__42746));
    LocalMux I__10019 (
            .O(N__42746),
            .I(N__42741));
    InMux I__10018 (
            .O(N__42745),
            .I(N__42736));
    InMux I__10017 (
            .O(N__42744),
            .I(N__42736));
    Sp12to4 I__10016 (
            .O(N__42741),
            .I(N__42731));
    LocalMux I__10015 (
            .O(N__42736),
            .I(N__42731));
    Span12Mux_s7_v I__10014 (
            .O(N__42731),
            .I(N__42726));
    InMux I__10013 (
            .O(N__42730),
            .I(N__42723));
    InMux I__10012 (
            .O(N__42729),
            .I(N__42720));
    Odrv12 I__10011 (
            .O(N__42726),
            .I(n14_adj_2615));
    LocalMux I__10010 (
            .O(N__42723),
            .I(n14_adj_2615));
    LocalMux I__10009 (
            .O(N__42720),
            .I(n14_adj_2615));
    CascadeMux I__10008 (
            .O(N__42713),
            .I(N__42709));
    InMux I__10007 (
            .O(N__42712),
            .I(N__42701));
    InMux I__10006 (
            .O(N__42709),
            .I(N__42701));
    CascadeMux I__10005 (
            .O(N__42708),
            .I(N__42698));
    CascadeMux I__10004 (
            .O(N__42707),
            .I(N__42693));
    InMux I__10003 (
            .O(N__42706),
            .I(N__42689));
    LocalMux I__10002 (
            .O(N__42701),
            .I(N__42686));
    InMux I__10001 (
            .O(N__42698),
            .I(N__42683));
    InMux I__10000 (
            .O(N__42697),
            .I(N__42678));
    InMux I__9999 (
            .O(N__42696),
            .I(N__42678));
    InMux I__9998 (
            .O(N__42693),
            .I(N__42675));
    CascadeMux I__9997 (
            .O(N__42692),
            .I(N__42672));
    LocalMux I__9996 (
            .O(N__42689),
            .I(N__42669));
    Span4Mux_h I__9995 (
            .O(N__42686),
            .I(N__42660));
    LocalMux I__9994 (
            .O(N__42683),
            .I(N__42660));
    LocalMux I__9993 (
            .O(N__42678),
            .I(N__42660));
    LocalMux I__9992 (
            .O(N__42675),
            .I(N__42660));
    InMux I__9991 (
            .O(N__42672),
            .I(N__42657));
    Span4Mux_v I__9990 (
            .O(N__42669),
            .I(N__42653));
    Span4Mux_v I__9989 (
            .O(N__42660),
            .I(N__42650));
    LocalMux I__9988 (
            .O(N__42657),
            .I(N__42647));
    InMux I__9987 (
            .O(N__42656),
            .I(N__42644));
    Odrv4 I__9986 (
            .O(N__42653),
            .I(n9631));
    Odrv4 I__9985 (
            .O(N__42650),
            .I(n9631));
    Odrv4 I__9984 (
            .O(N__42647),
            .I(n9631));
    LocalMux I__9983 (
            .O(N__42644),
            .I(n9631));
    CascadeMux I__9982 (
            .O(N__42635),
            .I(N__42632));
    InMux I__9981 (
            .O(N__42632),
            .I(N__42629));
    LocalMux I__9980 (
            .O(N__42629),
            .I(N__42625));
    InMux I__9979 (
            .O(N__42628),
            .I(N__42622));
    Odrv4 I__9978 (
            .O(N__42625),
            .I(tx_transmit_N_2239_6));
    LocalMux I__9977 (
            .O(N__42622),
            .I(tx_transmit_N_2239_6));
    CascadeMux I__9976 (
            .O(N__42617),
            .I(N__42613));
    InMux I__9975 (
            .O(N__42616),
            .I(N__42610));
    InMux I__9974 (
            .O(N__42613),
            .I(N__42607));
    LocalMux I__9973 (
            .O(N__42610),
            .I(byte_transmit_counter_6));
    LocalMux I__9972 (
            .O(N__42607),
            .I(byte_transmit_counter_6));
    InMux I__9971 (
            .O(N__42602),
            .I(N__42598));
    InMux I__9970 (
            .O(N__42601),
            .I(N__42595));
    LocalMux I__9969 (
            .O(N__42598),
            .I(\c0.n149 ));
    LocalMux I__9968 (
            .O(N__42595),
            .I(\c0.n149 ));
    CascadeMux I__9967 (
            .O(N__42590),
            .I(N__42587));
    InMux I__9966 (
            .O(N__42587),
            .I(N__42584));
    LocalMux I__9965 (
            .O(N__42584),
            .I(\c0.n17741 ));
    CascadeMux I__9964 (
            .O(N__42581),
            .I(N__42576));
    CascadeMux I__9963 (
            .O(N__42580),
            .I(N__42563));
    InMux I__9962 (
            .O(N__42579),
            .I(N__42556));
    InMux I__9961 (
            .O(N__42576),
            .I(N__42556));
    InMux I__9960 (
            .O(N__42575),
            .I(N__42546));
    InMux I__9959 (
            .O(N__42574),
            .I(N__42546));
    InMux I__9958 (
            .O(N__42573),
            .I(N__42541));
    InMux I__9957 (
            .O(N__42572),
            .I(N__42541));
    InMux I__9956 (
            .O(N__42571),
            .I(N__42538));
    InMux I__9955 (
            .O(N__42570),
            .I(N__42535));
    InMux I__9954 (
            .O(N__42569),
            .I(N__42532));
    InMux I__9953 (
            .O(N__42568),
            .I(N__42529));
    InMux I__9952 (
            .O(N__42567),
            .I(N__42526));
    InMux I__9951 (
            .O(N__42566),
            .I(N__42521));
    InMux I__9950 (
            .O(N__42563),
            .I(N__42521));
    InMux I__9949 (
            .O(N__42562),
            .I(N__42516));
    InMux I__9948 (
            .O(N__42561),
            .I(N__42516));
    LocalMux I__9947 (
            .O(N__42556),
            .I(N__42513));
    InMux I__9946 (
            .O(N__42555),
            .I(N__42510));
    InMux I__9945 (
            .O(N__42554),
            .I(N__42507));
    InMux I__9944 (
            .O(N__42553),
            .I(N__42504));
    InMux I__9943 (
            .O(N__42552),
            .I(N__42499));
    InMux I__9942 (
            .O(N__42551),
            .I(N__42499));
    LocalMux I__9941 (
            .O(N__42546),
            .I(N__42496));
    LocalMux I__9940 (
            .O(N__42541),
            .I(N__42493));
    LocalMux I__9939 (
            .O(N__42538),
            .I(N__42488));
    LocalMux I__9938 (
            .O(N__42535),
            .I(N__42488));
    LocalMux I__9937 (
            .O(N__42532),
            .I(n29));
    LocalMux I__9936 (
            .O(N__42529),
            .I(n29));
    LocalMux I__9935 (
            .O(N__42526),
            .I(n29));
    LocalMux I__9934 (
            .O(N__42521),
            .I(n29));
    LocalMux I__9933 (
            .O(N__42516),
            .I(n29));
    Odrv4 I__9932 (
            .O(N__42513),
            .I(n29));
    LocalMux I__9931 (
            .O(N__42510),
            .I(n29));
    LocalMux I__9930 (
            .O(N__42507),
            .I(n29));
    LocalMux I__9929 (
            .O(N__42504),
            .I(n29));
    LocalMux I__9928 (
            .O(N__42499),
            .I(n29));
    Odrv4 I__9927 (
            .O(N__42496),
            .I(n29));
    Odrv4 I__9926 (
            .O(N__42493),
            .I(n29));
    Odrv4 I__9925 (
            .O(N__42488),
            .I(n29));
    CascadeMux I__9924 (
            .O(N__42461),
            .I(N__42458));
    InMux I__9923 (
            .O(N__42458),
            .I(N__42455));
    LocalMux I__9922 (
            .O(N__42455),
            .I(N__42452));
    Odrv4 I__9921 (
            .O(N__42452),
            .I(\c0.n7268 ));
    InMux I__9920 (
            .O(N__42449),
            .I(N__42445));
    InMux I__9919 (
            .O(N__42448),
            .I(N__42442));
    LocalMux I__9918 (
            .O(N__42445),
            .I(N__42439));
    LocalMux I__9917 (
            .O(N__42442),
            .I(N__42424));
    Span4Mux_h I__9916 (
            .O(N__42439),
            .I(N__42421));
    InMux I__9915 (
            .O(N__42438),
            .I(N__42416));
    InMux I__9914 (
            .O(N__42437),
            .I(N__42416));
    InMux I__9913 (
            .O(N__42436),
            .I(N__42407));
    InMux I__9912 (
            .O(N__42435),
            .I(N__42407));
    InMux I__9911 (
            .O(N__42434),
            .I(N__42407));
    InMux I__9910 (
            .O(N__42433),
            .I(N__42407));
    InMux I__9909 (
            .O(N__42432),
            .I(N__42400));
    InMux I__9908 (
            .O(N__42431),
            .I(N__42400));
    InMux I__9907 (
            .O(N__42430),
            .I(N__42400));
    InMux I__9906 (
            .O(N__42429),
            .I(N__42393));
    InMux I__9905 (
            .O(N__42428),
            .I(N__42393));
    InMux I__9904 (
            .O(N__42427),
            .I(N__42393));
    Odrv4 I__9903 (
            .O(N__42424),
            .I(\c0.n1314 ));
    Odrv4 I__9902 (
            .O(N__42421),
            .I(\c0.n1314 ));
    LocalMux I__9901 (
            .O(N__42416),
            .I(\c0.n1314 ));
    LocalMux I__9900 (
            .O(N__42407),
            .I(\c0.n1314 ));
    LocalMux I__9899 (
            .O(N__42400),
            .I(\c0.n1314 ));
    LocalMux I__9898 (
            .O(N__42393),
            .I(\c0.n1314 ));
    InMux I__9897 (
            .O(N__42380),
            .I(N__42376));
    InMux I__9896 (
            .O(N__42379),
            .I(N__42371));
    LocalMux I__9895 (
            .O(N__42376),
            .I(N__42368));
    InMux I__9894 (
            .O(N__42375),
            .I(N__42363));
    InMux I__9893 (
            .O(N__42374),
            .I(N__42363));
    LocalMux I__9892 (
            .O(N__42371),
            .I(\c0.delay_counter_7 ));
    Odrv4 I__9891 (
            .O(N__42368),
            .I(\c0.delay_counter_7 ));
    LocalMux I__9890 (
            .O(N__42363),
            .I(\c0.delay_counter_7 ));
    InMux I__9889 (
            .O(N__42356),
            .I(N__42350));
    InMux I__9888 (
            .O(N__42355),
            .I(N__42347));
    InMux I__9887 (
            .O(N__42354),
            .I(N__42342));
    InMux I__9886 (
            .O(N__42353),
            .I(N__42342));
    LocalMux I__9885 (
            .O(N__42350),
            .I(\c0.delay_counter_11 ));
    LocalMux I__9884 (
            .O(N__42347),
            .I(\c0.delay_counter_11 ));
    LocalMux I__9883 (
            .O(N__42342),
            .I(\c0.delay_counter_11 ));
    InMux I__9882 (
            .O(N__42335),
            .I(N__42330));
    CascadeMux I__9881 (
            .O(N__42334),
            .I(N__42326));
    InMux I__9880 (
            .O(N__42333),
            .I(N__42323));
    LocalMux I__9879 (
            .O(N__42330),
            .I(N__42320));
    InMux I__9878 (
            .O(N__42329),
            .I(N__42315));
    InMux I__9877 (
            .O(N__42326),
            .I(N__42315));
    LocalMux I__9876 (
            .O(N__42323),
            .I(N__42312));
    Span4Mux_h I__9875 (
            .O(N__42320),
            .I(N__42309));
    LocalMux I__9874 (
            .O(N__42315),
            .I(\c0.delay_counter_8 ));
    Odrv4 I__9873 (
            .O(N__42312),
            .I(\c0.delay_counter_8 ));
    Odrv4 I__9872 (
            .O(N__42309),
            .I(\c0.delay_counter_8 ));
    CascadeMux I__9871 (
            .O(N__42302),
            .I(N__42297));
    InMux I__9870 (
            .O(N__42301),
            .I(N__42293));
    InMux I__9869 (
            .O(N__42300),
            .I(N__42290));
    InMux I__9868 (
            .O(N__42297),
            .I(N__42287));
    InMux I__9867 (
            .O(N__42296),
            .I(N__42284));
    LocalMux I__9866 (
            .O(N__42293),
            .I(\c0.delay_counter_5 ));
    LocalMux I__9865 (
            .O(N__42290),
            .I(\c0.delay_counter_5 ));
    LocalMux I__9864 (
            .O(N__42287),
            .I(\c0.delay_counter_5 ));
    LocalMux I__9863 (
            .O(N__42284),
            .I(\c0.delay_counter_5 ));
    CascadeMux I__9862 (
            .O(N__42275),
            .I(\c0.n10_adj_2532_cascade_ ));
    InMux I__9861 (
            .O(N__42272),
            .I(N__42269));
    LocalMux I__9860 (
            .O(N__42269),
            .I(N__42266));
    Odrv4 I__9859 (
            .O(N__42266),
            .I(\c0.n14_adj_2533 ));
    InMux I__9858 (
            .O(N__42263),
            .I(N__42260));
    LocalMux I__9857 (
            .O(N__42260),
            .I(N__42257));
    Span4Mux_v I__9856 (
            .O(N__42257),
            .I(N__42254));
    Odrv4 I__9855 (
            .O(N__42254),
            .I(n17306));
    CascadeMux I__9854 (
            .O(N__42251),
            .I(n17306_cascade_));
    InMux I__9853 (
            .O(N__42248),
            .I(N__42245));
    LocalMux I__9852 (
            .O(N__42245),
            .I(N__42242));
    Span12Mux_s4_v I__9851 (
            .O(N__42242),
            .I(N__42237));
    InMux I__9850 (
            .O(N__42241),
            .I(N__42234));
    InMux I__9849 (
            .O(N__42240),
            .I(N__42231));
    Odrv12 I__9848 (
            .O(N__42237),
            .I(\c0.n17387 ));
    LocalMux I__9847 (
            .O(N__42234),
            .I(\c0.n17387 ));
    LocalMux I__9846 (
            .O(N__42231),
            .I(\c0.n17387 ));
    InMux I__9845 (
            .O(N__42224),
            .I(N__42221));
    LocalMux I__9844 (
            .O(N__42221),
            .I(\c0.n6_adj_2534 ));
    InMux I__9843 (
            .O(N__42218),
            .I(N__42215));
    LocalMux I__9842 (
            .O(N__42215),
            .I(N__42212));
    Span4Mux_h I__9841 (
            .O(N__42212),
            .I(N__42209));
    Odrv4 I__9840 (
            .O(N__42209),
            .I(tx_data_4_N_keep));
    InMux I__9839 (
            .O(N__42206),
            .I(N__42202));
    InMux I__9838 (
            .O(N__42205),
            .I(N__42199));
    LocalMux I__9837 (
            .O(N__42202),
            .I(N__42196));
    LocalMux I__9836 (
            .O(N__42199),
            .I(r_Tx_Data_4));
    Odrv4 I__9835 (
            .O(N__42196),
            .I(r_Tx_Data_4));
    CascadeMux I__9834 (
            .O(N__42191),
            .I(\c0.n16_adj_2445_cascade_ ));
    CascadeMux I__9833 (
            .O(N__42188),
            .I(\c0.n19_adj_2446_cascade_ ));
    InMux I__9832 (
            .O(N__42185),
            .I(N__42180));
    InMux I__9831 (
            .O(N__42184),
            .I(N__42177));
    InMux I__9830 (
            .O(N__42183),
            .I(N__42172));
    LocalMux I__9829 (
            .O(N__42180),
            .I(N__42167));
    LocalMux I__9828 (
            .O(N__42177),
            .I(N__42167));
    InMux I__9827 (
            .O(N__42176),
            .I(N__42162));
    InMux I__9826 (
            .O(N__42175),
            .I(N__42162));
    LocalMux I__9825 (
            .O(N__42172),
            .I(\c0.n8550 ));
    Odrv4 I__9824 (
            .O(N__42167),
            .I(\c0.n8550 ));
    LocalMux I__9823 (
            .O(N__42162),
            .I(\c0.n8550 ));
    InMux I__9822 (
            .O(N__42155),
            .I(N__42151));
    InMux I__9821 (
            .O(N__42154),
            .I(N__42148));
    LocalMux I__9820 (
            .O(N__42151),
            .I(n96));
    LocalMux I__9819 (
            .O(N__42148),
            .I(n96));
    InMux I__9818 (
            .O(N__42143),
            .I(N__42139));
    InMux I__9817 (
            .O(N__42142),
            .I(N__42136));
    LocalMux I__9816 (
            .O(N__42139),
            .I(n6878));
    LocalMux I__9815 (
            .O(N__42136),
            .I(n6878));
    CascadeMux I__9814 (
            .O(N__42131),
            .I(n17672_cascade_));
    InMux I__9813 (
            .O(N__42128),
            .I(N__42123));
    InMux I__9812 (
            .O(N__42127),
            .I(N__42120));
    InMux I__9811 (
            .O(N__42126),
            .I(N__42117));
    LocalMux I__9810 (
            .O(N__42123),
            .I(\c0.n113 ));
    LocalMux I__9809 (
            .O(N__42120),
            .I(\c0.n113 ));
    LocalMux I__9808 (
            .O(N__42117),
            .I(\c0.n113 ));
    InMux I__9807 (
            .O(N__42110),
            .I(N__42103));
    InMux I__9806 (
            .O(N__42109),
            .I(N__42103));
    InMux I__9805 (
            .O(N__42108),
            .I(N__42100));
    LocalMux I__9804 (
            .O(N__42103),
            .I(n17364));
    LocalMux I__9803 (
            .O(N__42100),
            .I(n17364));
    InMux I__9802 (
            .O(N__42095),
            .I(N__42092));
    LocalMux I__9801 (
            .O(N__42092),
            .I(N__42089));
    Span4Mux_h I__9800 (
            .O(N__42089),
            .I(N__42086));
    Odrv4 I__9799 (
            .O(N__42086),
            .I(\c0.n18009 ));
    InMux I__9798 (
            .O(N__42083),
            .I(N__42078));
    InMux I__9797 (
            .O(N__42082),
            .I(N__42075));
    InMux I__9796 (
            .O(N__42081),
            .I(N__42072));
    LocalMux I__9795 (
            .O(N__42078),
            .I(N__42069));
    LocalMux I__9794 (
            .O(N__42075),
            .I(N__42066));
    LocalMux I__9793 (
            .O(N__42072),
            .I(N__42058));
    Span4Mux_h I__9792 (
            .O(N__42069),
            .I(N__42058));
    Span4Mux_v I__9791 (
            .O(N__42066),
            .I(N__42058));
    InMux I__9790 (
            .O(N__42065),
            .I(N__42055));
    Odrv4 I__9789 (
            .O(N__42058),
            .I(\c0.delay_counter_12 ));
    LocalMux I__9788 (
            .O(N__42055),
            .I(\c0.delay_counter_12 ));
    InMux I__9787 (
            .O(N__42050),
            .I(N__42044));
    InMux I__9786 (
            .O(N__42049),
            .I(N__42041));
    InMux I__9785 (
            .O(N__42048),
            .I(N__42038));
    InMux I__9784 (
            .O(N__42047),
            .I(N__42035));
    LocalMux I__9783 (
            .O(N__42044),
            .I(N__42032));
    LocalMux I__9782 (
            .O(N__42041),
            .I(N__42029));
    LocalMux I__9781 (
            .O(N__42038),
            .I(N__42026));
    LocalMux I__9780 (
            .O(N__42035),
            .I(N__42023));
    Odrv12 I__9779 (
            .O(N__42032),
            .I(n119));
    Odrv4 I__9778 (
            .O(N__42029),
            .I(n119));
    Odrv4 I__9777 (
            .O(N__42026),
            .I(n119));
    Odrv12 I__9776 (
            .O(N__42023),
            .I(n119));
    CascadeMux I__9775 (
            .O(N__42014),
            .I(UART_TRANSMITTER_state_7_N_1749_2_cascade_));
    InMux I__9774 (
            .O(N__42011),
            .I(N__42008));
    LocalMux I__9773 (
            .O(N__42008),
            .I(n18032));
    InMux I__9772 (
            .O(N__42005),
            .I(N__42000));
    InMux I__9771 (
            .O(N__42004),
            .I(N__41995));
    InMux I__9770 (
            .O(N__42003),
            .I(N__41995));
    LocalMux I__9769 (
            .O(N__42000),
            .I(n8488));
    LocalMux I__9768 (
            .O(N__41995),
            .I(n8488));
    InMux I__9767 (
            .O(N__41990),
            .I(N__41985));
    InMux I__9766 (
            .O(N__41989),
            .I(N__41980));
    InMux I__9765 (
            .O(N__41988),
            .I(N__41980));
    LocalMux I__9764 (
            .O(N__41985),
            .I(n17709));
    LocalMux I__9763 (
            .O(N__41980),
            .I(n17709));
    CascadeMux I__9762 (
            .O(N__41975),
            .I(N__41971));
    CascadeMux I__9761 (
            .O(N__41974),
            .I(N__41968));
    InMux I__9760 (
            .O(N__41971),
            .I(N__41965));
    InMux I__9759 (
            .O(N__41968),
            .I(N__41961));
    LocalMux I__9758 (
            .O(N__41965),
            .I(N__41957));
    InMux I__9757 (
            .O(N__41964),
            .I(N__41954));
    LocalMux I__9756 (
            .O(N__41961),
            .I(N__41951));
    InMux I__9755 (
            .O(N__41960),
            .I(N__41948));
    Span4Mux_h I__9754 (
            .O(N__41957),
            .I(N__41945));
    LocalMux I__9753 (
            .O(N__41954),
            .I(\c0.delay_counter_6 ));
    Odrv12 I__9752 (
            .O(N__41951),
            .I(\c0.delay_counter_6 ));
    LocalMux I__9751 (
            .O(N__41948),
            .I(\c0.delay_counter_6 ));
    Odrv4 I__9750 (
            .O(N__41945),
            .I(\c0.delay_counter_6 ));
    CascadeMux I__9749 (
            .O(N__41936),
            .I(N__41932));
    InMux I__9748 (
            .O(N__41935),
            .I(N__41928));
    InMux I__9747 (
            .O(N__41932),
            .I(N__41924));
    InMux I__9746 (
            .O(N__41931),
            .I(N__41921));
    LocalMux I__9745 (
            .O(N__41928),
            .I(N__41918));
    InMux I__9744 (
            .O(N__41927),
            .I(N__41915));
    LocalMux I__9743 (
            .O(N__41924),
            .I(N__41910));
    LocalMux I__9742 (
            .O(N__41921),
            .I(N__41910));
    Span4Mux_h I__9741 (
            .O(N__41918),
            .I(N__41907));
    LocalMux I__9740 (
            .O(N__41915),
            .I(\c0.delay_counter_9 ));
    Odrv4 I__9739 (
            .O(N__41910),
            .I(\c0.delay_counter_9 ));
    Odrv4 I__9738 (
            .O(N__41907),
            .I(\c0.delay_counter_9 ));
    InMux I__9737 (
            .O(N__41900),
            .I(N__41897));
    LocalMux I__9736 (
            .O(N__41897),
            .I(N__41894));
    Span4Mux_h I__9735 (
            .O(N__41894),
            .I(N__41891));
    Odrv4 I__9734 (
            .O(N__41891),
            .I(\c0.n17753 ));
    CascadeMux I__9733 (
            .O(N__41888),
            .I(\c0.n17662_cascade_ ));
    InMux I__9732 (
            .O(N__41885),
            .I(N__41882));
    LocalMux I__9731 (
            .O(N__41882),
            .I(N__41878));
    CascadeMux I__9730 (
            .O(N__41881),
            .I(N__41875));
    Span4Mux_h I__9729 (
            .O(N__41878),
            .I(N__41872));
    InMux I__9728 (
            .O(N__41875),
            .I(N__41869));
    Odrv4 I__9727 (
            .O(N__41872),
            .I(rand_setpoint_23));
    LocalMux I__9726 (
            .O(N__41869),
            .I(rand_setpoint_23));
    CascadeMux I__9725 (
            .O(N__41864),
            .I(\c0.n2041_cascade_ ));
    InMux I__9724 (
            .O(N__41861),
            .I(N__41858));
    LocalMux I__9723 (
            .O(N__41858),
            .I(N__41855));
    Span4Mux_s2_v I__9722 (
            .O(N__41855),
            .I(N__41852));
    Odrv4 I__9721 (
            .O(N__41852),
            .I(\c0.n17974 ));
    InMux I__9720 (
            .O(N__41849),
            .I(N__41846));
    LocalMux I__9719 (
            .O(N__41846),
            .I(N__41842));
    CascadeMux I__9718 (
            .O(N__41845),
            .I(N__41839));
    Span4Mux_s1_v I__9717 (
            .O(N__41842),
            .I(N__41836));
    InMux I__9716 (
            .O(N__41839),
            .I(N__41833));
    Odrv4 I__9715 (
            .O(N__41836),
            .I(rand_setpoint_16));
    LocalMux I__9714 (
            .O(N__41833),
            .I(rand_setpoint_16));
    CascadeMux I__9713 (
            .O(N__41828),
            .I(\c0.n17693_cascade_ ));
    InMux I__9712 (
            .O(N__41825),
            .I(N__41822));
    LocalMux I__9711 (
            .O(N__41822),
            .I(N__41818));
    InMux I__9710 (
            .O(N__41821),
            .I(N__41815));
    Span4Mux_h I__9709 (
            .O(N__41818),
            .I(N__41810));
    LocalMux I__9708 (
            .O(N__41815),
            .I(N__41810));
    Odrv4 I__9707 (
            .O(N__41810),
            .I(\c0.data_out_6_0 ));
    InMux I__9706 (
            .O(N__41807),
            .I(N__41804));
    LocalMux I__9705 (
            .O(N__41804),
            .I(N__41801));
    Span4Mux_v I__9704 (
            .O(N__41801),
            .I(N__41798));
    Span4Mux_h I__9703 (
            .O(N__41798),
            .I(N__41794));
    InMux I__9702 (
            .O(N__41797),
            .I(N__41789));
    Span4Mux_h I__9701 (
            .O(N__41794),
            .I(N__41786));
    CascadeMux I__9700 (
            .O(N__41793),
            .I(N__41783));
    InMux I__9699 (
            .O(N__41792),
            .I(N__41780));
    LocalMux I__9698 (
            .O(N__41789),
            .I(N__41775));
    Sp12to4 I__9697 (
            .O(N__41786),
            .I(N__41775));
    InMux I__9696 (
            .O(N__41783),
            .I(N__41772));
    LocalMux I__9695 (
            .O(N__41780),
            .I(N__41769));
    Span12Mux_v I__9694 (
            .O(N__41775),
            .I(N__41766));
    LocalMux I__9693 (
            .O(N__41772),
            .I(data_out_1_7));
    Odrv4 I__9692 (
            .O(N__41769),
            .I(data_out_1_7));
    Odrv12 I__9691 (
            .O(N__41766),
            .I(data_out_1_7));
    InMux I__9690 (
            .O(N__41759),
            .I(N__41756));
    LocalMux I__9689 (
            .O(N__41756),
            .I(N__41752));
    InMux I__9688 (
            .O(N__41755),
            .I(N__41749));
    Odrv12 I__9687 (
            .O(N__41752),
            .I(\c0.n17578 ));
    LocalMux I__9686 (
            .O(N__41749),
            .I(\c0.n17578 ));
    InMux I__9685 (
            .O(N__41744),
            .I(N__41740));
    InMux I__9684 (
            .O(N__41743),
            .I(N__41735));
    LocalMux I__9683 (
            .O(N__41740),
            .I(N__41732));
    InMux I__9682 (
            .O(N__41739),
            .I(N__41727));
    InMux I__9681 (
            .O(N__41738),
            .I(N__41727));
    LocalMux I__9680 (
            .O(N__41735),
            .I(N__41722));
    Span4Mux_h I__9679 (
            .O(N__41732),
            .I(N__41722));
    LocalMux I__9678 (
            .O(N__41727),
            .I(\c0.delay_counter_10 ));
    Odrv4 I__9677 (
            .O(N__41722),
            .I(\c0.delay_counter_10 ));
    InMux I__9676 (
            .O(N__41717),
            .I(N__41713));
    CascadeMux I__9675 (
            .O(N__41716),
            .I(N__41710));
    LocalMux I__9674 (
            .O(N__41713),
            .I(N__41707));
    InMux I__9673 (
            .O(N__41710),
            .I(N__41704));
    Odrv12 I__9672 (
            .O(N__41707),
            .I(rand_setpoint_12));
    LocalMux I__9671 (
            .O(N__41704),
            .I(rand_setpoint_12));
    CascadeMux I__9670 (
            .O(N__41699),
            .I(\c0.n17931_cascade_ ));
    CascadeMux I__9669 (
            .O(N__41696),
            .I(N__41693));
    InMux I__9668 (
            .O(N__41693),
            .I(N__41690));
    LocalMux I__9667 (
            .O(N__41690),
            .I(N__41686));
    InMux I__9666 (
            .O(N__41689),
            .I(N__41683));
    Span4Mux_h I__9665 (
            .O(N__41686),
            .I(N__41678));
    LocalMux I__9664 (
            .O(N__41683),
            .I(N__41678));
    Span4Mux_s2_v I__9663 (
            .O(N__41678),
            .I(N__41675));
    Odrv4 I__9662 (
            .O(N__41675),
            .I(\c0.n17400 ));
    InMux I__9661 (
            .O(N__41672),
            .I(N__41669));
    LocalMux I__9660 (
            .O(N__41669),
            .I(N__41665));
    InMux I__9659 (
            .O(N__41668),
            .I(N__41662));
    Odrv12 I__9658 (
            .O(N__41665),
            .I(\c0.data_out_7__4__N_550 ));
    LocalMux I__9657 (
            .O(N__41662),
            .I(\c0.data_out_7__4__N_550 ));
    InMux I__9656 (
            .O(N__41657),
            .I(N__41653));
    InMux I__9655 (
            .O(N__41656),
            .I(N__41650));
    LocalMux I__9654 (
            .O(N__41653),
            .I(N__41645));
    LocalMux I__9653 (
            .O(N__41650),
            .I(N__41642));
    InMux I__9652 (
            .O(N__41649),
            .I(N__41637));
    InMux I__9651 (
            .O(N__41648),
            .I(N__41637));
    Span4Mux_h I__9650 (
            .O(N__41645),
            .I(N__41634));
    Span4Mux_h I__9649 (
            .O(N__41642),
            .I(N__41631));
    LocalMux I__9648 (
            .O(N__41637),
            .I(\c0.data_out_7_4 ));
    Odrv4 I__9647 (
            .O(N__41634),
            .I(\c0.data_out_7_4 ));
    Odrv4 I__9646 (
            .O(N__41631),
            .I(\c0.data_out_7_4 ));
    InMux I__9645 (
            .O(N__41624),
            .I(N__41616));
    InMux I__9644 (
            .O(N__41623),
            .I(N__41616));
    InMux I__9643 (
            .O(N__41622),
            .I(N__41611));
    InMux I__9642 (
            .O(N__41621),
            .I(N__41608));
    LocalMux I__9641 (
            .O(N__41616),
            .I(N__41605));
    InMux I__9640 (
            .O(N__41615),
            .I(N__41600));
    InMux I__9639 (
            .O(N__41614),
            .I(N__41600));
    LocalMux I__9638 (
            .O(N__41611),
            .I(data_out_5__4__N_959));
    LocalMux I__9637 (
            .O(N__41608),
            .I(data_out_5__4__N_959));
    Odrv4 I__9636 (
            .O(N__41605),
            .I(data_out_5__4__N_959));
    LocalMux I__9635 (
            .O(N__41600),
            .I(data_out_5__4__N_959));
    InMux I__9634 (
            .O(N__41591),
            .I(N__41588));
    LocalMux I__9633 (
            .O(N__41588),
            .I(N__41584));
    CascadeMux I__9632 (
            .O(N__41587),
            .I(N__41581));
    Span4Mux_h I__9631 (
            .O(N__41584),
            .I(N__41578));
    InMux I__9630 (
            .O(N__41581),
            .I(N__41575));
    Odrv4 I__9629 (
            .O(N__41578),
            .I(rand_setpoint_28));
    LocalMux I__9628 (
            .O(N__41575),
            .I(rand_setpoint_28));
    CascadeMux I__9627 (
            .O(N__41570),
            .I(\c0.n17967_cascade_ ));
    CascadeMux I__9626 (
            .O(N__41567),
            .I(N__41564));
    InMux I__9625 (
            .O(N__41564),
            .I(N__41561));
    LocalMux I__9624 (
            .O(N__41561),
            .I(N__41558));
    Odrv4 I__9623 (
            .O(N__41558),
            .I(\c0.n6_adj_2467 ));
    InMux I__9622 (
            .O(N__41555),
            .I(N__41552));
    LocalMux I__9621 (
            .O(N__41552),
            .I(N__41549));
    Odrv4 I__9620 (
            .O(N__41549),
            .I(\c0.n9276 ));
    CascadeMux I__9619 (
            .O(N__41546),
            .I(N__41542));
    InMux I__9618 (
            .O(N__41545),
            .I(N__41538));
    InMux I__9617 (
            .O(N__41542),
            .I(N__41535));
    InMux I__9616 (
            .O(N__41541),
            .I(N__41532));
    LocalMux I__9615 (
            .O(N__41538),
            .I(\c0.n8634 ));
    LocalMux I__9614 (
            .O(N__41535),
            .I(\c0.n8634 ));
    LocalMux I__9613 (
            .O(N__41532),
            .I(\c0.n8634 ));
    CascadeMux I__9612 (
            .O(N__41525),
            .I(\c0.n9276_cascade_ ));
    InMux I__9611 (
            .O(N__41522),
            .I(N__41519));
    LocalMux I__9610 (
            .O(N__41519),
            .I(N__41516));
    Span4Mux_v I__9609 (
            .O(N__41516),
            .I(N__41513));
    Odrv4 I__9608 (
            .O(N__41513),
            .I(\c0.data_out_7__1__N_626 ));
    CascadeMux I__9607 (
            .O(N__41510),
            .I(\c0.n17623_cascade_ ));
    InMux I__9606 (
            .O(N__41507),
            .I(N__41504));
    LocalMux I__9605 (
            .O(N__41504),
            .I(N__41501));
    Span4Mux_v I__9604 (
            .O(N__41501),
            .I(N__41497));
    CascadeMux I__9603 (
            .O(N__41500),
            .I(N__41494));
    Span4Mux_h I__9602 (
            .O(N__41497),
            .I(N__41491));
    InMux I__9601 (
            .O(N__41494),
            .I(N__41488));
    Odrv4 I__9600 (
            .O(N__41491),
            .I(rand_setpoint_8));
    LocalMux I__9599 (
            .O(N__41488),
            .I(rand_setpoint_8));
    CascadeMux I__9598 (
            .O(N__41483),
            .I(\c0.n17916_cascade_ ));
    InMux I__9597 (
            .O(N__41480),
            .I(N__41477));
    LocalMux I__9596 (
            .O(N__41477),
            .I(N__41473));
    InMux I__9595 (
            .O(N__41476),
            .I(N__41470));
    Span4Mux_h I__9594 (
            .O(N__41473),
            .I(N__41467));
    LocalMux I__9593 (
            .O(N__41470),
            .I(N__41464));
    Span4Mux_v I__9592 (
            .O(N__41467),
            .I(N__41461));
    Span4Mux_h I__9591 (
            .O(N__41464),
            .I(N__41458));
    Odrv4 I__9590 (
            .O(N__41461),
            .I(\c0.data_out_7_0 ));
    Odrv4 I__9589 (
            .O(N__41458),
            .I(\c0.data_out_7_0 ));
    CascadeMux I__9588 (
            .O(N__41453),
            .I(N__41450));
    InMux I__9587 (
            .O(N__41450),
            .I(N__41447));
    LocalMux I__9586 (
            .O(N__41447),
            .I(N__41444));
    Span4Mux_v I__9585 (
            .O(N__41444),
            .I(N__41441));
    Span4Mux_v I__9584 (
            .O(N__41441),
            .I(N__41438));
    Odrv4 I__9583 (
            .O(N__41438),
            .I(\c0.n8486 ));
    CascadeMux I__9582 (
            .O(N__41435),
            .I(\c0.n8486_cascade_ ));
    InMux I__9581 (
            .O(N__41432),
            .I(N__41429));
    LocalMux I__9580 (
            .O(N__41429),
            .I(N__41426));
    Odrv12 I__9579 (
            .O(N__41426),
            .I(\c0.n16450 ));
    InMux I__9578 (
            .O(N__41423),
            .I(N__41420));
    LocalMux I__9577 (
            .O(N__41420),
            .I(N__41417));
    Span4Mux_v I__9576 (
            .O(N__41417),
            .I(N__41414));
    Odrv4 I__9575 (
            .O(N__41414),
            .I(n4_adj_2612));
    InMux I__9574 (
            .O(N__41411),
            .I(N__41407));
    CascadeMux I__9573 (
            .O(N__41410),
            .I(N__41404));
    LocalMux I__9572 (
            .O(N__41407),
            .I(N__41401));
    InMux I__9571 (
            .O(N__41404),
            .I(N__41398));
    Odrv12 I__9570 (
            .O(N__41401),
            .I(rand_setpoint_13));
    LocalMux I__9569 (
            .O(N__41398),
            .I(rand_setpoint_13));
    CascadeMux I__9568 (
            .O(N__41393),
            .I(\c0.n17925_cascade_ ));
    InMux I__9567 (
            .O(N__41390),
            .I(N__41387));
    LocalMux I__9566 (
            .O(N__41387),
            .I(\c0.n18068 ));
    InMux I__9565 (
            .O(N__41384),
            .I(N__41381));
    LocalMux I__9564 (
            .O(N__41381),
            .I(\c0.n5_adj_2490 ));
    InMux I__9563 (
            .O(N__41378),
            .I(N__41375));
    LocalMux I__9562 (
            .O(N__41375),
            .I(\c0.data_out_10_4 ));
    InMux I__9561 (
            .O(N__41372),
            .I(N__41369));
    LocalMux I__9560 (
            .O(N__41369),
            .I(\c0.n18067 ));
    InMux I__9559 (
            .O(N__41366),
            .I(N__41363));
    LocalMux I__9558 (
            .O(N__41363),
            .I(\c0.n18092 ));
    InMux I__9557 (
            .O(N__41360),
            .I(N__41357));
    LocalMux I__9556 (
            .O(N__41357),
            .I(N__41354));
    Odrv4 I__9555 (
            .O(N__41354),
            .I(\c0.n18094 ));
    InMux I__9554 (
            .O(N__41351),
            .I(N__41348));
    LocalMux I__9553 (
            .O(N__41348),
            .I(N__41345));
    Span4Mux_h I__9552 (
            .O(N__41345),
            .I(N__41342));
    Span4Mux_v I__9551 (
            .O(N__41342),
            .I(N__41339));
    Odrv4 I__9550 (
            .O(N__41339),
            .I(\c0.n18096 ));
    InMux I__9549 (
            .O(N__41336),
            .I(N__41333));
    LocalMux I__9548 (
            .O(N__41333),
            .I(N__41330));
    Span4Mux_h I__9547 (
            .O(N__41330),
            .I(N__41327));
    Odrv4 I__9546 (
            .O(N__41327),
            .I(\c0.n18088 ));
    InMux I__9545 (
            .O(N__41324),
            .I(N__41321));
    LocalMux I__9544 (
            .O(N__41321),
            .I(N__41317));
    InMux I__9543 (
            .O(N__41320),
            .I(N__41314));
    Span4Mux_h I__9542 (
            .O(N__41317),
            .I(N__41311));
    LocalMux I__9541 (
            .O(N__41314),
            .I(byte_transmit_counter_5));
    Odrv4 I__9540 (
            .O(N__41311),
            .I(byte_transmit_counter_5));
    InMux I__9539 (
            .O(N__41306),
            .I(N__41303));
    LocalMux I__9538 (
            .O(N__41303),
            .I(N__41300));
    Span4Mux_h I__9537 (
            .O(N__41300),
            .I(N__41296));
    InMux I__9536 (
            .O(N__41299),
            .I(N__41293));
    Odrv4 I__9535 (
            .O(N__41296),
            .I(tx_transmit_N_2239_5));
    LocalMux I__9534 (
            .O(N__41293),
            .I(tx_transmit_N_2239_5));
    InMux I__9533 (
            .O(N__41288),
            .I(\c0.n16354 ));
    InMux I__9532 (
            .O(N__41285),
            .I(\c0.n16355 ));
    InMux I__9531 (
            .O(N__41282),
            .I(N__41278));
    InMux I__9530 (
            .O(N__41281),
            .I(N__41275));
    LocalMux I__9529 (
            .O(N__41278),
            .I(byte_transmit_counter_7));
    LocalMux I__9528 (
            .O(N__41275),
            .I(byte_transmit_counter_7));
    InMux I__9527 (
            .O(N__41270),
            .I(\c0.n16356 ));
    InMux I__9526 (
            .O(N__41267),
            .I(N__41263));
    InMux I__9525 (
            .O(N__41266),
            .I(N__41260));
    LocalMux I__9524 (
            .O(N__41263),
            .I(tx_transmit_N_2239_7));
    LocalMux I__9523 (
            .O(N__41260),
            .I(tx_transmit_N_2239_7));
    InMux I__9522 (
            .O(N__41255),
            .I(N__41251));
    CascadeMux I__9521 (
            .O(N__41254),
            .I(N__41248));
    LocalMux I__9520 (
            .O(N__41251),
            .I(N__41245));
    InMux I__9519 (
            .O(N__41248),
            .I(N__41241));
    Span4Mux_h I__9518 (
            .O(N__41245),
            .I(N__41238));
    InMux I__9517 (
            .O(N__41244),
            .I(N__41234));
    LocalMux I__9516 (
            .O(N__41241),
            .I(N__41231));
    Span4Mux_v I__9515 (
            .O(N__41238),
            .I(N__41228));
    InMux I__9514 (
            .O(N__41237),
            .I(N__41225));
    LocalMux I__9513 (
            .O(N__41234),
            .I(data_out_3_4));
    Odrv4 I__9512 (
            .O(N__41231),
            .I(data_out_3_4));
    Odrv4 I__9511 (
            .O(N__41228),
            .I(data_out_3_4));
    LocalMux I__9510 (
            .O(N__41225),
            .I(data_out_3_4));
    CascadeMux I__9509 (
            .O(N__41216),
            .I(\c0.n18093_cascade_ ));
    CascadeMux I__9508 (
            .O(N__41213),
            .I(\c0.n18399_cascade_ ));
    CascadeMux I__9507 (
            .O(N__41210),
            .I(N__41206));
    InMux I__9506 (
            .O(N__41209),
            .I(N__41203));
    InMux I__9505 (
            .O(N__41206),
            .I(N__41200));
    LocalMux I__9504 (
            .O(N__41203),
            .I(tx_transmit_N_2239_4));
    LocalMux I__9503 (
            .O(N__41200),
            .I(tx_transmit_N_2239_4));
    InMux I__9502 (
            .O(N__41195),
            .I(N__41192));
    LocalMux I__9501 (
            .O(N__41192),
            .I(\c0.n5_adj_2447 ));
    CascadeMux I__9500 (
            .O(N__41189),
            .I(\c0.n17941_cascade_ ));
    InMux I__9499 (
            .O(N__41186),
            .I(N__41183));
    LocalMux I__9498 (
            .O(N__41183),
            .I(\c0.n18396 ));
    CascadeMux I__9497 (
            .O(N__41180),
            .I(n8529_cascade_));
    CascadeMux I__9496 (
            .O(N__41177),
            .I(\c0.n8550_cascade_ ));
    InMux I__9495 (
            .O(N__41174),
            .I(N__41171));
    LocalMux I__9494 (
            .O(N__41171),
            .I(n121_adj_2606));
    InMux I__9493 (
            .O(N__41168),
            .I(N__41165));
    LocalMux I__9492 (
            .O(N__41165),
            .I(n8529));
    CascadeMux I__9491 (
            .O(N__41162),
            .I(n121_adj_2606_cascade_));
    InMux I__9490 (
            .O(N__41159),
            .I(N__41156));
    LocalMux I__9489 (
            .O(N__41156),
            .I(N__41153));
    Odrv4 I__9488 (
            .O(N__41153),
            .I(n13_adj_2652));
    InMux I__9487 (
            .O(N__41150),
            .I(N__41147));
    LocalMux I__9486 (
            .O(N__41147),
            .I(\c0.n251 ));
    InMux I__9485 (
            .O(N__41144),
            .I(\c0.n16350 ));
    InMux I__9484 (
            .O(N__41141),
            .I(\c0.n16351 ));
    InMux I__9483 (
            .O(N__41138),
            .I(\c0.n16352 ));
    InMux I__9482 (
            .O(N__41135),
            .I(\c0.n16353 ));
    InMux I__9481 (
            .O(N__41132),
            .I(N__41129));
    LocalMux I__9480 (
            .O(N__41129),
            .I(N__41126));
    Odrv4 I__9479 (
            .O(N__41126),
            .I(\c0.n18008 ));
    InMux I__9478 (
            .O(N__41123),
            .I(N__41118));
    InMux I__9477 (
            .O(N__41122),
            .I(N__41115));
    InMux I__9476 (
            .O(N__41121),
            .I(N__41112));
    LocalMux I__9475 (
            .O(N__41118),
            .I(N__41107));
    LocalMux I__9474 (
            .O(N__41115),
            .I(N__41107));
    LocalMux I__9473 (
            .O(N__41112),
            .I(\c0.delay_counter_3 ));
    Odrv4 I__9472 (
            .O(N__41107),
            .I(\c0.delay_counter_3 ));
    InMux I__9471 (
            .O(N__41102),
            .I(N__41097));
    InMux I__9470 (
            .O(N__41101),
            .I(N__41092));
    InMux I__9469 (
            .O(N__41100),
            .I(N__41092));
    LocalMux I__9468 (
            .O(N__41097),
            .I(\c0.delay_counter_1 ));
    LocalMux I__9467 (
            .O(N__41092),
            .I(\c0.delay_counter_1 ));
    CascadeMux I__9466 (
            .O(N__41087),
            .I(N__41082));
    InMux I__9465 (
            .O(N__41086),
            .I(N__41079));
    InMux I__9464 (
            .O(N__41085),
            .I(N__41076));
    InMux I__9463 (
            .O(N__41082),
            .I(N__41073));
    LocalMux I__9462 (
            .O(N__41079),
            .I(\c0.delay_counter_2 ));
    LocalMux I__9461 (
            .O(N__41076),
            .I(\c0.delay_counter_2 ));
    LocalMux I__9460 (
            .O(N__41073),
            .I(\c0.delay_counter_2 ));
    InMux I__9459 (
            .O(N__41066),
            .I(N__41061));
    InMux I__9458 (
            .O(N__41065),
            .I(N__41058));
    InMux I__9457 (
            .O(N__41064),
            .I(N__41055));
    LocalMux I__9456 (
            .O(N__41061),
            .I(\c0.delay_counter_4 ));
    LocalMux I__9455 (
            .O(N__41058),
            .I(\c0.delay_counter_4 ));
    LocalMux I__9454 (
            .O(N__41055),
            .I(\c0.delay_counter_4 ));
    InMux I__9453 (
            .O(N__41048),
            .I(N__41044));
    InMux I__9452 (
            .O(N__41047),
            .I(N__41040));
    LocalMux I__9451 (
            .O(N__41044),
            .I(N__41037));
    InMux I__9450 (
            .O(N__41043),
            .I(N__41033));
    LocalMux I__9449 (
            .O(N__41040),
            .I(N__41028));
    Span4Mux_v I__9448 (
            .O(N__41037),
            .I(N__41028));
    InMux I__9447 (
            .O(N__41036),
            .I(N__41025));
    LocalMux I__9446 (
            .O(N__41033),
            .I(delay_counter_0));
    Odrv4 I__9445 (
            .O(N__41028),
            .I(delay_counter_0));
    LocalMux I__9444 (
            .O(N__41025),
            .I(delay_counter_0));
    InMux I__9443 (
            .O(N__41018),
            .I(N__41015));
    LocalMux I__9442 (
            .O(N__41015),
            .I(N__41012));
    Span4Mux_v I__9441 (
            .O(N__41012),
            .I(N__41006));
    CascadeMux I__9440 (
            .O(N__41011),
            .I(N__41003));
    CascadeMux I__9439 (
            .O(N__41010),
            .I(N__41000));
    InMux I__9438 (
            .O(N__41009),
            .I(N__40997));
    Sp12to4 I__9437 (
            .O(N__41006),
            .I(N__40994));
    InMux I__9436 (
            .O(N__41003),
            .I(N__40989));
    InMux I__9435 (
            .O(N__41000),
            .I(N__40989));
    LocalMux I__9434 (
            .O(N__40997),
            .I(delay_counter_13));
    Odrv12 I__9433 (
            .O(N__40994),
            .I(delay_counter_13));
    LocalMux I__9432 (
            .O(N__40989),
            .I(delay_counter_13));
    InMux I__9431 (
            .O(N__40982),
            .I(N__40978));
    InMux I__9430 (
            .O(N__40981),
            .I(N__40975));
    LocalMux I__9429 (
            .O(N__40978),
            .I(N__40969));
    LocalMux I__9428 (
            .O(N__40975),
            .I(N__40969));
    InMux I__9427 (
            .O(N__40974),
            .I(N__40965));
    Span4Mux_v I__9426 (
            .O(N__40969),
            .I(N__40962));
    InMux I__9425 (
            .O(N__40968),
            .I(N__40959));
    LocalMux I__9424 (
            .O(N__40965),
            .I(delay_counter_14));
    Odrv4 I__9423 (
            .O(N__40962),
            .I(delay_counter_14));
    LocalMux I__9422 (
            .O(N__40959),
            .I(delay_counter_14));
    InMux I__9421 (
            .O(N__40952),
            .I(N__40949));
    LocalMux I__9420 (
            .O(N__40949),
            .I(\c0.n7264 ));
    CascadeMux I__9419 (
            .O(N__40946),
            .I(n29_cascade_));
    InMux I__9418 (
            .O(N__40943),
            .I(N__40939));
    InMux I__9417 (
            .O(N__40942),
            .I(N__40936));
    LocalMux I__9416 (
            .O(N__40939),
            .I(data_in_12_6));
    LocalMux I__9415 (
            .O(N__40936),
            .I(data_in_12_6));
    CascadeMux I__9414 (
            .O(N__40931),
            .I(\c0.n149_cascade_ ));
    InMux I__9413 (
            .O(N__40928),
            .I(N__40925));
    LocalMux I__9412 (
            .O(N__40925),
            .I(N__40922));
    Span4Mux_h I__9411 (
            .O(N__40922),
            .I(N__40919));
    Odrv4 I__9410 (
            .O(N__40919),
            .I(\c0.n93 ));
    CascadeMux I__9409 (
            .O(N__40916),
            .I(N__40913));
    InMux I__9408 (
            .O(N__40913),
            .I(N__40910));
    LocalMux I__9407 (
            .O(N__40910),
            .I(n17958));
    InMux I__9406 (
            .O(N__40907),
            .I(N__40904));
    LocalMux I__9405 (
            .O(N__40904),
            .I(n43));
    CascadeMux I__9404 (
            .O(N__40901),
            .I(N__40898));
    InMux I__9403 (
            .O(N__40898),
            .I(N__40895));
    LocalMux I__9402 (
            .O(N__40895),
            .I(\c0.n7271 ));
    CascadeMux I__9401 (
            .O(N__40892),
            .I(N__40889));
    InMux I__9400 (
            .O(N__40889),
            .I(N__40886));
    LocalMux I__9399 (
            .O(N__40886),
            .I(N__40883));
    Odrv4 I__9398 (
            .O(N__40883),
            .I(\c0.n18105 ));
    InMux I__9397 (
            .O(N__40880),
            .I(N__40877));
    LocalMux I__9396 (
            .O(N__40877),
            .I(\c0.n18012 ));
    InMux I__9395 (
            .O(N__40874),
            .I(N__40871));
    LocalMux I__9394 (
            .O(N__40871),
            .I(N__40868));
    Odrv4 I__9393 (
            .O(N__40868),
            .I(\c0.n17936 ));
    InMux I__9392 (
            .O(N__40865),
            .I(N__40862));
    LocalMux I__9391 (
            .O(N__40862),
            .I(\c0.n7275 ));
    CascadeMux I__9390 (
            .O(N__40859),
            .I(N__40856));
    InMux I__9389 (
            .O(N__40856),
            .I(N__40853));
    LocalMux I__9388 (
            .O(N__40853),
            .I(\c0.n7274 ));
    InMux I__9387 (
            .O(N__40850),
            .I(N__40843));
    InMux I__9386 (
            .O(N__40849),
            .I(N__40838));
    InMux I__9385 (
            .O(N__40848),
            .I(N__40838));
    InMux I__9384 (
            .O(N__40847),
            .I(N__40835));
    CascadeMux I__9383 (
            .O(N__40846),
            .I(N__40832));
    LocalMux I__9382 (
            .O(N__40843),
            .I(N__40824));
    LocalMux I__9381 (
            .O(N__40838),
            .I(N__40824));
    LocalMux I__9380 (
            .O(N__40835),
            .I(N__40824));
    InMux I__9379 (
            .O(N__40832),
            .I(N__40819));
    InMux I__9378 (
            .O(N__40831),
            .I(N__40819));
    Odrv12 I__9377 (
            .O(N__40824),
            .I(data_out_6__7__N_678));
    LocalMux I__9376 (
            .O(N__40819),
            .I(data_out_6__7__N_678));
    CascadeMux I__9375 (
            .O(N__40814),
            .I(n96_cascade_));
    CascadeMux I__9374 (
            .O(N__40811),
            .I(n47_cascade_));
    InMux I__9373 (
            .O(N__40808),
            .I(N__40804));
    InMux I__9372 (
            .O(N__40807),
            .I(N__40801));
    LocalMux I__9371 (
            .O(N__40804),
            .I(n2615));
    LocalMux I__9370 (
            .O(N__40801),
            .I(n2615));
    CascadeMux I__9369 (
            .O(N__40796),
            .I(n41_cascade_));
    InMux I__9368 (
            .O(N__40793),
            .I(N__40789));
    InMux I__9367 (
            .O(N__40792),
            .I(N__40786));
    LocalMux I__9366 (
            .O(N__40789),
            .I(N__40783));
    LocalMux I__9365 (
            .O(N__40786),
            .I(N__40780));
    Span4Mux_h I__9364 (
            .O(N__40783),
            .I(N__40777));
    Odrv4 I__9363 (
            .O(N__40780),
            .I(\c0.data_out_5__3__N_964 ));
    Odrv4 I__9362 (
            .O(N__40777),
            .I(\c0.data_out_5__3__N_964 ));
    CascadeMux I__9361 (
            .O(N__40772),
            .I(\c0.data_out_5__3__N_964_cascade_ ));
    CascadeMux I__9360 (
            .O(N__40769),
            .I(\c0.data_out_6__3__N_785_cascade_ ));
    InMux I__9359 (
            .O(N__40766),
            .I(N__40762));
    CascadeMux I__9358 (
            .O(N__40765),
            .I(N__40759));
    LocalMux I__9357 (
            .O(N__40762),
            .I(N__40756));
    InMux I__9356 (
            .O(N__40759),
            .I(N__40753));
    Odrv4 I__9355 (
            .O(N__40756),
            .I(rand_setpoint_19));
    LocalMux I__9354 (
            .O(N__40753),
            .I(rand_setpoint_19));
    CascadeMux I__9353 (
            .O(N__40748),
            .I(\c0.n2181_cascade_ ));
    InMux I__9352 (
            .O(N__40745),
            .I(N__40733));
    InMux I__9351 (
            .O(N__40744),
            .I(N__40733));
    InMux I__9350 (
            .O(N__40743),
            .I(N__40733));
    InMux I__9349 (
            .O(N__40742),
            .I(N__40730));
    InMux I__9348 (
            .O(N__40741),
            .I(N__40725));
    InMux I__9347 (
            .O(N__40740),
            .I(N__40722));
    LocalMux I__9346 (
            .O(N__40733),
            .I(N__40717));
    LocalMux I__9345 (
            .O(N__40730),
            .I(N__40717));
    InMux I__9344 (
            .O(N__40729),
            .I(N__40712));
    InMux I__9343 (
            .O(N__40728),
            .I(N__40712));
    LocalMux I__9342 (
            .O(N__40725),
            .I(data_out_6__6__N_729));
    LocalMux I__9341 (
            .O(N__40722),
            .I(data_out_6__6__N_729));
    Odrv12 I__9340 (
            .O(N__40717),
            .I(data_out_6__6__N_729));
    LocalMux I__9339 (
            .O(N__40712),
            .I(data_out_6__6__N_729));
    CascadeMux I__9338 (
            .O(N__40703),
            .I(N__40698));
    InMux I__9337 (
            .O(N__40702),
            .I(N__40694));
    InMux I__9336 (
            .O(N__40701),
            .I(N__40690));
    InMux I__9335 (
            .O(N__40698),
            .I(N__40687));
    CascadeMux I__9334 (
            .O(N__40697),
            .I(N__40683));
    LocalMux I__9333 (
            .O(N__40694),
            .I(N__40680));
    InMux I__9332 (
            .O(N__40693),
            .I(N__40677));
    LocalMux I__9331 (
            .O(N__40690),
            .I(N__40674));
    LocalMux I__9330 (
            .O(N__40687),
            .I(N__40671));
    InMux I__9329 (
            .O(N__40686),
            .I(N__40666));
    InMux I__9328 (
            .O(N__40683),
            .I(N__40666));
    Odrv4 I__9327 (
            .O(N__40680),
            .I(data_out_2_0));
    LocalMux I__9326 (
            .O(N__40677),
            .I(data_out_2_0));
    Odrv4 I__9325 (
            .O(N__40674),
            .I(data_out_2_0));
    Odrv12 I__9324 (
            .O(N__40671),
            .I(data_out_2_0));
    LocalMux I__9323 (
            .O(N__40666),
            .I(data_out_2_0));
    InMux I__9322 (
            .O(N__40655),
            .I(N__40652));
    LocalMux I__9321 (
            .O(N__40652),
            .I(N__40649));
    Span4Mux_v I__9320 (
            .O(N__40649),
            .I(N__40646));
    Odrv4 I__9319 (
            .O(N__40646),
            .I(\c0.n2_adj_2483 ));
    InMux I__9318 (
            .O(N__40643),
            .I(N__40640));
    LocalMux I__9317 (
            .O(N__40640),
            .I(\c0.n17389 ));
    CascadeMux I__9316 (
            .O(N__40637),
            .I(\c0.n17389_cascade_ ));
    CascadeMux I__9315 (
            .O(N__40634),
            .I(\c0.n17600_cascade_ ));
    InMux I__9314 (
            .O(N__40631),
            .I(N__40628));
    LocalMux I__9313 (
            .O(N__40628),
            .I(N__40625));
    Span4Mux_h I__9312 (
            .O(N__40625),
            .I(N__40622));
    Odrv4 I__9311 (
            .O(N__40622),
            .I(\c0.n9658 ));
    CascadeMux I__9310 (
            .O(N__40619),
            .I(\c0.n17398_cascade_ ));
    InMux I__9309 (
            .O(N__40616),
            .I(N__40612));
    CascadeMux I__9308 (
            .O(N__40615),
            .I(N__40609));
    LocalMux I__9307 (
            .O(N__40612),
            .I(N__40606));
    InMux I__9306 (
            .O(N__40609),
            .I(N__40603));
    Odrv4 I__9305 (
            .O(N__40606),
            .I(rand_setpoint_20));
    LocalMux I__9304 (
            .O(N__40603),
            .I(rand_setpoint_20));
    CascadeMux I__9303 (
            .O(N__40598),
            .I(\c0.n2146_cascade_ ));
    CascadeMux I__9302 (
            .O(N__40595),
            .I(\c0.data_out_6__7__N_675_cascade_ ));
    InMux I__9301 (
            .O(N__40592),
            .I(N__40589));
    LocalMux I__9300 (
            .O(N__40589),
            .I(N__40585));
    CascadeMux I__9299 (
            .O(N__40588),
            .I(N__40582));
    Span4Mux_h I__9298 (
            .O(N__40585),
            .I(N__40579));
    InMux I__9297 (
            .O(N__40582),
            .I(N__40576));
    Odrv4 I__9296 (
            .O(N__40579),
            .I(rand_setpoint_15));
    LocalMux I__9295 (
            .O(N__40576),
            .I(rand_setpoint_15));
    CascadeMux I__9294 (
            .O(N__40571),
            .I(\c0.n17928_cascade_ ));
    InMux I__9293 (
            .O(N__40568),
            .I(N__40565));
    LocalMux I__9292 (
            .O(N__40565),
            .I(N__40562));
    Span4Mux_h I__9291 (
            .O(N__40562),
            .I(N__40558));
    InMux I__9290 (
            .O(N__40561),
            .I(N__40555));
    Odrv4 I__9289 (
            .O(N__40558),
            .I(rand_setpoint_14));
    LocalMux I__9288 (
            .O(N__40555),
            .I(rand_setpoint_14));
    InMux I__9287 (
            .O(N__40550),
            .I(N__40547));
    LocalMux I__9286 (
            .O(N__40547),
            .I(N__40544));
    Odrv4 I__9285 (
            .O(N__40544),
            .I(\c0.n17465 ));
    CascadeMux I__9284 (
            .O(N__40541),
            .I(\c0.n17906_cascade_ ));
    InMux I__9283 (
            .O(N__40538),
            .I(N__40535));
    LocalMux I__9282 (
            .O(N__40535),
            .I(N__40532));
    Span4Mux_h I__9281 (
            .O(N__40532),
            .I(N__40529));
    Odrv4 I__9280 (
            .O(N__40529),
            .I(\c0.n17921 ));
    InMux I__9279 (
            .O(N__40526),
            .I(N__40523));
    LocalMux I__9278 (
            .O(N__40523),
            .I(N__40520));
    Odrv4 I__9277 (
            .O(N__40520),
            .I(\c0.data_out_10_6 ));
    CascadeMux I__9276 (
            .O(N__40517),
            .I(\c0.n18393_cascade_ ));
    InMux I__9275 (
            .O(N__40514),
            .I(N__40511));
    LocalMux I__9274 (
            .O(N__40511),
            .I(tx_data_3_N_keep));
    InMux I__9273 (
            .O(N__40508),
            .I(N__40505));
    LocalMux I__9272 (
            .O(N__40505),
            .I(\c0.n18095 ));
    CascadeMux I__9271 (
            .O(N__40502),
            .I(N__40498));
    InMux I__9270 (
            .O(N__40501),
            .I(N__40493));
    InMux I__9269 (
            .O(N__40498),
            .I(N__40490));
    InMux I__9268 (
            .O(N__40497),
            .I(N__40485));
    InMux I__9267 (
            .O(N__40496),
            .I(N__40485));
    LocalMux I__9266 (
            .O(N__40493),
            .I(N__40482));
    LocalMux I__9265 (
            .O(N__40490),
            .I(N__40477));
    LocalMux I__9264 (
            .O(N__40485),
            .I(N__40477));
    Odrv4 I__9263 (
            .O(N__40482),
            .I(n9646));
    Odrv4 I__9262 (
            .O(N__40477),
            .I(n9646));
    InMux I__9261 (
            .O(N__40472),
            .I(N__40468));
    InMux I__9260 (
            .O(N__40471),
            .I(N__40465));
    LocalMux I__9259 (
            .O(N__40468),
            .I(n9920));
    LocalMux I__9258 (
            .O(N__40465),
            .I(n9920));
    CascadeMux I__9257 (
            .O(N__40460),
            .I(N__40456));
    CascadeMux I__9256 (
            .O(N__40459),
            .I(N__40453));
    InMux I__9255 (
            .O(N__40456),
            .I(N__40446));
    InMux I__9254 (
            .O(N__40453),
            .I(N__40446));
    InMux I__9253 (
            .O(N__40452),
            .I(N__40441));
    InMux I__9252 (
            .O(N__40451),
            .I(N__40438));
    LocalMux I__9251 (
            .O(N__40446),
            .I(N__40435));
    InMux I__9250 (
            .O(N__40445),
            .I(N__40430));
    InMux I__9249 (
            .O(N__40444),
            .I(N__40430));
    LocalMux I__9248 (
            .O(N__40441),
            .I(N__40427));
    LocalMux I__9247 (
            .O(N__40438),
            .I(N__40418));
    Span4Mux_h I__9246 (
            .O(N__40435),
            .I(N__40418));
    LocalMux I__9245 (
            .O(N__40430),
            .I(N__40418));
    Span4Mux_v I__9244 (
            .O(N__40427),
            .I(N__40418));
    Odrv4 I__9243 (
            .O(N__40418),
            .I(r_Bit_Index_0_adj_2627));
    InMux I__9242 (
            .O(N__40415),
            .I(N__40408));
    InMux I__9241 (
            .O(N__40414),
            .I(N__40408));
    InMux I__9240 (
            .O(N__40413),
            .I(N__40405));
    LocalMux I__9239 (
            .O(N__40408),
            .I(N__40397));
    LocalMux I__9238 (
            .O(N__40405),
            .I(N__40397));
    InMux I__9237 (
            .O(N__40404),
            .I(N__40394));
    InMux I__9236 (
            .O(N__40403),
            .I(N__40389));
    InMux I__9235 (
            .O(N__40402),
            .I(N__40389));
    Span4Mux_h I__9234 (
            .O(N__40397),
            .I(N__40386));
    LocalMux I__9233 (
            .O(N__40394),
            .I(r_SM_Main_2_N_2323_1));
    LocalMux I__9232 (
            .O(N__40389),
            .I(r_SM_Main_2_N_2323_1));
    Odrv4 I__9231 (
            .O(N__40386),
            .I(r_SM_Main_2_N_2323_1));
    CascadeMux I__9230 (
            .O(N__40379),
            .I(n4_adj_2653_cascade_));
    CascadeMux I__9229 (
            .O(N__40376),
            .I(N__40366));
    InMux I__9228 (
            .O(N__40375),
            .I(N__40363));
    InMux I__9227 (
            .O(N__40374),
            .I(N__40354));
    InMux I__9226 (
            .O(N__40373),
            .I(N__40354));
    InMux I__9225 (
            .O(N__40372),
            .I(N__40354));
    InMux I__9224 (
            .O(N__40371),
            .I(N__40354));
    CascadeMux I__9223 (
            .O(N__40370),
            .I(N__40351));
    CascadeMux I__9222 (
            .O(N__40369),
            .I(N__40347));
    InMux I__9221 (
            .O(N__40366),
            .I(N__40343));
    LocalMux I__9220 (
            .O(N__40363),
            .I(N__40340));
    LocalMux I__9219 (
            .O(N__40354),
            .I(N__40334));
    InMux I__9218 (
            .O(N__40351),
            .I(N__40329));
    InMux I__9217 (
            .O(N__40350),
            .I(N__40329));
    InMux I__9216 (
            .O(N__40347),
            .I(N__40326));
    InMux I__9215 (
            .O(N__40346),
            .I(N__40321));
    LocalMux I__9214 (
            .O(N__40343),
            .I(N__40316));
    Span4Mux_h I__9213 (
            .O(N__40340),
            .I(N__40316));
    InMux I__9212 (
            .O(N__40339),
            .I(N__40313));
    InMux I__9211 (
            .O(N__40338),
            .I(N__40308));
    InMux I__9210 (
            .O(N__40337),
            .I(N__40308));
    Span4Mux_h I__9209 (
            .O(N__40334),
            .I(N__40305));
    LocalMux I__9208 (
            .O(N__40329),
            .I(N__40302));
    LocalMux I__9207 (
            .O(N__40326),
            .I(N__40299));
    InMux I__9206 (
            .O(N__40325),
            .I(N__40294));
    InMux I__9205 (
            .O(N__40324),
            .I(N__40294));
    LocalMux I__9204 (
            .O(N__40321),
            .I(N__40281));
    Span4Mux_v I__9203 (
            .O(N__40316),
            .I(N__40281));
    LocalMux I__9202 (
            .O(N__40313),
            .I(N__40281));
    LocalMux I__9201 (
            .O(N__40308),
            .I(N__40278));
    Span4Mux_h I__9200 (
            .O(N__40305),
            .I(N__40273));
    Span4Mux_h I__9199 (
            .O(N__40302),
            .I(N__40273));
    Span4Mux_v I__9198 (
            .O(N__40299),
            .I(N__40268));
    LocalMux I__9197 (
            .O(N__40294),
            .I(N__40268));
    InMux I__9196 (
            .O(N__40293),
            .I(N__40259));
    InMux I__9195 (
            .O(N__40292),
            .I(N__40259));
    InMux I__9194 (
            .O(N__40291),
            .I(N__40259));
    InMux I__9193 (
            .O(N__40290),
            .I(N__40259));
    InMux I__9192 (
            .O(N__40289),
            .I(N__40254));
    InMux I__9191 (
            .O(N__40288),
            .I(N__40254));
    Odrv4 I__9190 (
            .O(N__40281),
            .I(r_SM_Main_2));
    Odrv12 I__9189 (
            .O(N__40278),
            .I(r_SM_Main_2));
    Odrv4 I__9188 (
            .O(N__40273),
            .I(r_SM_Main_2));
    Odrv4 I__9187 (
            .O(N__40268),
            .I(r_SM_Main_2));
    LocalMux I__9186 (
            .O(N__40259),
            .I(r_SM_Main_2));
    LocalMux I__9185 (
            .O(N__40254),
            .I(r_SM_Main_2));
    CascadeMux I__9184 (
            .O(N__40241),
            .I(N__40234));
    CascadeMux I__9183 (
            .O(N__40240),
            .I(N__40231));
    InMux I__9182 (
            .O(N__40239),
            .I(N__40226));
    InMux I__9181 (
            .O(N__40238),
            .I(N__40226));
    CascadeMux I__9180 (
            .O(N__40237),
            .I(N__40223));
    InMux I__9179 (
            .O(N__40234),
            .I(N__40216));
    InMux I__9178 (
            .O(N__40231),
            .I(N__40216));
    LocalMux I__9177 (
            .O(N__40226),
            .I(N__40210));
    InMux I__9176 (
            .O(N__40223),
            .I(N__40207));
    CascadeMux I__9175 (
            .O(N__40222),
            .I(N__40203));
    InMux I__9174 (
            .O(N__40221),
            .I(N__40200));
    LocalMux I__9173 (
            .O(N__40216),
            .I(N__40197));
    InMux I__9172 (
            .O(N__40215),
            .I(N__40194));
    InMux I__9171 (
            .O(N__40214),
            .I(N__40191));
    InMux I__9170 (
            .O(N__40213),
            .I(N__40188));
    Span4Mux_h I__9169 (
            .O(N__40210),
            .I(N__40183));
    LocalMux I__9168 (
            .O(N__40207),
            .I(N__40183));
    InMux I__9167 (
            .O(N__40206),
            .I(N__40178));
    InMux I__9166 (
            .O(N__40203),
            .I(N__40178));
    LocalMux I__9165 (
            .O(N__40200),
            .I(r_SM_Main_0));
    Odrv12 I__9164 (
            .O(N__40197),
            .I(r_SM_Main_0));
    LocalMux I__9163 (
            .O(N__40194),
            .I(r_SM_Main_0));
    LocalMux I__9162 (
            .O(N__40191),
            .I(r_SM_Main_0));
    LocalMux I__9161 (
            .O(N__40188),
            .I(r_SM_Main_0));
    Odrv4 I__9160 (
            .O(N__40183),
            .I(r_SM_Main_0));
    LocalMux I__9159 (
            .O(N__40178),
            .I(r_SM_Main_0));
    CascadeMux I__9158 (
            .O(N__40163),
            .I(N__40156));
    CascadeMux I__9157 (
            .O(N__40162),
            .I(N__40150));
    CascadeMux I__9156 (
            .O(N__40161),
            .I(N__40147));
    InMux I__9155 (
            .O(N__40160),
            .I(N__40142));
    InMux I__9154 (
            .O(N__40159),
            .I(N__40137));
    InMux I__9153 (
            .O(N__40156),
            .I(N__40137));
    InMux I__9152 (
            .O(N__40155),
            .I(N__40134));
    InMux I__9151 (
            .O(N__40154),
            .I(N__40130));
    InMux I__9150 (
            .O(N__40153),
            .I(N__40123));
    InMux I__9149 (
            .O(N__40150),
            .I(N__40123));
    InMux I__9148 (
            .O(N__40147),
            .I(N__40123));
    InMux I__9147 (
            .O(N__40146),
            .I(N__40120));
    InMux I__9146 (
            .O(N__40145),
            .I(N__40117));
    LocalMux I__9145 (
            .O(N__40142),
            .I(N__40112));
    LocalMux I__9144 (
            .O(N__40137),
            .I(N__40112));
    LocalMux I__9143 (
            .O(N__40134),
            .I(N__40109));
    CascadeMux I__9142 (
            .O(N__40133),
            .I(N__40104));
    LocalMux I__9141 (
            .O(N__40130),
            .I(N__40096));
    LocalMux I__9140 (
            .O(N__40123),
            .I(N__40096));
    LocalMux I__9139 (
            .O(N__40120),
            .I(N__40091));
    LocalMux I__9138 (
            .O(N__40117),
            .I(N__40091));
    Span4Mux_v I__9137 (
            .O(N__40112),
            .I(N__40086));
    Span4Mux_h I__9136 (
            .O(N__40109),
            .I(N__40086));
    InMux I__9135 (
            .O(N__40108),
            .I(N__40077));
    InMux I__9134 (
            .O(N__40107),
            .I(N__40077));
    InMux I__9133 (
            .O(N__40104),
            .I(N__40077));
    InMux I__9132 (
            .O(N__40103),
            .I(N__40077));
    InMux I__9131 (
            .O(N__40102),
            .I(N__40072));
    InMux I__9130 (
            .O(N__40101),
            .I(N__40072));
    Odrv4 I__9129 (
            .O(N__40096),
            .I(r_SM_Main_1));
    Odrv4 I__9128 (
            .O(N__40091),
            .I(r_SM_Main_1));
    Odrv4 I__9127 (
            .O(N__40086),
            .I(r_SM_Main_1));
    LocalMux I__9126 (
            .O(N__40077),
            .I(r_SM_Main_1));
    LocalMux I__9125 (
            .O(N__40072),
            .I(r_SM_Main_1));
    InMux I__9124 (
            .O(N__40061),
            .I(N__40058));
    LocalMux I__9123 (
            .O(N__40058),
            .I(\c0.tx_active_prev ));
    InMux I__9122 (
            .O(N__40055),
            .I(N__40051));
    InMux I__9121 (
            .O(N__40054),
            .I(N__40048));
    LocalMux I__9120 (
            .O(N__40051),
            .I(\c0.n17349 ));
    LocalMux I__9119 (
            .O(N__40048),
            .I(\c0.n17349 ));
    InMux I__9118 (
            .O(N__40043),
            .I(N__40040));
    LocalMux I__9117 (
            .O(N__40040),
            .I(\c0.n17937 ));
    CascadeMux I__9116 (
            .O(N__40037),
            .I(\c0.n18390_cascade_ ));
    InMux I__9115 (
            .O(N__40034),
            .I(\c0.n16311 ));
    InMux I__9114 (
            .O(N__40031),
            .I(N__40028));
    LocalMux I__9113 (
            .O(N__40028),
            .I(N__40025));
    Odrv4 I__9112 (
            .O(N__40025),
            .I(\c0.n18011 ));
    InMux I__9111 (
            .O(N__40022),
            .I(bfn_12_25_0_));
    InMux I__9110 (
            .O(N__40019),
            .I(N__40016));
    LocalMux I__9109 (
            .O(N__40016),
            .I(\c0.n7266 ));
    InMux I__9108 (
            .O(N__40013),
            .I(\c0.n16313 ));
    CascadeMux I__9107 (
            .O(N__40010),
            .I(N__40007));
    InMux I__9106 (
            .O(N__40007),
            .I(N__40004));
    LocalMux I__9105 (
            .O(N__40004),
            .I(N__40001));
    Odrv4 I__9104 (
            .O(N__40001),
            .I(\c0.n7265 ));
    InMux I__9103 (
            .O(N__39998),
            .I(\c0.n16314 ));
    InMux I__9102 (
            .O(N__39995),
            .I(\c0.n16315 ));
    InMux I__9101 (
            .O(N__39992),
            .I(\c0.n16316 ));
    InMux I__9100 (
            .O(N__39989),
            .I(\c0.n16317 ));
    InMux I__9099 (
            .O(N__39986),
            .I(\c0.n16318 ));
    InMux I__9098 (
            .O(N__39983),
            .I(N__39980));
    LocalMux I__9097 (
            .O(N__39980),
            .I(\c0.n25_adj_2517 ));
    CascadeMux I__9096 (
            .O(N__39977),
            .I(\c0.n1314_cascade_ ));
    InMux I__9095 (
            .O(N__39974),
            .I(bfn_12_24_0_));
    InMux I__9094 (
            .O(N__39971),
            .I(\c0.n16305 ));
    InMux I__9093 (
            .O(N__39968),
            .I(N__39965));
    LocalMux I__9092 (
            .O(N__39965),
            .I(\c0.n7273 ));
    InMux I__9091 (
            .O(N__39962),
            .I(\c0.n16306 ));
    CascadeMux I__9090 (
            .O(N__39959),
            .I(N__39956));
    InMux I__9089 (
            .O(N__39956),
            .I(N__39953));
    LocalMux I__9088 (
            .O(N__39953),
            .I(\c0.n7272 ));
    InMux I__9087 (
            .O(N__39950),
            .I(\c0.n16307 ));
    InMux I__9086 (
            .O(N__39947),
            .I(\c0.n16308 ));
    InMux I__9085 (
            .O(N__39944),
            .I(\c0.n16309 ));
    InMux I__9084 (
            .O(N__39941),
            .I(N__39938));
    LocalMux I__9083 (
            .O(N__39938),
            .I(\c0.n7269 ));
    InMux I__9082 (
            .O(N__39935),
            .I(\c0.n16310 ));
    InMux I__9081 (
            .O(N__39932),
            .I(N__39928));
    InMux I__9080 (
            .O(N__39931),
            .I(N__39925));
    LocalMux I__9079 (
            .O(N__39928),
            .I(N__39922));
    LocalMux I__9078 (
            .O(N__39925),
            .I(N__39919));
    Span4Mux_h I__9077 (
            .O(N__39922),
            .I(N__39915));
    Span4Mux_h I__9076 (
            .O(N__39919),
            .I(N__39912));
    InMux I__9075 (
            .O(N__39918),
            .I(N__39909));
    Span4Mux_h I__9074 (
            .O(N__39915),
            .I(N__39906));
    Odrv4 I__9073 (
            .O(N__39912),
            .I(\c0.data_in_6_1 ));
    LocalMux I__9072 (
            .O(N__39909),
            .I(\c0.data_in_6_1 ));
    Odrv4 I__9071 (
            .O(N__39906),
            .I(\c0.data_in_6_1 ));
    CascadeMux I__9070 (
            .O(N__39899),
            .I(N__39896));
    InMux I__9069 (
            .O(N__39896),
            .I(N__39893));
    LocalMux I__9068 (
            .O(N__39893),
            .I(N__39889));
    CascadeMux I__9067 (
            .O(N__39892),
            .I(N__39886));
    Span4Mux_v I__9066 (
            .O(N__39889),
            .I(N__39882));
    InMux I__9065 (
            .O(N__39886),
            .I(N__39879));
    InMux I__9064 (
            .O(N__39885),
            .I(N__39875));
    Span4Mux_s1_h I__9063 (
            .O(N__39882),
            .I(N__39872));
    LocalMux I__9062 (
            .O(N__39879),
            .I(N__39869));
    InMux I__9061 (
            .O(N__39878),
            .I(N__39866));
    LocalMux I__9060 (
            .O(N__39875),
            .I(N__39863));
    Span4Mux_h I__9059 (
            .O(N__39872),
            .I(N__39858));
    Span4Mux_v I__9058 (
            .O(N__39869),
            .I(N__39858));
    LocalMux I__9057 (
            .O(N__39866),
            .I(N__39853));
    Span4Mux_v I__9056 (
            .O(N__39863),
            .I(N__39853));
    Span4Mux_h I__9055 (
            .O(N__39858),
            .I(N__39850));
    Odrv4 I__9054 (
            .O(N__39853),
            .I(data_in_5_1));
    Odrv4 I__9053 (
            .O(N__39850),
            .I(data_in_5_1));
    InMux I__9052 (
            .O(N__39845),
            .I(N__39841));
    InMux I__9051 (
            .O(N__39844),
            .I(N__39838));
    LocalMux I__9050 (
            .O(N__39841),
            .I(N__39835));
    LocalMux I__9049 (
            .O(N__39838),
            .I(N__39831));
    Span4Mux_h I__9048 (
            .O(N__39835),
            .I(N__39828));
    InMux I__9047 (
            .O(N__39834),
            .I(N__39825));
    Span4Mux_h I__9046 (
            .O(N__39831),
            .I(N__39822));
    Span4Mux_h I__9045 (
            .O(N__39828),
            .I(N__39819));
    LocalMux I__9044 (
            .O(N__39825),
            .I(data_in_10_6));
    Odrv4 I__9043 (
            .O(N__39822),
            .I(data_in_10_6));
    Odrv4 I__9042 (
            .O(N__39819),
            .I(data_in_10_6));
    InMux I__9041 (
            .O(N__39812),
            .I(N__39808));
    InMux I__9040 (
            .O(N__39811),
            .I(N__39805));
    LocalMux I__9039 (
            .O(N__39808),
            .I(data_in_11_6));
    LocalMux I__9038 (
            .O(N__39805),
            .I(data_in_11_6));
    InMux I__9037 (
            .O(N__39800),
            .I(N__39797));
    LocalMux I__9036 (
            .O(N__39797),
            .I(N__39794));
    Odrv4 I__9035 (
            .O(N__39794),
            .I(\c0.n17755 ));
    CascadeMux I__9034 (
            .O(N__39791),
            .I(\c0.n17525_cascade_ ));
    InMux I__9033 (
            .O(N__39788),
            .I(N__39785));
    LocalMux I__9032 (
            .O(N__39785),
            .I(N__39782));
    Odrv4 I__9031 (
            .O(N__39782),
            .I(\c0.rx.n9553 ));
    InMux I__9030 (
            .O(N__39779),
            .I(N__39775));
    InMux I__9029 (
            .O(N__39778),
            .I(N__39768));
    LocalMux I__9028 (
            .O(N__39775),
            .I(N__39765));
    InMux I__9027 (
            .O(N__39774),
            .I(N__39758));
    InMux I__9026 (
            .O(N__39773),
            .I(N__39758));
    InMux I__9025 (
            .O(N__39772),
            .I(N__39758));
    CascadeMux I__9024 (
            .O(N__39771),
            .I(N__39755));
    LocalMux I__9023 (
            .O(N__39768),
            .I(N__39749));
    Span4Mux_s2_v I__9022 (
            .O(N__39765),
            .I(N__39744));
    LocalMux I__9021 (
            .O(N__39758),
            .I(N__39744));
    InMux I__9020 (
            .O(N__39755),
            .I(N__39735));
    InMux I__9019 (
            .O(N__39754),
            .I(N__39735));
    InMux I__9018 (
            .O(N__39753),
            .I(N__39735));
    InMux I__9017 (
            .O(N__39752),
            .I(N__39735));
    Span4Mux_v I__9016 (
            .O(N__39749),
            .I(N__39732));
    Span4Mux_h I__9015 (
            .O(N__39744),
            .I(N__39729));
    LocalMux I__9014 (
            .O(N__39735),
            .I(N__39726));
    Odrv4 I__9013 (
            .O(N__39732),
            .I(\c0.rx.r_SM_Main_2 ));
    Odrv4 I__9012 (
            .O(N__39729),
            .I(\c0.rx.r_SM_Main_2 ));
    Odrv4 I__9011 (
            .O(N__39726),
            .I(\c0.rx.r_SM_Main_2 ));
    CascadeMux I__9010 (
            .O(N__39719),
            .I(N__39714));
    InMux I__9009 (
            .O(N__39718),
            .I(N__39707));
    InMux I__9008 (
            .O(N__39717),
            .I(N__39704));
    InMux I__9007 (
            .O(N__39714),
            .I(N__39697));
    InMux I__9006 (
            .O(N__39713),
            .I(N__39697));
    InMux I__9005 (
            .O(N__39712),
            .I(N__39697));
    InMux I__9004 (
            .O(N__39711),
            .I(N__39694));
    InMux I__9003 (
            .O(N__39710),
            .I(N__39691));
    LocalMux I__9002 (
            .O(N__39707),
            .I(N__39684));
    LocalMux I__9001 (
            .O(N__39704),
            .I(N__39675));
    LocalMux I__9000 (
            .O(N__39697),
            .I(N__39675));
    LocalMux I__8999 (
            .O(N__39694),
            .I(N__39675));
    LocalMux I__8998 (
            .O(N__39691),
            .I(N__39675));
    InMux I__8997 (
            .O(N__39690),
            .I(N__39666));
    InMux I__8996 (
            .O(N__39689),
            .I(N__39666));
    InMux I__8995 (
            .O(N__39688),
            .I(N__39666));
    InMux I__8994 (
            .O(N__39687),
            .I(N__39666));
    Span4Mux_v I__8993 (
            .O(N__39684),
            .I(N__39661));
    Span4Mux_s3_v I__8992 (
            .O(N__39675),
            .I(N__39661));
    LocalMux I__8991 (
            .O(N__39666),
            .I(\c0.rx.r_SM_Main_1 ));
    Odrv4 I__8990 (
            .O(N__39661),
            .I(\c0.rx.r_SM_Main_1 ));
    InMux I__8989 (
            .O(N__39656),
            .I(N__39651));
    InMux I__8988 (
            .O(N__39655),
            .I(N__39645));
    InMux I__8987 (
            .O(N__39654),
            .I(N__39645));
    LocalMux I__8986 (
            .O(N__39651),
            .I(N__39642));
    CascadeMux I__8985 (
            .O(N__39650),
            .I(N__39638));
    LocalMux I__8984 (
            .O(N__39645),
            .I(N__39635));
    Span4Mux_s2_v I__8983 (
            .O(N__39642),
            .I(N__39632));
    InMux I__8982 (
            .O(N__39641),
            .I(N__39626));
    InMux I__8981 (
            .O(N__39638),
            .I(N__39626));
    Span4Mux_h I__8980 (
            .O(N__39635),
            .I(N__39623));
    Sp12to4 I__8979 (
            .O(N__39632),
            .I(N__39620));
    InMux I__8978 (
            .O(N__39631),
            .I(N__39617));
    LocalMux I__8977 (
            .O(N__39626),
            .I(\c0.rx.r_SM_Main_2_N_2380_2 ));
    Odrv4 I__8976 (
            .O(N__39623),
            .I(\c0.rx.r_SM_Main_2_N_2380_2 ));
    Odrv12 I__8975 (
            .O(N__39620),
            .I(\c0.rx.r_SM_Main_2_N_2380_2 ));
    LocalMux I__8974 (
            .O(N__39617),
            .I(\c0.rx.r_SM_Main_2_N_2380_2 ));
    SRMux I__8973 (
            .O(N__39608),
            .I(N__39605));
    LocalMux I__8972 (
            .O(N__39605),
            .I(N__39602));
    Span4Mux_s2_v I__8971 (
            .O(N__39602),
            .I(N__39599));
    Span4Mux_h I__8970 (
            .O(N__39599),
            .I(N__39596));
    Span4Mux_s2_v I__8969 (
            .O(N__39596),
            .I(N__39593));
    Odrv4 I__8968 (
            .O(N__39593),
            .I(\c0.rx.n17351 ));
    InMux I__8967 (
            .O(N__39590),
            .I(N__39581));
    InMux I__8966 (
            .O(N__39589),
            .I(N__39572));
    InMux I__8965 (
            .O(N__39588),
            .I(N__39572));
    InMux I__8964 (
            .O(N__39587),
            .I(N__39572));
    InMux I__8963 (
            .O(N__39586),
            .I(N__39572));
    InMux I__8962 (
            .O(N__39585),
            .I(N__39566));
    InMux I__8961 (
            .O(N__39584),
            .I(N__39566));
    LocalMux I__8960 (
            .O(N__39581),
            .I(N__39560));
    LocalMux I__8959 (
            .O(N__39572),
            .I(N__39560));
    InMux I__8958 (
            .O(N__39571),
            .I(N__39557));
    LocalMux I__8957 (
            .O(N__39566),
            .I(N__39553));
    InMux I__8956 (
            .O(N__39565),
            .I(N__39550));
    Span4Mux_h I__8955 (
            .O(N__39560),
            .I(N__39547));
    LocalMux I__8954 (
            .O(N__39557),
            .I(N__39544));
    InMux I__8953 (
            .O(N__39556),
            .I(N__39541));
    Span4Mux_h I__8952 (
            .O(N__39553),
            .I(N__39536));
    LocalMux I__8951 (
            .O(N__39550),
            .I(N__39536));
    Span4Mux_h I__8950 (
            .O(N__39547),
            .I(N__39533));
    Span12Mux_v I__8949 (
            .O(N__39544),
            .I(N__39528));
    LocalMux I__8948 (
            .O(N__39541),
            .I(N__39528));
    Odrv4 I__8947 (
            .O(N__39536),
            .I(\c0.rx.r_SM_Main_0 ));
    Odrv4 I__8946 (
            .O(N__39533),
            .I(\c0.rx.r_SM_Main_0 ));
    Odrv12 I__8945 (
            .O(N__39528),
            .I(\c0.rx.r_SM_Main_0 ));
    InMux I__8944 (
            .O(N__39521),
            .I(N__39518));
    LocalMux I__8943 (
            .O(N__39518),
            .I(N__39515));
    Span4Mux_h I__8942 (
            .O(N__39515),
            .I(N__39512));
    Odrv4 I__8941 (
            .O(N__39512),
            .I(\c0.rx.n17376 ));
    CascadeMux I__8940 (
            .O(N__39509),
            .I(\c0.data_out_6__2__N_803_cascade_ ));
    InMux I__8939 (
            .O(N__39506),
            .I(N__39502));
    CascadeMux I__8938 (
            .O(N__39505),
            .I(N__39499));
    LocalMux I__8937 (
            .O(N__39502),
            .I(N__39496));
    InMux I__8936 (
            .O(N__39499),
            .I(N__39493));
    Odrv4 I__8935 (
            .O(N__39496),
            .I(rand_setpoint_18));
    LocalMux I__8934 (
            .O(N__39493),
            .I(rand_setpoint_18));
    CascadeMux I__8933 (
            .O(N__39488),
            .I(\c0.n2216_cascade_ ));
    InMux I__8932 (
            .O(N__39485),
            .I(N__39481));
    InMux I__8931 (
            .O(N__39484),
            .I(N__39478));
    LocalMux I__8930 (
            .O(N__39481),
            .I(N__39475));
    LocalMux I__8929 (
            .O(N__39478),
            .I(N__39470));
    Span4Mux_v I__8928 (
            .O(N__39475),
            .I(N__39470));
    Odrv4 I__8927 (
            .O(N__39470),
            .I(\c0.data_out_6_2 ));
    InMux I__8926 (
            .O(N__39467),
            .I(N__39464));
    LocalMux I__8925 (
            .O(N__39464),
            .I(N__39460));
    CascadeMux I__8924 (
            .O(N__39463),
            .I(N__39457));
    Span4Mux_h I__8923 (
            .O(N__39460),
            .I(N__39454));
    InMux I__8922 (
            .O(N__39457),
            .I(N__39451));
    Odrv4 I__8921 (
            .O(N__39454),
            .I(rand_setpoint_26));
    LocalMux I__8920 (
            .O(N__39451),
            .I(rand_setpoint_26));
    InMux I__8919 (
            .O(N__39446),
            .I(N__39443));
    LocalMux I__8918 (
            .O(N__39443),
            .I(\c0.data_out_6__2__N_803 ));
    CascadeMux I__8917 (
            .O(N__39440),
            .I(\c0.n17964_cascade_ ));
    InMux I__8916 (
            .O(N__39437),
            .I(N__39433));
    CascadeMux I__8915 (
            .O(N__39436),
            .I(N__39430));
    LocalMux I__8914 (
            .O(N__39433),
            .I(N__39427));
    InMux I__8913 (
            .O(N__39430),
            .I(N__39424));
    Odrv4 I__8912 (
            .O(N__39427),
            .I(rand_setpoint_0));
    LocalMux I__8911 (
            .O(N__39424),
            .I(rand_setpoint_0));
    CascadeMux I__8910 (
            .O(N__39419),
            .I(\c0.n8953_cascade_ ));
    InMux I__8909 (
            .O(N__39416),
            .I(N__39413));
    LocalMux I__8908 (
            .O(N__39413),
            .I(N__39409));
    CascadeMux I__8907 (
            .O(N__39412),
            .I(N__39406));
    Span4Mux_h I__8906 (
            .O(N__39409),
            .I(N__39403));
    InMux I__8905 (
            .O(N__39406),
            .I(N__39400));
    Odrv4 I__8904 (
            .O(N__39403),
            .I(rand_setpoint_5));
    LocalMux I__8903 (
            .O(N__39400),
            .I(rand_setpoint_5));
    InMux I__8902 (
            .O(N__39395),
            .I(N__39392));
    LocalMux I__8901 (
            .O(N__39392),
            .I(N__39389));
    Sp12to4 I__8900 (
            .O(N__39389),
            .I(N__39386));
    Odrv12 I__8899 (
            .O(N__39386),
            .I(\c0.n5 ));
    InMux I__8898 (
            .O(N__39383),
            .I(N__39380));
    LocalMux I__8897 (
            .O(N__39380),
            .I(\c0.n17972 ));
    InMux I__8896 (
            .O(N__39377),
            .I(N__39374));
    LocalMux I__8895 (
            .O(N__39374),
            .I(\c0.n18501 ));
    CascadeMux I__8894 (
            .O(N__39371),
            .I(tx_data_0_N_keep_cascade_));
    InMux I__8893 (
            .O(N__39368),
            .I(N__39364));
    InMux I__8892 (
            .O(N__39367),
            .I(N__39361));
    LocalMux I__8891 (
            .O(N__39364),
            .I(N__39358));
    LocalMux I__8890 (
            .O(N__39361),
            .I(r_Tx_Data_0));
    Odrv12 I__8889 (
            .O(N__39358),
            .I(r_Tx_Data_0));
    InMux I__8888 (
            .O(N__39353),
            .I(N__39350));
    LocalMux I__8887 (
            .O(N__39350),
            .I(N__39346));
    InMux I__8886 (
            .O(N__39349),
            .I(N__39343));
    Span4Mux_v I__8885 (
            .O(N__39346),
            .I(N__39340));
    LocalMux I__8884 (
            .O(N__39343),
            .I(data_in_15_5));
    Odrv4 I__8883 (
            .O(N__39340),
            .I(data_in_15_5));
    InMux I__8882 (
            .O(N__39335),
            .I(N__39332));
    LocalMux I__8881 (
            .O(N__39332),
            .I(N__39328));
    InMux I__8880 (
            .O(N__39331),
            .I(N__39325));
    Odrv12 I__8879 (
            .O(N__39328),
            .I(data_in_14_5));
    LocalMux I__8878 (
            .O(N__39325),
            .I(data_in_14_5));
    InMux I__8877 (
            .O(N__39320),
            .I(N__39317));
    LocalMux I__8876 (
            .O(N__39317),
            .I(n4958));
    InMux I__8875 (
            .O(N__39314),
            .I(N__39308));
    InMux I__8874 (
            .O(N__39313),
            .I(N__39308));
    LocalMux I__8873 (
            .O(N__39308),
            .I(N__39304));
    InMux I__8872 (
            .O(N__39307),
            .I(N__39301));
    Span4Mux_h I__8871 (
            .O(N__39304),
            .I(N__39297));
    LocalMux I__8870 (
            .O(N__39301),
            .I(N__39294));
    InMux I__8869 (
            .O(N__39300),
            .I(N__39291));
    Span4Mux_h I__8868 (
            .O(N__39297),
            .I(N__39287));
    Span4Mux_v I__8867 (
            .O(N__39294),
            .I(N__39282));
    LocalMux I__8866 (
            .O(N__39291),
            .I(N__39279));
    InMux I__8865 (
            .O(N__39290),
            .I(N__39276));
    Sp12to4 I__8864 (
            .O(N__39287),
            .I(N__39273));
    InMux I__8863 (
            .O(N__39286),
            .I(N__39270));
    InMux I__8862 (
            .O(N__39285),
            .I(N__39267));
    Span4Mux_h I__8861 (
            .O(N__39282),
            .I(N__39262));
    Span4Mux_v I__8860 (
            .O(N__39279),
            .I(N__39262));
    LocalMux I__8859 (
            .O(N__39276),
            .I(r_Bit_Index_2_adj_2625));
    Odrv12 I__8858 (
            .O(N__39273),
            .I(r_Bit_Index_2_adj_2625));
    LocalMux I__8857 (
            .O(N__39270),
            .I(r_Bit_Index_2_adj_2625));
    LocalMux I__8856 (
            .O(N__39267),
            .I(r_Bit_Index_2_adj_2625));
    Odrv4 I__8855 (
            .O(N__39262),
            .I(r_Bit_Index_2_adj_2625));
    CascadeMux I__8854 (
            .O(N__39251),
            .I(n4958_cascade_));
    CascadeMux I__8853 (
            .O(N__39248),
            .I(n9920_cascade_));
    InMux I__8852 (
            .O(N__39245),
            .I(N__39242));
    LocalMux I__8851 (
            .O(N__39242),
            .I(N__39237));
    InMux I__8850 (
            .O(N__39241),
            .I(N__39231));
    InMux I__8849 (
            .O(N__39240),
            .I(N__39231));
    Span4Mux_h I__8848 (
            .O(N__39237),
            .I(N__39225));
    InMux I__8847 (
            .O(N__39236),
            .I(N__39222));
    LocalMux I__8846 (
            .O(N__39231),
            .I(N__39219));
    InMux I__8845 (
            .O(N__39230),
            .I(N__39216));
    InMux I__8844 (
            .O(N__39229),
            .I(N__39211));
    InMux I__8843 (
            .O(N__39228),
            .I(N__39211));
    Span4Mux_h I__8842 (
            .O(N__39225),
            .I(N__39206));
    LocalMux I__8841 (
            .O(N__39222),
            .I(N__39206));
    Span12Mux_v I__8840 (
            .O(N__39219),
            .I(N__39203));
    LocalMux I__8839 (
            .O(N__39216),
            .I(r_Bit_Index_1_adj_2626));
    LocalMux I__8838 (
            .O(N__39211),
            .I(r_Bit_Index_1_adj_2626));
    Odrv4 I__8837 (
            .O(N__39206),
            .I(r_Bit_Index_1_adj_2626));
    Odrv12 I__8836 (
            .O(N__39203),
            .I(r_Bit_Index_1_adj_2626));
    InMux I__8835 (
            .O(N__39194),
            .I(N__39191));
    LocalMux I__8834 (
            .O(N__39191),
            .I(N__39187));
    InMux I__8833 (
            .O(N__39190),
            .I(N__39184));
    Odrv4 I__8832 (
            .O(N__39187),
            .I(data_in_15_0));
    LocalMux I__8831 (
            .O(N__39184),
            .I(data_in_15_0));
    InMux I__8830 (
            .O(N__39179),
            .I(N__39176));
    LocalMux I__8829 (
            .O(N__39176),
            .I(N__39172));
    InMux I__8828 (
            .O(N__39175),
            .I(N__39169));
    Odrv4 I__8827 (
            .O(N__39172),
            .I(data_in_14_0));
    LocalMux I__8826 (
            .O(N__39169),
            .I(data_in_14_0));
    CascadeMux I__8825 (
            .O(N__39164),
            .I(N__39161));
    InMux I__8824 (
            .O(N__39161),
            .I(N__39157));
    CascadeMux I__8823 (
            .O(N__39160),
            .I(N__39154));
    LocalMux I__8822 (
            .O(N__39157),
            .I(N__39151));
    InMux I__8821 (
            .O(N__39154),
            .I(N__39148));
    Odrv12 I__8820 (
            .O(N__39151),
            .I(rand_setpoint_1));
    LocalMux I__8819 (
            .O(N__39148),
            .I(rand_setpoint_1));
    InMux I__8818 (
            .O(N__39143),
            .I(N__39140));
    LocalMux I__8817 (
            .O(N__39140),
            .I(n18438));
    CascadeMux I__8816 (
            .O(N__39137),
            .I(N__39134));
    InMux I__8815 (
            .O(N__39134),
            .I(N__39131));
    LocalMux I__8814 (
            .O(N__39131),
            .I(N__39127));
    InMux I__8813 (
            .O(N__39130),
            .I(N__39119));
    Span4Mux_v I__8812 (
            .O(N__39127),
            .I(N__39116));
    InMux I__8811 (
            .O(N__39126),
            .I(N__39113));
    InMux I__8810 (
            .O(N__39125),
            .I(N__39108));
    InMux I__8809 (
            .O(N__39124),
            .I(N__39108));
    CascadeMux I__8808 (
            .O(N__39123),
            .I(N__39104));
    InMux I__8807 (
            .O(N__39122),
            .I(N__39101));
    LocalMux I__8806 (
            .O(N__39119),
            .I(N__39096));
    Span4Mux_h I__8805 (
            .O(N__39116),
            .I(N__39096));
    LocalMux I__8804 (
            .O(N__39113),
            .I(N__39091));
    LocalMux I__8803 (
            .O(N__39108),
            .I(N__39091));
    InMux I__8802 (
            .O(N__39107),
            .I(N__39086));
    InMux I__8801 (
            .O(N__39104),
            .I(N__39086));
    LocalMux I__8800 (
            .O(N__39101),
            .I(r_Bit_Index_1));
    Odrv4 I__8799 (
            .O(N__39096),
            .I(r_Bit_Index_1));
    Odrv4 I__8798 (
            .O(N__39091),
            .I(r_Bit_Index_1));
    LocalMux I__8797 (
            .O(N__39086),
            .I(r_Bit_Index_1));
    InMux I__8796 (
            .O(N__39077),
            .I(N__39074));
    LocalMux I__8795 (
            .O(N__39074),
            .I(N__39071));
    Odrv4 I__8794 (
            .O(N__39071),
            .I(n18441));
    InMux I__8793 (
            .O(N__39068),
            .I(N__39065));
    LocalMux I__8792 (
            .O(N__39065),
            .I(N__39061));
    InMux I__8791 (
            .O(N__39064),
            .I(N__39058));
    Odrv4 I__8790 (
            .O(N__39061),
            .I(data_in_13_0));
    LocalMux I__8789 (
            .O(N__39058),
            .I(data_in_13_0));
    InMux I__8788 (
            .O(N__39053),
            .I(N__39049));
    InMux I__8787 (
            .O(N__39052),
            .I(N__39046));
    LocalMux I__8786 (
            .O(N__39049),
            .I(r_Tx_Data_3));
    LocalMux I__8785 (
            .O(N__39046),
            .I(r_Tx_Data_3));
    InMux I__8784 (
            .O(N__39041),
            .I(N__39037));
    InMux I__8783 (
            .O(N__39040),
            .I(N__39034));
    LocalMux I__8782 (
            .O(N__39037),
            .I(data_in_20_1));
    LocalMux I__8781 (
            .O(N__39034),
            .I(data_in_20_1));
    InMux I__8780 (
            .O(N__39029),
            .I(N__39023));
    InMux I__8779 (
            .O(N__39028),
            .I(N__39023));
    LocalMux I__8778 (
            .O(N__39023),
            .I(data_in_19_1));
    InMux I__8777 (
            .O(N__39020),
            .I(N__39016));
    InMux I__8776 (
            .O(N__39019),
            .I(N__39013));
    LocalMux I__8775 (
            .O(N__39016),
            .I(data_in_17_0));
    LocalMux I__8774 (
            .O(N__39013),
            .I(data_in_17_0));
    InMux I__8773 (
            .O(N__39008),
            .I(N__39002));
    InMux I__8772 (
            .O(N__39007),
            .I(N__39002));
    LocalMux I__8771 (
            .O(N__39002),
            .I(data_in_16_0));
    CascadeMux I__8770 (
            .O(N__38999),
            .I(n17737_cascade_));
    InMux I__8769 (
            .O(N__38996),
            .I(N__38993));
    LocalMux I__8768 (
            .O(N__38993),
            .I(n17312));
    CascadeMux I__8767 (
            .O(N__38990),
            .I(n17312_cascade_));
    CascadeMux I__8766 (
            .O(N__38987),
            .I(n14_adj_2615_cascade_));
    InMux I__8765 (
            .O(N__38984),
            .I(N__38980));
    InMux I__8764 (
            .O(N__38983),
            .I(N__38977));
    LocalMux I__8763 (
            .O(N__38980),
            .I(data_in_17_1));
    LocalMux I__8762 (
            .O(N__38977),
            .I(data_in_17_1));
    InMux I__8761 (
            .O(N__38972),
            .I(N__38969));
    LocalMux I__8760 (
            .O(N__38969),
            .I(N__38966));
    Span4Mux_h I__8759 (
            .O(N__38966),
            .I(N__38962));
    InMux I__8758 (
            .O(N__38965),
            .I(N__38959));
    Odrv4 I__8757 (
            .O(N__38962),
            .I(data_in_16_1));
    LocalMux I__8756 (
            .O(N__38959),
            .I(data_in_16_1));
    InMux I__8755 (
            .O(N__38954),
            .I(N__38951));
    LocalMux I__8754 (
            .O(N__38951),
            .I(N__38947));
    InMux I__8753 (
            .O(N__38950),
            .I(N__38944));
    Span4Mux_h I__8752 (
            .O(N__38947),
            .I(N__38940));
    LocalMux I__8751 (
            .O(N__38944),
            .I(N__38937));
    InMux I__8750 (
            .O(N__38943),
            .I(N__38934));
    Odrv4 I__8749 (
            .O(N__38940),
            .I(n17757));
    Odrv4 I__8748 (
            .O(N__38937),
            .I(n17757));
    LocalMux I__8747 (
            .O(N__38934),
            .I(n17757));
    CascadeMux I__8746 (
            .O(N__38927),
            .I(N__38922));
    CascadeMux I__8745 (
            .O(N__38926),
            .I(N__38919));
    CascadeMux I__8744 (
            .O(N__38925),
            .I(N__38915));
    InMux I__8743 (
            .O(N__38922),
            .I(N__38912));
    InMux I__8742 (
            .O(N__38919),
            .I(N__38907));
    InMux I__8741 (
            .O(N__38918),
            .I(N__38907));
    InMux I__8740 (
            .O(N__38915),
            .I(N__38902));
    LocalMux I__8739 (
            .O(N__38912),
            .I(N__38899));
    LocalMux I__8738 (
            .O(N__38907),
            .I(N__38896));
    InMux I__8737 (
            .O(N__38906),
            .I(N__38893));
    InMux I__8736 (
            .O(N__38905),
            .I(N__38890));
    LocalMux I__8735 (
            .O(N__38902),
            .I(N__38887));
    Span4Mux_v I__8734 (
            .O(N__38899),
            .I(N__38880));
    Span4Mux_h I__8733 (
            .O(N__38896),
            .I(N__38880));
    LocalMux I__8732 (
            .O(N__38893),
            .I(N__38880));
    LocalMux I__8731 (
            .O(N__38890),
            .I(r_Bit_Index_0));
    Odrv4 I__8730 (
            .O(N__38887),
            .I(r_Bit_Index_0));
    Odrv4 I__8729 (
            .O(N__38880),
            .I(r_Bit_Index_0));
    InMux I__8728 (
            .O(N__38873),
            .I(N__38869));
    InMux I__8727 (
            .O(N__38872),
            .I(N__38866));
    LocalMux I__8726 (
            .O(N__38869),
            .I(data_in_18_1));
    LocalMux I__8725 (
            .O(N__38866),
            .I(data_in_18_1));
    InMux I__8724 (
            .O(N__38861),
            .I(N__38855));
    InMux I__8723 (
            .O(N__38860),
            .I(N__38855));
    LocalMux I__8722 (
            .O(N__38855),
            .I(data_in_19_3));
    InMux I__8721 (
            .O(N__38852),
            .I(N__38846));
    InMux I__8720 (
            .O(N__38851),
            .I(N__38846));
    LocalMux I__8719 (
            .O(N__38846),
            .I(data_in_18_3));
    InMux I__8718 (
            .O(N__38843),
            .I(N__38839));
    InMux I__8717 (
            .O(N__38842),
            .I(N__38836));
    LocalMux I__8716 (
            .O(N__38839),
            .I(N__38833));
    LocalMux I__8715 (
            .O(N__38836),
            .I(data_in_12_0));
    Odrv4 I__8714 (
            .O(N__38833),
            .I(data_in_12_0));
    InMux I__8713 (
            .O(N__38828),
            .I(N__38825));
    LocalMux I__8712 (
            .O(N__38825),
            .I(N__38821));
    InMux I__8711 (
            .O(N__38824),
            .I(N__38818));
    Odrv4 I__8710 (
            .O(N__38821),
            .I(data_in_12_3));
    LocalMux I__8709 (
            .O(N__38818),
            .I(data_in_12_3));
    InMux I__8708 (
            .O(N__38813),
            .I(N__38810));
    LocalMux I__8707 (
            .O(N__38810),
            .I(n18462));
    InMux I__8706 (
            .O(N__38807),
            .I(N__38804));
    LocalMux I__8705 (
            .O(N__38804),
            .I(n18465));
    InMux I__8704 (
            .O(N__38801),
            .I(N__38797));
    InMux I__8703 (
            .O(N__38800),
            .I(N__38794));
    LocalMux I__8702 (
            .O(N__38797),
            .I(N__38791));
    LocalMux I__8701 (
            .O(N__38794),
            .I(N__38787));
    Span4Mux_v I__8700 (
            .O(N__38791),
            .I(N__38784));
    InMux I__8699 (
            .O(N__38790),
            .I(N__38781));
    Span4Mux_h I__8698 (
            .O(N__38787),
            .I(N__38778));
    Span4Mux_h I__8697 (
            .O(N__38784),
            .I(N__38775));
    LocalMux I__8696 (
            .O(N__38781),
            .I(data_in_9_6));
    Odrv4 I__8695 (
            .O(N__38778),
            .I(data_in_9_6));
    Odrv4 I__8694 (
            .O(N__38775),
            .I(data_in_9_6));
    CascadeMux I__8693 (
            .O(N__38768),
            .I(N__38765));
    InMux I__8692 (
            .O(N__38765),
            .I(N__38762));
    LocalMux I__8691 (
            .O(N__38762),
            .I(N__38758));
    InMux I__8690 (
            .O(N__38761),
            .I(N__38755));
    Span4Mux_v I__8689 (
            .O(N__38758),
            .I(N__38752));
    LocalMux I__8688 (
            .O(N__38755),
            .I(N__38749));
    Span4Mux_h I__8687 (
            .O(N__38752),
            .I(N__38744));
    Span4Mux_h I__8686 (
            .O(N__38749),
            .I(N__38744));
    Span4Mux_h I__8685 (
            .O(N__38744),
            .I(N__38740));
    InMux I__8684 (
            .O(N__38743),
            .I(N__38737));
    Odrv4 I__8683 (
            .O(N__38740),
            .I(data_in_8_6));
    LocalMux I__8682 (
            .O(N__38737),
            .I(data_in_8_6));
    InMux I__8681 (
            .O(N__38732),
            .I(N__38729));
    LocalMux I__8680 (
            .O(N__38729),
            .I(N__38726));
    Span4Mux_h I__8679 (
            .O(N__38726),
            .I(N__38722));
    InMux I__8678 (
            .O(N__38725),
            .I(N__38719));
    Odrv4 I__8677 (
            .O(N__38722),
            .I(data_in_16_5));
    LocalMux I__8676 (
            .O(N__38719),
            .I(data_in_16_5));
    InMux I__8675 (
            .O(N__38714),
            .I(N__38710));
    InMux I__8674 (
            .O(N__38713),
            .I(N__38707));
    LocalMux I__8673 (
            .O(N__38710),
            .I(data_in_14_3));
    LocalMux I__8672 (
            .O(N__38707),
            .I(data_in_14_3));
    InMux I__8671 (
            .O(N__38702),
            .I(N__38696));
    InMux I__8670 (
            .O(N__38701),
            .I(N__38696));
    LocalMux I__8669 (
            .O(N__38696),
            .I(data_in_13_3));
    CascadeMux I__8668 (
            .O(N__38693),
            .I(\c0.n18429_cascade_ ));
    InMux I__8667 (
            .O(N__38690),
            .I(N__38687));
    LocalMux I__8666 (
            .O(N__38687),
            .I(N__38684));
    Odrv4 I__8665 (
            .O(N__38684),
            .I(tx_data_7_N_keep));
    CascadeMux I__8664 (
            .O(N__38681),
            .I(\c0.n18017_cascade_ ));
    InMux I__8663 (
            .O(N__38678),
            .I(N__38675));
    LocalMux I__8662 (
            .O(N__38675),
            .I(\c0.n18426 ));
    InMux I__8661 (
            .O(N__38672),
            .I(N__38668));
    InMux I__8660 (
            .O(N__38671),
            .I(N__38665));
    LocalMux I__8659 (
            .O(N__38668),
            .I(data_in_17_3));
    LocalMux I__8658 (
            .O(N__38665),
            .I(data_in_17_3));
    CascadeMux I__8657 (
            .O(N__38660),
            .I(N__38657));
    InMux I__8656 (
            .O(N__38657),
            .I(N__38654));
    LocalMux I__8655 (
            .O(N__38654),
            .I(N__38651));
    Span4Mux_h I__8654 (
            .O(N__38651),
            .I(N__38648));
    Odrv4 I__8653 (
            .O(N__38648),
            .I(\c0.n5_adj_2499 ));
    CascadeMux I__8652 (
            .O(N__38645),
            .I(\c0.n18378_cascade_ ));
    CascadeMux I__8651 (
            .O(N__38642),
            .I(\c0.n18381_cascade_ ));
    InMux I__8650 (
            .O(N__38639),
            .I(N__38636));
    LocalMux I__8649 (
            .O(N__38636),
            .I(tx_data_2_N_keep));
    InMux I__8648 (
            .O(N__38633),
            .I(N__38630));
    LocalMux I__8647 (
            .O(N__38630),
            .I(N__38627));
    Span4Mux_h I__8646 (
            .O(N__38627),
            .I(N__38623));
    InMux I__8645 (
            .O(N__38626),
            .I(N__38620));
    Odrv4 I__8644 (
            .O(N__38623),
            .I(data_in_20_3));
    LocalMux I__8643 (
            .O(N__38620),
            .I(data_in_20_3));
    InMux I__8642 (
            .O(N__38615),
            .I(N__38612));
    LocalMux I__8641 (
            .O(N__38612),
            .I(N__38609));
    Span4Mux_v I__8640 (
            .O(N__38609),
            .I(N__38605));
    InMux I__8639 (
            .O(N__38608),
            .I(N__38602));
    Odrv4 I__8638 (
            .O(N__38605),
            .I(data_in_13_5));
    LocalMux I__8637 (
            .O(N__38602),
            .I(data_in_13_5));
    InMux I__8636 (
            .O(N__38597),
            .I(N__38591));
    InMux I__8635 (
            .O(N__38596),
            .I(N__38591));
    LocalMux I__8634 (
            .O(N__38591),
            .I(data_in_12_4));
    InMux I__8633 (
            .O(N__38588),
            .I(N__38582));
    InMux I__8632 (
            .O(N__38587),
            .I(N__38582));
    LocalMux I__8631 (
            .O(N__38582),
            .I(data_in_13_4));
    InMux I__8630 (
            .O(N__38579),
            .I(N__38573));
    InMux I__8629 (
            .O(N__38578),
            .I(N__38573));
    LocalMux I__8628 (
            .O(N__38573),
            .I(data_in_14_4));
    InMux I__8627 (
            .O(N__38570),
            .I(N__38566));
    InMux I__8626 (
            .O(N__38569),
            .I(N__38563));
    LocalMux I__8625 (
            .O(N__38566),
            .I(data_in_11_3));
    LocalMux I__8624 (
            .O(N__38563),
            .I(data_in_11_3));
    InMux I__8623 (
            .O(N__38558),
            .I(N__38554));
    InMux I__8622 (
            .O(N__38557),
            .I(N__38551));
    LocalMux I__8621 (
            .O(N__38554),
            .I(data_in_15_4));
    LocalMux I__8620 (
            .O(N__38551),
            .I(data_in_15_4));
    InMux I__8619 (
            .O(N__38546),
            .I(N__38543));
    LocalMux I__8618 (
            .O(N__38543),
            .I(N__38540));
    Span4Mux_v I__8617 (
            .O(N__38540),
            .I(N__38537));
    Span4Mux_v I__8616 (
            .O(N__38537),
            .I(N__38533));
    InMux I__8615 (
            .O(N__38536),
            .I(N__38530));
    Odrv4 I__8614 (
            .O(N__38533),
            .I(data_in_17_4));
    LocalMux I__8613 (
            .O(N__38530),
            .I(data_in_17_4));
    InMux I__8612 (
            .O(N__38525),
            .I(N__38521));
    InMux I__8611 (
            .O(N__38524),
            .I(N__38518));
    LocalMux I__8610 (
            .O(N__38521),
            .I(data_in_16_4));
    LocalMux I__8609 (
            .O(N__38518),
            .I(data_in_16_4));
    CascadeMux I__8608 (
            .O(N__38513),
            .I(N__38510));
    InMux I__8607 (
            .O(N__38510),
            .I(N__38507));
    LocalMux I__8606 (
            .O(N__38507),
            .I(N__38503));
    InMux I__8605 (
            .O(N__38506),
            .I(N__38500));
    Span4Mux_h I__8604 (
            .O(N__38503),
            .I(N__38497));
    LocalMux I__8603 (
            .O(N__38500),
            .I(N__38494));
    Span4Mux_h I__8602 (
            .O(N__38497),
            .I(N__38490));
    Span4Mux_h I__8601 (
            .O(N__38494),
            .I(N__38487));
    InMux I__8600 (
            .O(N__38493),
            .I(N__38484));
    Odrv4 I__8599 (
            .O(N__38490),
            .I(data_in_4_1));
    Odrv4 I__8598 (
            .O(N__38487),
            .I(data_in_4_1));
    LocalMux I__8597 (
            .O(N__38484),
            .I(data_in_4_1));
    CascadeMux I__8596 (
            .O(N__38477),
            .I(\c0.n18089_cascade_ ));
    InMux I__8595 (
            .O(N__38474),
            .I(N__38471));
    LocalMux I__8594 (
            .O(N__38471),
            .I(N__38468));
    Span4Mux_s2_v I__8593 (
            .O(N__38468),
            .I(N__38465));
    Span4Mux_h I__8592 (
            .O(N__38465),
            .I(N__38461));
    InMux I__8591 (
            .O(N__38464),
            .I(N__38458));
    Odrv4 I__8590 (
            .O(N__38461),
            .I(data_in_19_2));
    LocalMux I__8589 (
            .O(N__38458),
            .I(data_in_19_2));
    InMux I__8588 (
            .O(N__38453),
            .I(N__38450));
    LocalMux I__8587 (
            .O(N__38450),
            .I(N__38447));
    Span4Mux_s3_v I__8586 (
            .O(N__38447),
            .I(N__38444));
    Span4Mux_h I__8585 (
            .O(N__38444),
            .I(N__38440));
    InMux I__8584 (
            .O(N__38443),
            .I(N__38437));
    Odrv4 I__8583 (
            .O(N__38440),
            .I(data_in_20_4));
    LocalMux I__8582 (
            .O(N__38437),
            .I(data_in_20_4));
    InMux I__8581 (
            .O(N__38432),
            .I(N__38426));
    InMux I__8580 (
            .O(N__38431),
            .I(N__38426));
    LocalMux I__8579 (
            .O(N__38426),
            .I(data_in_19_4));
    InMux I__8578 (
            .O(N__38423),
            .I(N__38417));
    InMux I__8577 (
            .O(N__38422),
            .I(N__38417));
    LocalMux I__8576 (
            .O(N__38417),
            .I(data_in_18_4));
    InMux I__8575 (
            .O(N__38414),
            .I(N__38408));
    InMux I__8574 (
            .O(N__38413),
            .I(N__38408));
    LocalMux I__8573 (
            .O(N__38408),
            .I(data_in_18_2));
    InMux I__8572 (
            .O(N__38405),
            .I(N__38402));
    LocalMux I__8571 (
            .O(N__38402),
            .I(N__38399));
    Span4Mux_h I__8570 (
            .O(N__38399),
            .I(N__38395));
    InMux I__8569 (
            .O(N__38398),
            .I(N__38392));
    Span4Mux_v I__8568 (
            .O(N__38395),
            .I(N__38389));
    LocalMux I__8567 (
            .O(N__38392),
            .I(data_in_17_2));
    Odrv4 I__8566 (
            .O(N__38389),
            .I(data_in_17_2));
    InMux I__8565 (
            .O(N__38384),
            .I(N__38381));
    LocalMux I__8564 (
            .O(N__38381),
            .I(N__38378));
    Span4Mux_v I__8563 (
            .O(N__38378),
            .I(N__38374));
    InMux I__8562 (
            .O(N__38377),
            .I(N__38371));
    Span4Mux_h I__8561 (
            .O(N__38374),
            .I(N__38368));
    LocalMux I__8560 (
            .O(N__38371),
            .I(N__38365));
    Span4Mux_h I__8559 (
            .O(N__38368),
            .I(N__38361));
    Span12Mux_v I__8558 (
            .O(N__38365),
            .I(N__38358));
    InMux I__8557 (
            .O(N__38364),
            .I(N__38355));
    Odrv4 I__8556 (
            .O(N__38361),
            .I(data_in_8_4));
    Odrv12 I__8555 (
            .O(N__38358),
            .I(data_in_8_4));
    LocalMux I__8554 (
            .O(N__38355),
            .I(data_in_8_4));
    InMux I__8553 (
            .O(N__38348),
            .I(N__38343));
    InMux I__8552 (
            .O(N__38347),
            .I(N__38338));
    InMux I__8551 (
            .O(N__38346),
            .I(N__38338));
    LocalMux I__8550 (
            .O(N__38343),
            .I(N__38335));
    LocalMux I__8549 (
            .O(N__38338),
            .I(data_in_9_4));
    Odrv12 I__8548 (
            .O(N__38335),
            .I(data_in_9_4));
    InMux I__8547 (
            .O(N__38330),
            .I(N__38327));
    LocalMux I__8546 (
            .O(N__38327),
            .I(N__38322));
    InMux I__8545 (
            .O(N__38326),
            .I(N__38317));
    InMux I__8544 (
            .O(N__38325),
            .I(N__38317));
    Span4Mux_h I__8543 (
            .O(N__38322),
            .I(N__38314));
    LocalMux I__8542 (
            .O(N__38317),
            .I(data_in_10_4));
    Odrv4 I__8541 (
            .O(N__38314),
            .I(data_in_10_4));
    InMux I__8540 (
            .O(N__38309),
            .I(N__38303));
    InMux I__8539 (
            .O(N__38308),
            .I(N__38303));
    LocalMux I__8538 (
            .O(N__38303),
            .I(data_in_11_4));
    CascadeMux I__8537 (
            .O(N__38300),
            .I(\c0.rx.n18000_cascade_ ));
    CascadeMux I__8536 (
            .O(N__38297),
            .I(N__38294));
    InMux I__8535 (
            .O(N__38294),
            .I(N__38291));
    LocalMux I__8534 (
            .O(N__38291),
            .I(N__38288));
    Span4Mux_h I__8533 (
            .O(N__38288),
            .I(N__38285));
    Odrv4 I__8532 (
            .O(N__38285),
            .I(\c0.rx.n18594 ));
    CascadeMux I__8531 (
            .O(N__38282),
            .I(N__38278));
    InMux I__8530 (
            .O(N__38281),
            .I(N__38275));
    InMux I__8529 (
            .O(N__38278),
            .I(N__38272));
    LocalMux I__8528 (
            .O(N__38275),
            .I(rand_setpoint_27));
    LocalMux I__8527 (
            .O(N__38272),
            .I(rand_setpoint_27));
    CascadeMux I__8526 (
            .O(N__38267),
            .I(\c0.n17966_cascade_ ));
    InMux I__8525 (
            .O(N__38264),
            .I(N__38260));
    InMux I__8524 (
            .O(N__38263),
            .I(N__38257));
    LocalMux I__8523 (
            .O(N__38260),
            .I(rand_setpoint_29));
    LocalMux I__8522 (
            .O(N__38257),
            .I(rand_setpoint_29));
    CascadeMux I__8521 (
            .O(N__38252),
            .I(\c0.n17970_cascade_ ));
    CascadeMux I__8520 (
            .O(N__38249),
            .I(N__38245));
    InMux I__8519 (
            .O(N__38248),
            .I(N__38242));
    InMux I__8518 (
            .O(N__38245),
            .I(N__38239));
    LocalMux I__8517 (
            .O(N__38242),
            .I(rand_setpoint_24));
    LocalMux I__8516 (
            .O(N__38239),
            .I(rand_setpoint_24));
    CascadeMux I__8515 (
            .O(N__38234),
            .I(\c0.n17957_cascade_ ));
    CascadeMux I__8514 (
            .O(N__38231),
            .I(N__38228));
    InMux I__8513 (
            .O(N__38228),
            .I(N__38224));
    InMux I__8512 (
            .O(N__38227),
            .I(N__38221));
    LocalMux I__8511 (
            .O(N__38224),
            .I(rand_setpoint_22));
    LocalMux I__8510 (
            .O(N__38221),
            .I(rand_setpoint_22));
    CascadeMux I__8509 (
            .O(N__38216),
            .I(N__38212));
    InMux I__8508 (
            .O(N__38215),
            .I(N__38209));
    InMux I__8507 (
            .O(N__38212),
            .I(N__38206));
    LocalMux I__8506 (
            .O(N__38209),
            .I(rand_setpoint_4));
    LocalMux I__8505 (
            .O(N__38206),
            .I(rand_setpoint_4));
    InMux I__8504 (
            .O(N__38201),
            .I(N__38195));
    InMux I__8503 (
            .O(N__38200),
            .I(N__38195));
    LocalMux I__8502 (
            .O(N__38195),
            .I(data_in_15_6));
    CascadeMux I__8501 (
            .O(N__38192),
            .I(N__38188));
    InMux I__8500 (
            .O(N__38191),
            .I(N__38185));
    InMux I__8499 (
            .O(N__38188),
            .I(N__38182));
    LocalMux I__8498 (
            .O(N__38185),
            .I(rand_setpoint_11));
    LocalMux I__8497 (
            .O(N__38182),
            .I(rand_setpoint_11));
    InMux I__8496 (
            .O(N__38177),
            .I(N__38173));
    CascadeMux I__8495 (
            .O(N__38176),
            .I(N__38170));
    LocalMux I__8494 (
            .O(N__38173),
            .I(N__38167));
    InMux I__8493 (
            .O(N__38170),
            .I(N__38164));
    Odrv4 I__8492 (
            .O(N__38167),
            .I(rand_setpoint_25));
    LocalMux I__8491 (
            .O(N__38164),
            .I(rand_setpoint_25));
    InMux I__8490 (
            .O(N__38159),
            .I(N__38156));
    LocalMux I__8489 (
            .O(N__38156),
            .I(N__38152));
    InMux I__8488 (
            .O(N__38155),
            .I(N__38149));
    Span4Mux_h I__8487 (
            .O(N__38152),
            .I(N__38146));
    LocalMux I__8486 (
            .O(N__38149),
            .I(rand_setpoint_30));
    Odrv4 I__8485 (
            .O(N__38146),
            .I(rand_setpoint_30));
    InMux I__8484 (
            .O(N__38141),
            .I(N__38137));
    InMux I__8483 (
            .O(N__38140),
            .I(N__38134));
    LocalMux I__8482 (
            .O(N__38137),
            .I(N__38131));
    LocalMux I__8481 (
            .O(N__38134),
            .I(rand_setpoint_31));
    Odrv4 I__8480 (
            .O(N__38131),
            .I(rand_setpoint_31));
    CascadeMux I__8479 (
            .O(N__38126),
            .I(N__38122));
    InMux I__8478 (
            .O(N__38125),
            .I(N__38119));
    InMux I__8477 (
            .O(N__38122),
            .I(N__38116));
    LocalMux I__8476 (
            .O(N__38119),
            .I(rand_setpoint_10));
    LocalMux I__8475 (
            .O(N__38116),
            .I(rand_setpoint_10));
    InMux I__8474 (
            .O(N__38111),
            .I(N__38107));
    CascadeMux I__8473 (
            .O(N__38110),
            .I(N__38103));
    LocalMux I__8472 (
            .O(N__38107),
            .I(N__38097));
    CascadeMux I__8471 (
            .O(N__38106),
            .I(N__38093));
    InMux I__8470 (
            .O(N__38103),
            .I(N__38090));
    InMux I__8469 (
            .O(N__38102),
            .I(N__38087));
    InMux I__8468 (
            .O(N__38101),
            .I(N__38084));
    InMux I__8467 (
            .O(N__38100),
            .I(N__38081));
    Span4Mux_h I__8466 (
            .O(N__38097),
            .I(N__38078));
    InMux I__8465 (
            .O(N__38096),
            .I(N__38073));
    InMux I__8464 (
            .O(N__38093),
            .I(N__38073));
    LocalMux I__8463 (
            .O(N__38090),
            .I(r_Clock_Count_5_adj_2619));
    LocalMux I__8462 (
            .O(N__38087),
            .I(r_Clock_Count_5_adj_2619));
    LocalMux I__8461 (
            .O(N__38084),
            .I(r_Clock_Count_5_adj_2619));
    LocalMux I__8460 (
            .O(N__38081),
            .I(r_Clock_Count_5_adj_2619));
    Odrv4 I__8459 (
            .O(N__38078),
            .I(r_Clock_Count_5_adj_2619));
    LocalMux I__8458 (
            .O(N__38073),
            .I(r_Clock_Count_5_adj_2619));
    InMux I__8457 (
            .O(N__38060),
            .I(N__38057));
    LocalMux I__8456 (
            .O(N__38057),
            .I(N__38051));
    InMux I__8455 (
            .O(N__38056),
            .I(N__38046));
    InMux I__8454 (
            .O(N__38055),
            .I(N__38043));
    InMux I__8453 (
            .O(N__38054),
            .I(N__38040));
    Span4Mux_h I__8452 (
            .O(N__38051),
            .I(N__38037));
    InMux I__8451 (
            .O(N__38050),
            .I(N__38032));
    InMux I__8450 (
            .O(N__38049),
            .I(N__38032));
    LocalMux I__8449 (
            .O(N__38046),
            .I(\c0.rx.r_Clock_Count_7 ));
    LocalMux I__8448 (
            .O(N__38043),
            .I(\c0.rx.r_Clock_Count_7 ));
    LocalMux I__8447 (
            .O(N__38040),
            .I(\c0.rx.r_Clock_Count_7 ));
    Odrv4 I__8446 (
            .O(N__38037),
            .I(\c0.rx.r_Clock_Count_7 ));
    LocalMux I__8445 (
            .O(N__38032),
            .I(\c0.rx.r_Clock_Count_7 ));
    CascadeMux I__8444 (
            .O(N__38021),
            .I(N__38017));
    CascadeMux I__8443 (
            .O(N__38020),
            .I(N__38014));
    InMux I__8442 (
            .O(N__38017),
            .I(N__38011));
    InMux I__8441 (
            .O(N__38014),
            .I(N__38008));
    LocalMux I__8440 (
            .O(N__38011),
            .I(N__38005));
    LocalMux I__8439 (
            .O(N__38008),
            .I(\c0.rx.n97 ));
    Odrv12 I__8438 (
            .O(N__38005),
            .I(\c0.rx.n97 ));
    InMux I__8437 (
            .O(N__38000),
            .I(N__37994));
    InMux I__8436 (
            .O(N__37999),
            .I(N__37989));
    InMux I__8435 (
            .O(N__37998),
            .I(N__37986));
    InMux I__8434 (
            .O(N__37997),
            .I(N__37983));
    LocalMux I__8433 (
            .O(N__37994),
            .I(N__37980));
    InMux I__8432 (
            .O(N__37993),
            .I(N__37975));
    InMux I__8431 (
            .O(N__37992),
            .I(N__37975));
    LocalMux I__8430 (
            .O(N__37989),
            .I(\c0.rx.r_Clock_Count_6 ));
    LocalMux I__8429 (
            .O(N__37986),
            .I(\c0.rx.r_Clock_Count_6 ));
    LocalMux I__8428 (
            .O(N__37983),
            .I(\c0.rx.r_Clock_Count_6 ));
    Odrv12 I__8427 (
            .O(N__37980),
            .I(\c0.rx.r_Clock_Count_6 ));
    LocalMux I__8426 (
            .O(N__37975),
            .I(\c0.rx.r_Clock_Count_6 ));
    CascadeMux I__8425 (
            .O(N__37964),
            .I(\c0.rx.r_SM_Main_2_N_2380_2_cascade_ ));
    InMux I__8424 (
            .O(N__37961),
            .I(N__37958));
    LocalMux I__8423 (
            .O(N__37958),
            .I(\c0.n18498 ));
    CascadeMux I__8422 (
            .O(N__37955),
            .I(\c0.n2_adj_2487_cascade_ ));
    InMux I__8421 (
            .O(N__37952),
            .I(N__37949));
    LocalMux I__8420 (
            .O(N__37949),
            .I(n4_adj_2649));
    CascadeMux I__8419 (
            .O(N__37946),
            .I(N__37942));
    InMux I__8418 (
            .O(N__37945),
            .I(N__37938));
    InMux I__8417 (
            .O(N__37942),
            .I(N__37933));
    InMux I__8416 (
            .O(N__37941),
            .I(N__37933));
    LocalMux I__8415 (
            .O(N__37938),
            .I(N__37930));
    LocalMux I__8414 (
            .O(N__37933),
            .I(N__37927));
    Odrv12 I__8413 (
            .O(N__37930),
            .I(n8562));
    Odrv4 I__8412 (
            .O(N__37927),
            .I(n8562));
    CascadeMux I__8411 (
            .O(N__37922),
            .I(n4_adj_2649_cascade_));
    InMux I__8410 (
            .O(N__37919),
            .I(N__37911));
    InMux I__8409 (
            .O(N__37918),
            .I(N__37902));
    InMux I__8408 (
            .O(N__37917),
            .I(N__37902));
    InMux I__8407 (
            .O(N__37916),
            .I(N__37902));
    InMux I__8406 (
            .O(N__37915),
            .I(N__37899));
    InMux I__8405 (
            .O(N__37914),
            .I(N__37896));
    LocalMux I__8404 (
            .O(N__37911),
            .I(N__37891));
    InMux I__8403 (
            .O(N__37910),
            .I(N__37888));
    InMux I__8402 (
            .O(N__37909),
            .I(N__37885));
    LocalMux I__8401 (
            .O(N__37902),
            .I(N__37882));
    LocalMux I__8400 (
            .O(N__37899),
            .I(N__37877));
    LocalMux I__8399 (
            .O(N__37896),
            .I(N__37877));
    CascadeMux I__8398 (
            .O(N__37895),
            .I(N__37873));
    InMux I__8397 (
            .O(N__37894),
            .I(N__37870));
    Span4Mux_h I__8396 (
            .O(N__37891),
            .I(N__37867));
    LocalMux I__8395 (
            .O(N__37888),
            .I(N__37862));
    LocalMux I__8394 (
            .O(N__37885),
            .I(N__37862));
    Span4Mux_h I__8393 (
            .O(N__37882),
            .I(N__37859));
    Span4Mux_h I__8392 (
            .O(N__37877),
            .I(N__37856));
    InMux I__8391 (
            .O(N__37876),
            .I(N__37851));
    InMux I__8390 (
            .O(N__37873),
            .I(N__37851));
    LocalMux I__8389 (
            .O(N__37870),
            .I(r_Rx_Data));
    Odrv4 I__8388 (
            .O(N__37867),
            .I(r_Rx_Data));
    Odrv12 I__8387 (
            .O(N__37862),
            .I(r_Rx_Data));
    Odrv4 I__8386 (
            .O(N__37859),
            .I(r_Rx_Data));
    Odrv4 I__8385 (
            .O(N__37856),
            .I(r_Rx_Data));
    LocalMux I__8384 (
            .O(N__37851),
            .I(r_Rx_Data));
    InMux I__8383 (
            .O(N__37838),
            .I(N__37835));
    LocalMux I__8382 (
            .O(N__37835),
            .I(N__37831));
    InMux I__8381 (
            .O(N__37834),
            .I(N__37828));
    Odrv4 I__8380 (
            .O(N__37831),
            .I(rx_data_0));
    LocalMux I__8379 (
            .O(N__37828),
            .I(rx_data_0));
    InMux I__8378 (
            .O(N__37823),
            .I(N__37820));
    LocalMux I__8377 (
            .O(N__37820),
            .I(N__37816));
    InMux I__8376 (
            .O(N__37819),
            .I(N__37813));
    Odrv12 I__8375 (
            .O(N__37816),
            .I(data_in_20_0));
    LocalMux I__8374 (
            .O(N__37813),
            .I(data_in_20_0));
    InMux I__8373 (
            .O(N__37808),
            .I(N__37805));
    LocalMux I__8372 (
            .O(N__37805),
            .I(N__37801));
    InMux I__8371 (
            .O(N__37804),
            .I(N__37798));
    Odrv4 I__8370 (
            .O(N__37801),
            .I(data_in_17_6));
    LocalMux I__8369 (
            .O(N__37798),
            .I(data_in_17_6));
    InMux I__8368 (
            .O(N__37793),
            .I(N__37787));
    InMux I__8367 (
            .O(N__37792),
            .I(N__37787));
    LocalMux I__8366 (
            .O(N__37787),
            .I(data_in_16_6));
    InMux I__8365 (
            .O(N__37784),
            .I(N__37781));
    LocalMux I__8364 (
            .O(N__37781),
            .I(N__37778));
    Odrv4 I__8363 (
            .O(N__37778),
            .I(\c0.n6_adj_2448 ));
    InMux I__8362 (
            .O(N__37775),
            .I(N__37771));
    InMux I__8361 (
            .O(N__37774),
            .I(N__37768));
    LocalMux I__8360 (
            .O(N__37771),
            .I(data_in_19_6));
    LocalMux I__8359 (
            .O(N__37768),
            .I(data_in_19_6));
    InMux I__8358 (
            .O(N__37763),
            .I(N__37757));
    InMux I__8357 (
            .O(N__37762),
            .I(N__37757));
    LocalMux I__8356 (
            .O(N__37757),
            .I(data_in_18_6));
    CascadeMux I__8355 (
            .O(N__37754),
            .I(N__37750));
    InMux I__8354 (
            .O(N__37753),
            .I(N__37747));
    InMux I__8353 (
            .O(N__37750),
            .I(N__37744));
    LocalMux I__8352 (
            .O(N__37747),
            .I(rx_data_1));
    LocalMux I__8351 (
            .O(N__37744),
            .I(rx_data_1));
    InMux I__8350 (
            .O(N__37739),
            .I(N__37735));
    CascadeMux I__8349 (
            .O(N__37738),
            .I(N__37732));
    LocalMux I__8348 (
            .O(N__37735),
            .I(N__37729));
    InMux I__8347 (
            .O(N__37732),
            .I(N__37726));
    Odrv4 I__8346 (
            .O(N__37729),
            .I(rand_setpoint_2));
    LocalMux I__8345 (
            .O(N__37726),
            .I(rand_setpoint_2));
    InMux I__8344 (
            .O(N__37721),
            .I(N__37718));
    LocalMux I__8343 (
            .O(N__37718),
            .I(N__37714));
    InMux I__8342 (
            .O(N__37717),
            .I(N__37711));
    Odrv12 I__8341 (
            .O(N__37714),
            .I(data_in_19_5));
    LocalMux I__8340 (
            .O(N__37711),
            .I(data_in_19_5));
    InMux I__8339 (
            .O(N__37706),
            .I(N__37703));
    LocalMux I__8338 (
            .O(N__37703),
            .I(N__37699));
    InMux I__8337 (
            .O(N__37702),
            .I(N__37696));
    Odrv4 I__8336 (
            .O(N__37699),
            .I(rx_data_5));
    LocalMux I__8335 (
            .O(N__37696),
            .I(rx_data_5));
    InMux I__8334 (
            .O(N__37691),
            .I(N__37685));
    InMux I__8333 (
            .O(N__37690),
            .I(N__37685));
    LocalMux I__8332 (
            .O(N__37685),
            .I(data_in_20_5));
    InMux I__8331 (
            .O(N__37682),
            .I(N__37679));
    LocalMux I__8330 (
            .O(N__37679),
            .I(N__37676));
    Odrv4 I__8329 (
            .O(N__37676),
            .I(\c0.n17911 ));
    CascadeMux I__8328 (
            .O(N__37673),
            .I(N__37670));
    InMux I__8327 (
            .O(N__37670),
            .I(N__37667));
    LocalMux I__8326 (
            .O(N__37667),
            .I(\c0.n5_adj_2488 ));
    CascadeMux I__8325 (
            .O(N__37664),
            .I(\c0.n17556_cascade_ ));
    InMux I__8324 (
            .O(N__37661),
            .I(N__37657));
    InMux I__8323 (
            .O(N__37660),
            .I(N__37653));
    LocalMux I__8322 (
            .O(N__37657),
            .I(N__37649));
    InMux I__8321 (
            .O(N__37656),
            .I(N__37645));
    LocalMux I__8320 (
            .O(N__37653),
            .I(N__37642));
    InMux I__8319 (
            .O(N__37652),
            .I(N__37639));
    Span4Mux_h I__8318 (
            .O(N__37649),
            .I(N__37636));
    InMux I__8317 (
            .O(N__37648),
            .I(N__37633));
    LocalMux I__8316 (
            .O(N__37645),
            .I(N__37630));
    Sp12to4 I__8315 (
            .O(N__37642),
            .I(N__37625));
    LocalMux I__8314 (
            .O(N__37639),
            .I(N__37625));
    Odrv4 I__8313 (
            .O(N__37636),
            .I(data_in_1_4));
    LocalMux I__8312 (
            .O(N__37633),
            .I(data_in_1_4));
    Odrv12 I__8311 (
            .O(N__37630),
            .I(data_in_1_4));
    Odrv12 I__8310 (
            .O(N__37625),
            .I(data_in_1_4));
    InMux I__8309 (
            .O(N__37616),
            .I(N__37613));
    LocalMux I__8308 (
            .O(N__37613),
            .I(N__37609));
    CascadeMux I__8307 (
            .O(N__37612),
            .I(N__37605));
    Span4Mux_v I__8306 (
            .O(N__37609),
            .I(N__37601));
    InMux I__8305 (
            .O(N__37608),
            .I(N__37598));
    InMux I__8304 (
            .O(N__37605),
            .I(N__37595));
    InMux I__8303 (
            .O(N__37604),
            .I(N__37592));
    Span4Mux_h I__8302 (
            .O(N__37601),
            .I(N__37589));
    LocalMux I__8301 (
            .O(N__37598),
            .I(N__37586));
    LocalMux I__8300 (
            .O(N__37595),
            .I(N__37583));
    LocalMux I__8299 (
            .O(N__37592),
            .I(data_in_0_5));
    Odrv4 I__8298 (
            .O(N__37589),
            .I(data_in_0_5));
    Odrv12 I__8297 (
            .O(N__37586),
            .I(data_in_0_5));
    Odrv12 I__8296 (
            .O(N__37583),
            .I(data_in_0_5));
    CascadeMux I__8295 (
            .O(N__37574),
            .I(N__37570));
    InMux I__8294 (
            .O(N__37573),
            .I(N__37567));
    InMux I__8293 (
            .O(N__37570),
            .I(N__37563));
    LocalMux I__8292 (
            .O(N__37567),
            .I(N__37560));
    InMux I__8291 (
            .O(N__37566),
            .I(N__37557));
    LocalMux I__8290 (
            .O(N__37563),
            .I(N__37554));
    Span4Mux_v I__8289 (
            .O(N__37560),
            .I(N__37547));
    LocalMux I__8288 (
            .O(N__37557),
            .I(N__37547));
    Span4Mux_h I__8287 (
            .O(N__37554),
            .I(N__37544));
    CascadeMux I__8286 (
            .O(N__37553),
            .I(N__37541));
    InMux I__8285 (
            .O(N__37552),
            .I(N__37538));
    Span4Mux_h I__8284 (
            .O(N__37547),
            .I(N__37533));
    Span4Mux_v I__8283 (
            .O(N__37544),
            .I(N__37533));
    InMux I__8282 (
            .O(N__37541),
            .I(N__37530));
    LocalMux I__8281 (
            .O(N__37538),
            .I(data_in_2_3));
    Odrv4 I__8280 (
            .O(N__37533),
            .I(data_in_2_3));
    LocalMux I__8279 (
            .O(N__37530),
            .I(data_in_2_3));
    InMux I__8278 (
            .O(N__37523),
            .I(N__37520));
    LocalMux I__8277 (
            .O(N__37520),
            .I(N__37515));
    InMux I__8276 (
            .O(N__37519),
            .I(N__37512));
    InMux I__8275 (
            .O(N__37518),
            .I(N__37509));
    Span4Mux_v I__8274 (
            .O(N__37515),
            .I(N__37504));
    LocalMux I__8273 (
            .O(N__37512),
            .I(N__37501));
    LocalMux I__8272 (
            .O(N__37509),
            .I(N__37498));
    InMux I__8271 (
            .O(N__37508),
            .I(N__37495));
    InMux I__8270 (
            .O(N__37507),
            .I(N__37492));
    Span4Mux_h I__8269 (
            .O(N__37504),
            .I(N__37489));
    Span4Mux_v I__8268 (
            .O(N__37501),
            .I(N__37486));
    Span12Mux_s6_h I__8267 (
            .O(N__37498),
            .I(N__37481));
    LocalMux I__8266 (
            .O(N__37495),
            .I(N__37481));
    LocalMux I__8265 (
            .O(N__37492),
            .I(data_in_3_2));
    Odrv4 I__8264 (
            .O(N__37489),
            .I(data_in_3_2));
    Odrv4 I__8263 (
            .O(N__37486),
            .I(data_in_3_2));
    Odrv12 I__8262 (
            .O(N__37481),
            .I(data_in_3_2));
    InMux I__8261 (
            .O(N__37472),
            .I(N__37469));
    LocalMux I__8260 (
            .O(N__37469),
            .I(N__37466));
    Span4Mux_h I__8259 (
            .O(N__37466),
            .I(N__37463));
    Span4Mux_h I__8258 (
            .O(N__37463),
            .I(N__37460));
    Odrv4 I__8257 (
            .O(N__37460),
            .I(\c0.n16_adj_2513 ));
    InMux I__8256 (
            .O(N__37457),
            .I(N__37454));
    LocalMux I__8255 (
            .O(N__37454),
            .I(N__37450));
    InMux I__8254 (
            .O(N__37453),
            .I(N__37447));
    Odrv4 I__8253 (
            .O(N__37450),
            .I(data_in_18_0));
    LocalMux I__8252 (
            .O(N__37447),
            .I(data_in_18_0));
    InMux I__8251 (
            .O(N__37442),
            .I(N__37437));
    InMux I__8250 (
            .O(N__37441),
            .I(N__37434));
    InMux I__8249 (
            .O(N__37440),
            .I(N__37431));
    LocalMux I__8248 (
            .O(N__37437),
            .I(N__37428));
    LocalMux I__8247 (
            .O(N__37434),
            .I(N__37425));
    LocalMux I__8246 (
            .O(N__37431),
            .I(n9796));
    Odrv4 I__8245 (
            .O(N__37428),
            .I(n9796));
    Odrv4 I__8244 (
            .O(N__37425),
            .I(n9796));
    InMux I__8243 (
            .O(N__37418),
            .I(N__37414));
    InMux I__8242 (
            .O(N__37417),
            .I(N__37411));
    LocalMux I__8241 (
            .O(N__37414),
            .I(N__37408));
    LocalMux I__8240 (
            .O(N__37411),
            .I(r_Tx_Data_7));
    Odrv12 I__8239 (
            .O(N__37408),
            .I(r_Tx_Data_7));
    CascadeMux I__8238 (
            .O(N__37403),
            .I(N__37399));
    InMux I__8237 (
            .O(N__37402),
            .I(N__37390));
    InMux I__8236 (
            .O(N__37399),
            .I(N__37390));
    InMux I__8235 (
            .O(N__37398),
            .I(N__37385));
    InMux I__8234 (
            .O(N__37397),
            .I(N__37385));
    InMux I__8233 (
            .O(N__37396),
            .I(N__37382));
    InMux I__8232 (
            .O(N__37395),
            .I(N__37379));
    LocalMux I__8231 (
            .O(N__37390),
            .I(N__37376));
    LocalMux I__8230 (
            .O(N__37385),
            .I(N__37373));
    LocalMux I__8229 (
            .O(N__37382),
            .I(r_Bit_Index_2));
    LocalMux I__8228 (
            .O(N__37379),
            .I(r_Bit_Index_2));
    Odrv12 I__8227 (
            .O(N__37376),
            .I(r_Bit_Index_2));
    Odrv4 I__8226 (
            .O(N__37373),
            .I(r_Bit_Index_2));
    InMux I__8225 (
            .O(N__37364),
            .I(N__37359));
    InMux I__8224 (
            .O(N__37363),
            .I(N__37354));
    InMux I__8223 (
            .O(N__37362),
            .I(N__37354));
    LocalMux I__8222 (
            .O(N__37359),
            .I(N__37351));
    LocalMux I__8221 (
            .O(N__37354),
            .I(n12_adj_2618));
    Odrv4 I__8220 (
            .O(N__37351),
            .I(n12_adj_2618));
    InMux I__8219 (
            .O(N__37346),
            .I(N__37343));
    LocalMux I__8218 (
            .O(N__37343),
            .I(N__37340));
    Span4Mux_h I__8217 (
            .O(N__37340),
            .I(N__37337));
    Odrv4 I__8216 (
            .O(N__37337),
            .I(n22));
    InMux I__8215 (
            .O(N__37334),
            .I(N__37331));
    LocalMux I__8214 (
            .O(N__37331),
            .I(N__37328));
    Odrv12 I__8213 (
            .O(N__37328),
            .I(n17950));
    InMux I__8212 (
            .O(N__37325),
            .I(N__37322));
    LocalMux I__8211 (
            .O(N__37322),
            .I(N__37316));
    InMux I__8210 (
            .O(N__37321),
            .I(N__37312));
    InMux I__8209 (
            .O(N__37320),
            .I(N__37309));
    InMux I__8208 (
            .O(N__37319),
            .I(N__37306));
    Span4Mux_h I__8207 (
            .O(N__37316),
            .I(N__37303));
    InMux I__8206 (
            .O(N__37315),
            .I(N__37300));
    LocalMux I__8205 (
            .O(N__37312),
            .I(N__37295));
    LocalMux I__8204 (
            .O(N__37309),
            .I(N__37295));
    LocalMux I__8203 (
            .O(N__37306),
            .I(r_Clock_Count_8));
    Odrv4 I__8202 (
            .O(N__37303),
            .I(r_Clock_Count_8));
    LocalMux I__8201 (
            .O(N__37300),
            .I(r_Clock_Count_8));
    Odrv4 I__8200 (
            .O(N__37295),
            .I(r_Clock_Count_8));
    InMux I__8199 (
            .O(N__37286),
            .I(N__37283));
    LocalMux I__8198 (
            .O(N__37283),
            .I(n17767));
    InMux I__8197 (
            .O(N__37280),
            .I(N__37277));
    LocalMux I__8196 (
            .O(N__37277),
            .I(\c0.tx.n17 ));
    InMux I__8195 (
            .O(N__37274),
            .I(N__37268));
    InMux I__8194 (
            .O(N__37273),
            .I(N__37268));
    LocalMux I__8193 (
            .O(N__37268),
            .I(r_Tx_Data_2));
    InMux I__8192 (
            .O(N__37265),
            .I(N__37262));
    LocalMux I__8191 (
            .O(N__37262),
            .I(N__37258));
    CascadeMux I__8190 (
            .O(N__37261),
            .I(N__37255));
    Span4Mux_h I__8189 (
            .O(N__37258),
            .I(N__37249));
    InMux I__8188 (
            .O(N__37255),
            .I(N__37246));
    InMux I__8187 (
            .O(N__37254),
            .I(N__37241));
    InMux I__8186 (
            .O(N__37253),
            .I(N__37241));
    InMux I__8185 (
            .O(N__37252),
            .I(N__37238));
    Odrv4 I__8184 (
            .O(N__37249),
            .I(r_Clock_Count_6));
    LocalMux I__8183 (
            .O(N__37246),
            .I(r_Clock_Count_6));
    LocalMux I__8182 (
            .O(N__37241),
            .I(r_Clock_Count_6));
    LocalMux I__8181 (
            .O(N__37238),
            .I(r_Clock_Count_6));
    InMux I__8180 (
            .O(N__37229),
            .I(N__37226));
    LocalMux I__8179 (
            .O(N__37226),
            .I(N__37223));
    Span4Mux_v I__8178 (
            .O(N__37223),
            .I(N__37219));
    InMux I__8177 (
            .O(N__37222),
            .I(N__37216));
    Span4Mux_h I__8176 (
            .O(N__37219),
            .I(N__37210));
    LocalMux I__8175 (
            .O(N__37216),
            .I(N__37210));
    InMux I__8174 (
            .O(N__37215),
            .I(N__37206));
    Span4Mux_v I__8173 (
            .O(N__37210),
            .I(N__37203));
    InMux I__8172 (
            .O(N__37209),
            .I(N__37200));
    LocalMux I__8171 (
            .O(N__37206),
            .I(N__37192));
    Sp12to4 I__8170 (
            .O(N__37203),
            .I(N__37192));
    LocalMux I__8169 (
            .O(N__37200),
            .I(N__37192));
    InMux I__8168 (
            .O(N__37199),
            .I(N__37189));
    Span12Mux_h I__8167 (
            .O(N__37192),
            .I(N__37186));
    LocalMux I__8166 (
            .O(N__37189),
            .I(r_Clock_Count_7));
    Odrv12 I__8165 (
            .O(N__37186),
            .I(r_Clock_Count_7));
    CascadeMux I__8164 (
            .O(N__37181),
            .I(n1_cascade_));
    CascadeMux I__8163 (
            .O(N__37178),
            .I(n3_adj_2650_cascade_));
    IoInMux I__8162 (
            .O(N__37175),
            .I(N__37172));
    LocalMux I__8161 (
            .O(N__37172),
            .I(N__37169));
    IoSpan4Mux I__8160 (
            .O(N__37169),
            .I(N__37166));
    Span4Mux_s0_v I__8159 (
            .O(N__37166),
            .I(N__37163));
    Span4Mux_h I__8158 (
            .O(N__37163),
            .I(N__37159));
    InMux I__8157 (
            .O(N__37162),
            .I(N__37156));
    Span4Mux_s0_v I__8156 (
            .O(N__37159),
            .I(N__37151));
    LocalMux I__8155 (
            .O(N__37156),
            .I(N__37151));
    Span4Mux_v I__8154 (
            .O(N__37151),
            .I(N__37148));
    Span4Mux_v I__8153 (
            .O(N__37148),
            .I(N__37145));
    Span4Mux_h I__8152 (
            .O(N__37145),
            .I(N__37141));
    InMux I__8151 (
            .O(N__37144),
            .I(N__37138));
    Odrv4 I__8150 (
            .O(N__37141),
            .I(tx_o_adj_2584));
    LocalMux I__8149 (
            .O(N__37138),
            .I(tx_o_adj_2584));
    InMux I__8148 (
            .O(N__37133),
            .I(N__37129));
    InMux I__8147 (
            .O(N__37132),
            .I(N__37126));
    LocalMux I__8146 (
            .O(N__37129),
            .I(data_in_18_7));
    LocalMux I__8145 (
            .O(N__37126),
            .I(data_in_18_7));
    InMux I__8144 (
            .O(N__37121),
            .I(N__37118));
    LocalMux I__8143 (
            .O(N__37118),
            .I(N__37114));
    InMux I__8142 (
            .O(N__37117),
            .I(N__37111));
    Odrv4 I__8141 (
            .O(N__37114),
            .I(rx_data_7));
    LocalMux I__8140 (
            .O(N__37111),
            .I(rx_data_7));
    InMux I__8139 (
            .O(N__37106),
            .I(N__37103));
    LocalMux I__8138 (
            .O(N__37103),
            .I(N__37099));
    InMux I__8137 (
            .O(N__37102),
            .I(N__37096));
    Odrv4 I__8136 (
            .O(N__37099),
            .I(data_in_16_3));
    LocalMux I__8135 (
            .O(N__37096),
            .I(data_in_16_3));
    InMux I__8134 (
            .O(N__37091),
            .I(N__37088));
    LocalMux I__8133 (
            .O(N__37088),
            .I(N__37084));
    InMux I__8132 (
            .O(N__37087),
            .I(N__37081));
    Odrv4 I__8131 (
            .O(N__37084),
            .I(data_in_15_3));
    LocalMux I__8130 (
            .O(N__37081),
            .I(data_in_15_3));
    InMux I__8129 (
            .O(N__37076),
            .I(N__37070));
    InMux I__8128 (
            .O(N__37075),
            .I(N__37070));
    LocalMux I__8127 (
            .O(N__37070),
            .I(data_in_20_7));
    InMux I__8126 (
            .O(N__37067),
            .I(N__37063));
    InMux I__8125 (
            .O(N__37066),
            .I(N__37060));
    LocalMux I__8124 (
            .O(N__37063),
            .I(data_in_19_7));
    LocalMux I__8123 (
            .O(N__37060),
            .I(data_in_19_7));
    InMux I__8122 (
            .O(N__37055),
            .I(N__37052));
    LocalMux I__8121 (
            .O(N__37052),
            .I(n12123));
    InMux I__8120 (
            .O(N__37049),
            .I(N__37046));
    LocalMux I__8119 (
            .O(N__37046),
            .I(n7080));
    InMux I__8118 (
            .O(N__37043),
            .I(N__37039));
    InMux I__8117 (
            .O(N__37042),
            .I(N__37036));
    LocalMux I__8116 (
            .O(N__37039),
            .I(N__37033));
    LocalMux I__8115 (
            .O(N__37036),
            .I(N__37029));
    Span4Mux_h I__8114 (
            .O(N__37033),
            .I(N__37026));
    InMux I__8113 (
            .O(N__37032),
            .I(N__37023));
    Odrv12 I__8112 (
            .O(N__37029),
            .I(data_in_8_1));
    Odrv4 I__8111 (
            .O(N__37026),
            .I(data_in_8_1));
    LocalMux I__8110 (
            .O(N__37023),
            .I(data_in_8_1));
    InMux I__8109 (
            .O(N__37016),
            .I(N__37012));
    InMux I__8108 (
            .O(N__37015),
            .I(N__37009));
    LocalMux I__8107 (
            .O(N__37012),
            .I(N__37005));
    LocalMux I__8106 (
            .O(N__37009),
            .I(N__37002));
    InMux I__8105 (
            .O(N__37008),
            .I(N__36999));
    Span4Mux_h I__8104 (
            .O(N__37005),
            .I(N__36996));
    Odrv4 I__8103 (
            .O(N__37002),
            .I(\c0.data_in_7_1 ));
    LocalMux I__8102 (
            .O(N__36999),
            .I(\c0.data_in_7_1 ));
    Odrv4 I__8101 (
            .O(N__36996),
            .I(\c0.data_in_7_1 ));
    CascadeMux I__8100 (
            .O(N__36989),
            .I(N__36986));
    InMux I__8099 (
            .O(N__36986),
            .I(N__36983));
    LocalMux I__8098 (
            .O(N__36983),
            .I(N__36979));
    InMux I__8097 (
            .O(N__36982),
            .I(N__36975));
    Span4Mux_v I__8096 (
            .O(N__36979),
            .I(N__36972));
    InMux I__8095 (
            .O(N__36978),
            .I(N__36969));
    LocalMux I__8094 (
            .O(N__36975),
            .I(data_in_10_3));
    Odrv4 I__8093 (
            .O(N__36972),
            .I(data_in_10_3));
    LocalMux I__8092 (
            .O(N__36969),
            .I(data_in_10_3));
    InMux I__8091 (
            .O(N__36962),
            .I(N__36958));
    CascadeMux I__8090 (
            .O(N__36961),
            .I(N__36955));
    LocalMux I__8089 (
            .O(N__36958),
            .I(N__36952));
    InMux I__8088 (
            .O(N__36955),
            .I(N__36949));
    Span4Mux_v I__8087 (
            .O(N__36952),
            .I(N__36944));
    LocalMux I__8086 (
            .O(N__36949),
            .I(N__36941));
    InMux I__8085 (
            .O(N__36948),
            .I(N__36938));
    InMux I__8084 (
            .O(N__36947),
            .I(N__36935));
    Span4Mux_h I__8083 (
            .O(N__36944),
            .I(N__36930));
    Span4Mux_v I__8082 (
            .O(N__36941),
            .I(N__36930));
    LocalMux I__8081 (
            .O(N__36938),
            .I(data_in_6_7));
    LocalMux I__8080 (
            .O(N__36935),
            .I(data_in_6_7));
    Odrv4 I__8079 (
            .O(N__36930),
            .I(data_in_6_7));
    CascadeMux I__8078 (
            .O(N__36923),
            .I(N__36920));
    InMux I__8077 (
            .O(N__36920),
            .I(N__36917));
    LocalMux I__8076 (
            .O(N__36917),
            .I(N__36913));
    InMux I__8075 (
            .O(N__36916),
            .I(N__36909));
    Span4Mux_v I__8074 (
            .O(N__36913),
            .I(N__36906));
    CascadeMux I__8073 (
            .O(N__36912),
            .I(N__36903));
    LocalMux I__8072 (
            .O(N__36909),
            .I(N__36899));
    Span4Mux_h I__8071 (
            .O(N__36906),
            .I(N__36896));
    InMux I__8070 (
            .O(N__36903),
            .I(N__36893));
    InMux I__8069 (
            .O(N__36902),
            .I(N__36890));
    Span4Mux_h I__8068 (
            .O(N__36899),
            .I(N__36887));
    Span4Mux_h I__8067 (
            .O(N__36896),
            .I(N__36884));
    LocalMux I__8066 (
            .O(N__36893),
            .I(N__36881));
    LocalMux I__8065 (
            .O(N__36890),
            .I(data_in_5_7));
    Odrv4 I__8064 (
            .O(N__36887),
            .I(data_in_5_7));
    Odrv4 I__8063 (
            .O(N__36884),
            .I(data_in_5_7));
    Odrv12 I__8062 (
            .O(N__36881),
            .I(data_in_5_7));
    InMux I__8061 (
            .O(N__36872),
            .I(N__36868));
    CascadeMux I__8060 (
            .O(N__36871),
            .I(N__36865));
    LocalMux I__8059 (
            .O(N__36868),
            .I(N__36862));
    InMux I__8058 (
            .O(N__36865),
            .I(N__36859));
    Span4Mux_v I__8057 (
            .O(N__36862),
            .I(N__36852));
    LocalMux I__8056 (
            .O(N__36859),
            .I(N__36852));
    InMux I__8055 (
            .O(N__36858),
            .I(N__36849));
    InMux I__8054 (
            .O(N__36857),
            .I(N__36846));
    Span4Mux_h I__8053 (
            .O(N__36852),
            .I(N__36843));
    LocalMux I__8052 (
            .O(N__36849),
            .I(\c0.data_in_frame_10_1 ));
    LocalMux I__8051 (
            .O(N__36846),
            .I(\c0.data_in_frame_10_1 ));
    Odrv4 I__8050 (
            .O(N__36843),
            .I(\c0.data_in_frame_10_1 ));
    CascadeMux I__8049 (
            .O(N__36836),
            .I(N__36833));
    InMux I__8048 (
            .O(N__36833),
            .I(N__36828));
    InMux I__8047 (
            .O(N__36832),
            .I(N__36825));
    InMux I__8046 (
            .O(N__36831),
            .I(N__36822));
    LocalMux I__8045 (
            .O(N__36828),
            .I(N__36819));
    LocalMux I__8044 (
            .O(N__36825),
            .I(N__36814));
    LocalMux I__8043 (
            .O(N__36822),
            .I(N__36814));
    Span4Mux_h I__8042 (
            .O(N__36819),
            .I(N__36811));
    Odrv12 I__8041 (
            .O(N__36814),
            .I(\c0.data_in_frame_10_3 ));
    Odrv4 I__8040 (
            .O(N__36811),
            .I(\c0.data_in_frame_10_3 ));
    CascadeMux I__8039 (
            .O(N__36806),
            .I(N__36803));
    InMux I__8038 (
            .O(N__36803),
            .I(N__36800));
    LocalMux I__8037 (
            .O(N__36800),
            .I(N__36797));
    Span4Mux_h I__8036 (
            .O(N__36797),
            .I(N__36794));
    Span4Mux_h I__8035 (
            .O(N__36794),
            .I(N__36791));
    Span4Mux_v I__8034 (
            .O(N__36791),
            .I(N__36788));
    Odrv4 I__8033 (
            .O(N__36788),
            .I(\c0.n6 ));
    InMux I__8032 (
            .O(N__36785),
            .I(N__36782));
    LocalMux I__8031 (
            .O(N__36782),
            .I(N__36779));
    Span4Mux_v I__8030 (
            .O(N__36779),
            .I(N__36775));
    InMux I__8029 (
            .O(N__36778),
            .I(N__36772));
    Odrv4 I__8028 (
            .O(N__36775),
            .I(data_in_11_0));
    LocalMux I__8027 (
            .O(N__36772),
            .I(data_in_11_0));
    InMux I__8026 (
            .O(N__36767),
            .I(N__36764));
    LocalMux I__8025 (
            .O(N__36764),
            .I(n7086));
    InMux I__8024 (
            .O(N__36761),
            .I(N__36758));
    LocalMux I__8023 (
            .O(N__36758),
            .I(N__36755));
    Span4Mux_h I__8022 (
            .O(N__36755),
            .I(N__36751));
    InMux I__8021 (
            .O(N__36754),
            .I(N__36748));
    Odrv4 I__8020 (
            .O(N__36751),
            .I(data_in_15_1));
    LocalMux I__8019 (
            .O(N__36748),
            .I(data_in_15_1));
    InMux I__8018 (
            .O(N__36743),
            .I(N__36736));
    InMux I__8017 (
            .O(N__36742),
            .I(N__36736));
    CascadeMux I__8016 (
            .O(N__36741),
            .I(N__36733));
    LocalMux I__8015 (
            .O(N__36736),
            .I(N__36730));
    InMux I__8014 (
            .O(N__36733),
            .I(N__36726));
    Span4Mux_v I__8013 (
            .O(N__36730),
            .I(N__36723));
    InMux I__8012 (
            .O(N__36729),
            .I(N__36720));
    LocalMux I__8011 (
            .O(N__36726),
            .I(N__36717));
    IoSpan4Mux I__8010 (
            .O(N__36723),
            .I(N__36714));
    LocalMux I__8009 (
            .O(N__36720),
            .I(N__36711));
    Span4Mux_h I__8008 (
            .O(N__36717),
            .I(N__36708));
    IoSpan4Mux I__8007 (
            .O(N__36714),
            .I(N__36705));
    Span12Mux_h I__8006 (
            .O(N__36711),
            .I(N__36702));
    Span4Mux_s2_h I__8005 (
            .O(N__36708),
            .I(N__36699));
    Odrv4 I__8004 (
            .O(N__36705),
            .I(\c0.data_in_frame_9_1 ));
    Odrv12 I__8003 (
            .O(N__36702),
            .I(\c0.data_in_frame_9_1 ));
    Odrv4 I__8002 (
            .O(N__36699),
            .I(\c0.data_in_frame_9_1 ));
    InMux I__8001 (
            .O(N__36692),
            .I(N__36687));
    InMux I__8000 (
            .O(N__36691),
            .I(N__36682));
    InMux I__7999 (
            .O(N__36690),
            .I(N__36679));
    LocalMux I__7998 (
            .O(N__36687),
            .I(N__36676));
    InMux I__7997 (
            .O(N__36686),
            .I(N__36673));
    CascadeMux I__7996 (
            .O(N__36685),
            .I(N__36670));
    LocalMux I__7995 (
            .O(N__36682),
            .I(N__36667));
    LocalMux I__7994 (
            .O(N__36679),
            .I(N__36664));
    Span4Mux_h I__7993 (
            .O(N__36676),
            .I(N__36659));
    LocalMux I__7992 (
            .O(N__36673),
            .I(N__36659));
    InMux I__7991 (
            .O(N__36670),
            .I(N__36656));
    Span4Mux_v I__7990 (
            .O(N__36667),
            .I(N__36653));
    Span4Mux_v I__7989 (
            .O(N__36664),
            .I(N__36650));
    Span4Mux_v I__7988 (
            .O(N__36659),
            .I(N__36645));
    LocalMux I__7987 (
            .O(N__36656),
            .I(N__36645));
    Span4Mux_h I__7986 (
            .O(N__36653),
            .I(N__36642));
    Span4Mux_h I__7985 (
            .O(N__36650),
            .I(N__36637));
    Span4Mux_v I__7984 (
            .O(N__36645),
            .I(N__36637));
    Odrv4 I__7983 (
            .O(N__36642),
            .I(\c0.data_in_frame_10_7 ));
    Odrv4 I__7982 (
            .O(N__36637),
            .I(\c0.data_in_frame_10_7 ));
    InMux I__7981 (
            .O(N__36632),
            .I(N__36626));
    InMux I__7980 (
            .O(N__36631),
            .I(N__36626));
    LocalMux I__7979 (
            .O(N__36626),
            .I(N__36621));
    CascadeMux I__7978 (
            .O(N__36625),
            .I(N__36618));
    CascadeMux I__7977 (
            .O(N__36624),
            .I(N__36615));
    Span4Mux_h I__7976 (
            .O(N__36621),
            .I(N__36612));
    InMux I__7975 (
            .O(N__36618),
            .I(N__36609));
    InMux I__7974 (
            .O(N__36615),
            .I(N__36606));
    Span4Mux_v I__7973 (
            .O(N__36612),
            .I(N__36601));
    LocalMux I__7972 (
            .O(N__36609),
            .I(N__36601));
    LocalMux I__7971 (
            .O(N__36606),
            .I(N__36598));
    Span4Mux_v I__7970 (
            .O(N__36601),
            .I(N__36594));
    Span4Mux_h I__7969 (
            .O(N__36598),
            .I(N__36591));
    InMux I__7968 (
            .O(N__36597),
            .I(N__36588));
    Odrv4 I__7967 (
            .O(N__36594),
            .I(\c0.data_in_frame_9_5 ));
    Odrv4 I__7966 (
            .O(N__36591),
            .I(\c0.data_in_frame_9_5 ));
    LocalMux I__7965 (
            .O(N__36588),
            .I(\c0.data_in_frame_9_5 ));
    CascadeMux I__7964 (
            .O(N__36581),
            .I(N__36576));
    InMux I__7963 (
            .O(N__36580),
            .I(N__36573));
    InMux I__7962 (
            .O(N__36579),
            .I(N__36568));
    InMux I__7961 (
            .O(N__36576),
            .I(N__36568));
    LocalMux I__7960 (
            .O(N__36573),
            .I(N__36565));
    LocalMux I__7959 (
            .O(N__36568),
            .I(N__36562));
    Odrv12 I__7958 (
            .O(N__36565),
            .I(\c0.data_in_frame_9_3 ));
    Odrv4 I__7957 (
            .O(N__36562),
            .I(\c0.data_in_frame_9_3 ));
    CascadeMux I__7956 (
            .O(N__36557),
            .I(N__36553));
    InMux I__7955 (
            .O(N__36556),
            .I(N__36548));
    InMux I__7954 (
            .O(N__36553),
            .I(N__36548));
    LocalMux I__7953 (
            .O(N__36548),
            .I(N__36544));
    InMux I__7952 (
            .O(N__36547),
            .I(N__36541));
    Span4Mux_v I__7951 (
            .O(N__36544),
            .I(N__36538));
    LocalMux I__7950 (
            .O(N__36541),
            .I(N__36535));
    Span4Mux_h I__7949 (
            .O(N__36538),
            .I(N__36532));
    Span12Mux_s9_h I__7948 (
            .O(N__36535),
            .I(N__36529));
    Odrv4 I__7947 (
            .O(N__36532),
            .I(\c0.n8989 ));
    Odrv12 I__7946 (
            .O(N__36529),
            .I(\c0.n8989 ));
    InMux I__7945 (
            .O(N__36524),
            .I(N__36520));
    InMux I__7944 (
            .O(N__36523),
            .I(N__36517));
    LocalMux I__7943 (
            .O(N__36520),
            .I(N__36513));
    LocalMux I__7942 (
            .O(N__36517),
            .I(N__36510));
    InMux I__7941 (
            .O(N__36516),
            .I(N__36507));
    Span4Mux_v I__7940 (
            .O(N__36513),
            .I(N__36504));
    Odrv4 I__7939 (
            .O(N__36510),
            .I(data_in_10_2));
    LocalMux I__7938 (
            .O(N__36507),
            .I(data_in_10_2));
    Odrv4 I__7937 (
            .O(N__36504),
            .I(data_in_10_2));
    InMux I__7936 (
            .O(N__36497),
            .I(N__36494));
    LocalMux I__7935 (
            .O(N__36494),
            .I(N__36489));
    InMux I__7934 (
            .O(N__36493),
            .I(N__36486));
    InMux I__7933 (
            .O(N__36492),
            .I(N__36483));
    Span4Mux_v I__7932 (
            .O(N__36489),
            .I(N__36480));
    LocalMux I__7931 (
            .O(N__36486),
            .I(N__36477));
    LocalMux I__7930 (
            .O(N__36483),
            .I(data_in_9_2));
    Odrv4 I__7929 (
            .O(N__36480),
            .I(data_in_9_2));
    Odrv4 I__7928 (
            .O(N__36477),
            .I(data_in_9_2));
    CascadeMux I__7927 (
            .O(N__36470),
            .I(N__36467));
    InMux I__7926 (
            .O(N__36467),
            .I(N__36464));
    LocalMux I__7925 (
            .O(N__36464),
            .I(N__36460));
    InMux I__7924 (
            .O(N__36463),
            .I(N__36455));
    Span4Mux_v I__7923 (
            .O(N__36460),
            .I(N__36452));
    InMux I__7922 (
            .O(N__36459),
            .I(N__36449));
    InMux I__7921 (
            .O(N__36458),
            .I(N__36446));
    LocalMux I__7920 (
            .O(N__36455),
            .I(N__36443));
    Span4Mux_v I__7919 (
            .O(N__36452),
            .I(N__36438));
    LocalMux I__7918 (
            .O(N__36449),
            .I(N__36438));
    LocalMux I__7917 (
            .O(N__36446),
            .I(N__36434));
    Span12Mux_s4_h I__7916 (
            .O(N__36443),
            .I(N__36431));
    Span4Mux_h I__7915 (
            .O(N__36438),
            .I(N__36428));
    InMux I__7914 (
            .O(N__36437),
            .I(N__36425));
    Span4Mux_h I__7913 (
            .O(N__36434),
            .I(N__36422));
    Odrv12 I__7912 (
            .O(N__36431),
            .I(rand_data_28));
    Odrv4 I__7911 (
            .O(N__36428),
            .I(rand_data_28));
    LocalMux I__7910 (
            .O(N__36425),
            .I(rand_data_28));
    Odrv4 I__7909 (
            .O(N__36422),
            .I(rand_data_28));
    InMux I__7908 (
            .O(N__36413),
            .I(n16439));
    InMux I__7907 (
            .O(N__36410),
            .I(N__36403));
    InMux I__7906 (
            .O(N__36409),
            .I(N__36403));
    InMux I__7905 (
            .O(N__36408),
            .I(N__36400));
    LocalMux I__7904 (
            .O(N__36403),
            .I(N__36396));
    LocalMux I__7903 (
            .O(N__36400),
            .I(N__36393));
    CascadeMux I__7902 (
            .O(N__36399),
            .I(N__36390));
    Span4Mux_v I__7901 (
            .O(N__36396),
            .I(N__36387));
    Span4Mux_v I__7900 (
            .O(N__36393),
            .I(N__36384));
    InMux I__7899 (
            .O(N__36390),
            .I(N__36380));
    Span4Mux_h I__7898 (
            .O(N__36387),
            .I(N__36377));
    Span4Mux_v I__7897 (
            .O(N__36384),
            .I(N__36374));
    InMux I__7896 (
            .O(N__36383),
            .I(N__36371));
    LocalMux I__7895 (
            .O(N__36380),
            .I(N__36368));
    Odrv4 I__7894 (
            .O(N__36377),
            .I(rand_data_29));
    Odrv4 I__7893 (
            .O(N__36374),
            .I(rand_data_29));
    LocalMux I__7892 (
            .O(N__36371),
            .I(rand_data_29));
    Odrv12 I__7891 (
            .O(N__36368),
            .I(rand_data_29));
    InMux I__7890 (
            .O(N__36359),
            .I(n16440));
    InMux I__7889 (
            .O(N__36356),
            .I(N__36348));
    InMux I__7888 (
            .O(N__36355),
            .I(N__36348));
    InMux I__7887 (
            .O(N__36354),
            .I(N__36345));
    CascadeMux I__7886 (
            .O(N__36353),
            .I(N__36342));
    LocalMux I__7885 (
            .O(N__36348),
            .I(N__36339));
    LocalMux I__7884 (
            .O(N__36345),
            .I(N__36336));
    InMux I__7883 (
            .O(N__36342),
            .I(N__36332));
    Span4Mux_v I__7882 (
            .O(N__36339),
            .I(N__36329));
    Span12Mux_h I__7881 (
            .O(N__36336),
            .I(N__36326));
    InMux I__7880 (
            .O(N__36335),
            .I(N__36323));
    LocalMux I__7879 (
            .O(N__36332),
            .I(N__36320));
    Odrv4 I__7878 (
            .O(N__36329),
            .I(rand_data_30));
    Odrv12 I__7877 (
            .O(N__36326),
            .I(rand_data_30));
    LocalMux I__7876 (
            .O(N__36323),
            .I(rand_data_30));
    Odrv12 I__7875 (
            .O(N__36320),
            .I(rand_data_30));
    InMux I__7874 (
            .O(N__36311),
            .I(n16441));
    InMux I__7873 (
            .O(N__36308),
            .I(N__36301));
    InMux I__7872 (
            .O(N__36307),
            .I(N__36301));
    InMux I__7871 (
            .O(N__36306),
            .I(N__36298));
    LocalMux I__7870 (
            .O(N__36301),
            .I(N__36294));
    LocalMux I__7869 (
            .O(N__36298),
            .I(N__36291));
    InMux I__7868 (
            .O(N__36297),
            .I(N__36288));
    Span4Mux_v I__7867 (
            .O(N__36294),
            .I(N__36284));
    Span4Mux_h I__7866 (
            .O(N__36291),
            .I(N__36281));
    LocalMux I__7865 (
            .O(N__36288),
            .I(N__36278));
    InMux I__7864 (
            .O(N__36287),
            .I(N__36275));
    Span4Mux_v I__7863 (
            .O(N__36284),
            .I(N__36268));
    Span4Mux_v I__7862 (
            .O(N__36281),
            .I(N__36268));
    Span4Mux_h I__7861 (
            .O(N__36278),
            .I(N__36268));
    LocalMux I__7860 (
            .O(N__36275),
            .I(rand_data_31));
    Odrv4 I__7859 (
            .O(N__36268),
            .I(rand_data_31));
    InMux I__7858 (
            .O(N__36263),
            .I(n16442));
    InMux I__7857 (
            .O(N__36260),
            .I(N__36256));
    InMux I__7856 (
            .O(N__36259),
            .I(N__36253));
    LocalMux I__7855 (
            .O(N__36256),
            .I(N__36250));
    LocalMux I__7854 (
            .O(N__36253),
            .I(N__36247));
    Span4Mux_h I__7853 (
            .O(N__36250),
            .I(N__36244));
    Span4Mux_h I__7852 (
            .O(N__36247),
            .I(N__36239));
    Span4Mux_h I__7851 (
            .O(N__36244),
            .I(N__36236));
    InMux I__7850 (
            .O(N__36243),
            .I(N__36231));
    InMux I__7849 (
            .O(N__36242),
            .I(N__36231));
    Odrv4 I__7848 (
            .O(N__36239),
            .I(data_in_1_5));
    Odrv4 I__7847 (
            .O(N__36236),
            .I(data_in_1_5));
    LocalMux I__7846 (
            .O(N__36231),
            .I(data_in_1_5));
    InMux I__7845 (
            .O(N__36224),
            .I(N__36220));
    CascadeMux I__7844 (
            .O(N__36223),
            .I(N__36217));
    LocalMux I__7843 (
            .O(N__36220),
            .I(N__36214));
    InMux I__7842 (
            .O(N__36217),
            .I(N__36211));
    Span4Mux_v I__7841 (
            .O(N__36214),
            .I(N__36207));
    LocalMux I__7840 (
            .O(N__36211),
            .I(N__36204));
    InMux I__7839 (
            .O(N__36210),
            .I(N__36201));
    Span4Mux_h I__7838 (
            .O(N__36207),
            .I(N__36196));
    Span4Mux_v I__7837 (
            .O(N__36204),
            .I(N__36196));
    LocalMux I__7836 (
            .O(N__36201),
            .I(data_in_7_5));
    Odrv4 I__7835 (
            .O(N__36196),
            .I(data_in_7_5));
    InMux I__7834 (
            .O(N__36191),
            .I(N__36187));
    CascadeMux I__7833 (
            .O(N__36190),
            .I(N__36184));
    LocalMux I__7832 (
            .O(N__36187),
            .I(N__36181));
    InMux I__7831 (
            .O(N__36184),
            .I(N__36178));
    Span4Mux_v I__7830 (
            .O(N__36181),
            .I(N__36174));
    LocalMux I__7829 (
            .O(N__36178),
            .I(N__36171));
    InMux I__7828 (
            .O(N__36177),
            .I(N__36168));
    Span4Mux_h I__7827 (
            .O(N__36174),
            .I(N__36165));
    Span4Mux_h I__7826 (
            .O(N__36171),
            .I(N__36162));
    LocalMux I__7825 (
            .O(N__36168),
            .I(data_in_6_5));
    Odrv4 I__7824 (
            .O(N__36165),
            .I(data_in_6_5));
    Odrv4 I__7823 (
            .O(N__36162),
            .I(data_in_6_5));
    InMux I__7822 (
            .O(N__36155),
            .I(N__36152));
    LocalMux I__7821 (
            .O(N__36152),
            .I(N__36148));
    InMux I__7820 (
            .O(N__36151),
            .I(N__36145));
    Span4Mux_s2_h I__7819 (
            .O(N__36148),
            .I(N__36138));
    LocalMux I__7818 (
            .O(N__36145),
            .I(N__36138));
    InMux I__7817 (
            .O(N__36144),
            .I(N__36135));
    InMux I__7816 (
            .O(N__36143),
            .I(N__36132));
    Span4Mux_v I__7815 (
            .O(N__36138),
            .I(N__36128));
    LocalMux I__7814 (
            .O(N__36135),
            .I(N__36125));
    LocalMux I__7813 (
            .O(N__36132),
            .I(N__36122));
    InMux I__7812 (
            .O(N__36131),
            .I(N__36119));
    Span4Mux_s1_v I__7811 (
            .O(N__36128),
            .I(N__36114));
    Span4Mux_h I__7810 (
            .O(N__36125),
            .I(N__36114));
    Odrv4 I__7809 (
            .O(N__36122),
            .I(rand_data_20));
    LocalMux I__7808 (
            .O(N__36119),
            .I(rand_data_20));
    Odrv4 I__7807 (
            .O(N__36114),
            .I(rand_data_20));
    InMux I__7806 (
            .O(N__36107),
            .I(n16431));
    InMux I__7805 (
            .O(N__36104),
            .I(N__36101));
    LocalMux I__7804 (
            .O(N__36101),
            .I(N__36095));
    InMux I__7803 (
            .O(N__36100),
            .I(N__36092));
    InMux I__7802 (
            .O(N__36099),
            .I(N__36089));
    CascadeMux I__7801 (
            .O(N__36098),
            .I(N__36086));
    Span4Mux_h I__7800 (
            .O(N__36095),
            .I(N__36083));
    LocalMux I__7799 (
            .O(N__36092),
            .I(N__36080));
    LocalMux I__7798 (
            .O(N__36089),
            .I(N__36077));
    InMux I__7797 (
            .O(N__36086),
            .I(N__36073));
    Span4Mux_v I__7796 (
            .O(N__36083),
            .I(N__36070));
    Span4Mux_h I__7795 (
            .O(N__36080),
            .I(N__36067));
    Span4Mux_v I__7794 (
            .O(N__36077),
            .I(N__36064));
    InMux I__7793 (
            .O(N__36076),
            .I(N__36061));
    LocalMux I__7792 (
            .O(N__36073),
            .I(N__36058));
    Odrv4 I__7791 (
            .O(N__36070),
            .I(rand_data_21));
    Odrv4 I__7790 (
            .O(N__36067),
            .I(rand_data_21));
    Odrv4 I__7789 (
            .O(N__36064),
            .I(rand_data_21));
    LocalMux I__7788 (
            .O(N__36061),
            .I(rand_data_21));
    Odrv12 I__7787 (
            .O(N__36058),
            .I(rand_data_21));
    InMux I__7786 (
            .O(N__36047),
            .I(n16432));
    InMux I__7785 (
            .O(N__36044),
            .I(N__36035));
    InMux I__7784 (
            .O(N__36043),
            .I(N__36035));
    InMux I__7783 (
            .O(N__36042),
            .I(N__36035));
    LocalMux I__7782 (
            .O(N__36035),
            .I(N__36031));
    CascadeMux I__7781 (
            .O(N__36034),
            .I(N__36028));
    Sp12to4 I__7780 (
            .O(N__36031),
            .I(N__36024));
    InMux I__7779 (
            .O(N__36028),
            .I(N__36021));
    InMux I__7778 (
            .O(N__36027),
            .I(N__36018));
    Span12Mux_v I__7777 (
            .O(N__36024),
            .I(N__36013));
    LocalMux I__7776 (
            .O(N__36021),
            .I(N__36013));
    LocalMux I__7775 (
            .O(N__36018),
            .I(rand_data_22));
    Odrv12 I__7774 (
            .O(N__36013),
            .I(rand_data_22));
    InMux I__7773 (
            .O(N__36008),
            .I(n16433));
    InMux I__7772 (
            .O(N__36005),
            .I(N__36000));
    InMux I__7771 (
            .O(N__36004),
            .I(N__35995));
    InMux I__7770 (
            .O(N__36003),
            .I(N__35995));
    LocalMux I__7769 (
            .O(N__36000),
            .I(N__35992));
    LocalMux I__7768 (
            .O(N__35995),
            .I(N__35988));
    Span4Mux_h I__7767 (
            .O(N__35992),
            .I(N__35985));
    InMux I__7766 (
            .O(N__35991),
            .I(N__35982));
    Span4Mux_h I__7765 (
            .O(N__35988),
            .I(N__35979));
    Span4Mux_v I__7764 (
            .O(N__35985),
            .I(N__35975));
    LocalMux I__7763 (
            .O(N__35982),
            .I(N__35972));
    Span4Mux_v I__7762 (
            .O(N__35979),
            .I(N__35969));
    InMux I__7761 (
            .O(N__35978),
            .I(N__35966));
    Span4Mux_s1_h I__7760 (
            .O(N__35975),
            .I(N__35961));
    Span4Mux_h I__7759 (
            .O(N__35972),
            .I(N__35961));
    Odrv4 I__7758 (
            .O(N__35969),
            .I(rand_data_23));
    LocalMux I__7757 (
            .O(N__35966),
            .I(rand_data_23));
    Odrv4 I__7756 (
            .O(N__35961),
            .I(rand_data_23));
    InMux I__7755 (
            .O(N__35954),
            .I(n16434));
    InMux I__7754 (
            .O(N__35951),
            .I(N__35946));
    InMux I__7753 (
            .O(N__35950),
            .I(N__35943));
    InMux I__7752 (
            .O(N__35949),
            .I(N__35940));
    LocalMux I__7751 (
            .O(N__35946),
            .I(N__35936));
    LocalMux I__7750 (
            .O(N__35943),
            .I(N__35933));
    LocalMux I__7749 (
            .O(N__35940),
            .I(N__35930));
    InMux I__7748 (
            .O(N__35939),
            .I(N__35927));
    Span4Mux_v I__7747 (
            .O(N__35936),
            .I(N__35924));
    Span4Mux_h I__7746 (
            .O(N__35933),
            .I(N__35921));
    Span4Mux_h I__7745 (
            .O(N__35930),
            .I(N__35917));
    LocalMux I__7744 (
            .O(N__35927),
            .I(N__35914));
    Span4Mux_v I__7743 (
            .O(N__35924),
            .I(N__35911));
    Span4Mux_v I__7742 (
            .O(N__35921),
            .I(N__35908));
    InMux I__7741 (
            .O(N__35920),
            .I(N__35905));
    Span4Mux_v I__7740 (
            .O(N__35917),
            .I(N__35900));
    Span4Mux_h I__7739 (
            .O(N__35914),
            .I(N__35900));
    Odrv4 I__7738 (
            .O(N__35911),
            .I(rand_data_24));
    Odrv4 I__7737 (
            .O(N__35908),
            .I(rand_data_24));
    LocalMux I__7736 (
            .O(N__35905),
            .I(rand_data_24));
    Odrv4 I__7735 (
            .O(N__35900),
            .I(rand_data_24));
    InMux I__7734 (
            .O(N__35891),
            .I(bfn_9_32_0_));
    InMux I__7733 (
            .O(N__35888),
            .I(N__35883));
    InMux I__7732 (
            .O(N__35887),
            .I(N__35880));
    InMux I__7731 (
            .O(N__35886),
            .I(N__35877));
    LocalMux I__7730 (
            .O(N__35883),
            .I(N__35874));
    LocalMux I__7729 (
            .O(N__35880),
            .I(N__35871));
    LocalMux I__7728 (
            .O(N__35877),
            .I(N__35868));
    Span4Mux_h I__7727 (
            .O(N__35874),
            .I(N__35864));
    Span4Mux_h I__7726 (
            .O(N__35871),
            .I(N__35861));
    Span4Mux_v I__7725 (
            .O(N__35868),
            .I(N__35857));
    InMux I__7724 (
            .O(N__35867),
            .I(N__35854));
    Span4Mux_v I__7723 (
            .O(N__35864),
            .I(N__35851));
    Span4Mux_v I__7722 (
            .O(N__35861),
            .I(N__35848));
    InMux I__7721 (
            .O(N__35860),
            .I(N__35845));
    Sp12to4 I__7720 (
            .O(N__35857),
            .I(N__35840));
    LocalMux I__7719 (
            .O(N__35854),
            .I(N__35840));
    Odrv4 I__7718 (
            .O(N__35851),
            .I(rand_data_25));
    Odrv4 I__7717 (
            .O(N__35848),
            .I(rand_data_25));
    LocalMux I__7716 (
            .O(N__35845),
            .I(rand_data_25));
    Odrv12 I__7715 (
            .O(N__35840),
            .I(rand_data_25));
    InMux I__7714 (
            .O(N__35831),
            .I(n16436));
    InMux I__7713 (
            .O(N__35828),
            .I(N__35825));
    LocalMux I__7712 (
            .O(N__35825),
            .I(N__35822));
    Span4Mux_v I__7711 (
            .O(N__35822),
            .I(N__35818));
    InMux I__7710 (
            .O(N__35821),
            .I(N__35815));
    Span4Mux_s1_h I__7709 (
            .O(N__35818),
            .I(N__35810));
    LocalMux I__7708 (
            .O(N__35815),
            .I(N__35810));
    Span4Mux_v I__7707 (
            .O(N__35810),
            .I(N__35806));
    InMux I__7706 (
            .O(N__35809),
            .I(N__35803));
    Span4Mux_s1_h I__7705 (
            .O(N__35806),
            .I(N__35797));
    LocalMux I__7704 (
            .O(N__35803),
            .I(N__35797));
    InMux I__7703 (
            .O(N__35802),
            .I(N__35793));
    Span4Mux_h I__7702 (
            .O(N__35797),
            .I(N__35790));
    InMux I__7701 (
            .O(N__35796),
            .I(N__35787));
    LocalMux I__7700 (
            .O(N__35793),
            .I(N__35784));
    Odrv4 I__7699 (
            .O(N__35790),
            .I(rand_data_26));
    LocalMux I__7698 (
            .O(N__35787),
            .I(rand_data_26));
    Odrv12 I__7697 (
            .O(N__35784),
            .I(rand_data_26));
    InMux I__7696 (
            .O(N__35777),
            .I(n16437));
    InMux I__7695 (
            .O(N__35774),
            .I(N__35771));
    LocalMux I__7694 (
            .O(N__35771),
            .I(N__35766));
    InMux I__7693 (
            .O(N__35770),
            .I(N__35763));
    InMux I__7692 (
            .O(N__35769),
            .I(N__35760));
    Span4Mux_v I__7691 (
            .O(N__35766),
            .I(N__35756));
    LocalMux I__7690 (
            .O(N__35763),
            .I(N__35753));
    LocalMux I__7689 (
            .O(N__35760),
            .I(N__35750));
    InMux I__7688 (
            .O(N__35759),
            .I(N__35746));
    Span4Mux_v I__7687 (
            .O(N__35756),
            .I(N__35743));
    Span4Mux_h I__7686 (
            .O(N__35753),
            .I(N__35740));
    Span4Mux_h I__7685 (
            .O(N__35750),
            .I(N__35737));
    InMux I__7684 (
            .O(N__35749),
            .I(N__35734));
    LocalMux I__7683 (
            .O(N__35746),
            .I(N__35731));
    Odrv4 I__7682 (
            .O(N__35743),
            .I(rand_data_27));
    Odrv4 I__7681 (
            .O(N__35740),
            .I(rand_data_27));
    Odrv4 I__7680 (
            .O(N__35737),
            .I(rand_data_27));
    LocalMux I__7679 (
            .O(N__35734),
            .I(rand_data_27));
    Odrv12 I__7678 (
            .O(N__35731),
            .I(rand_data_27));
    InMux I__7677 (
            .O(N__35720),
            .I(n16438));
    InMux I__7676 (
            .O(N__35717),
            .I(N__35710));
    InMux I__7675 (
            .O(N__35716),
            .I(N__35710));
    InMux I__7674 (
            .O(N__35715),
            .I(N__35707));
    LocalMux I__7673 (
            .O(N__35710),
            .I(N__35701));
    LocalMux I__7672 (
            .O(N__35707),
            .I(N__35701));
    InMux I__7671 (
            .O(N__35706),
            .I(N__35698));
    Span4Mux_h I__7670 (
            .O(N__35701),
            .I(N__35693));
    LocalMux I__7669 (
            .O(N__35698),
            .I(N__35693));
    Span4Mux_v I__7668 (
            .O(N__35693),
            .I(N__35690));
    Span4Mux_s1_h I__7667 (
            .O(N__35690),
            .I(N__35686));
    InMux I__7666 (
            .O(N__35689),
            .I(N__35682));
    Span4Mux_h I__7665 (
            .O(N__35686),
            .I(N__35679));
    InMux I__7664 (
            .O(N__35685),
            .I(N__35676));
    LocalMux I__7663 (
            .O(N__35682),
            .I(N__35673));
    Odrv4 I__7662 (
            .O(N__35679),
            .I(rand_data_11));
    LocalMux I__7661 (
            .O(N__35676),
            .I(rand_data_11));
    Odrv12 I__7660 (
            .O(N__35673),
            .I(rand_data_11));
    InMux I__7659 (
            .O(N__35666),
            .I(n16422));
    CascadeMux I__7658 (
            .O(N__35663),
            .I(N__35659));
    InMux I__7657 (
            .O(N__35662),
            .I(N__35654));
    InMux I__7656 (
            .O(N__35659),
            .I(N__35651));
    InMux I__7655 (
            .O(N__35658),
            .I(N__35648));
    InMux I__7654 (
            .O(N__35657),
            .I(N__35644));
    LocalMux I__7653 (
            .O(N__35654),
            .I(N__35641));
    LocalMux I__7652 (
            .O(N__35651),
            .I(N__35636));
    LocalMux I__7651 (
            .O(N__35648),
            .I(N__35636));
    InMux I__7650 (
            .O(N__35647),
            .I(N__35633));
    LocalMux I__7649 (
            .O(N__35644),
            .I(N__35629));
    Span4Mux_v I__7648 (
            .O(N__35641),
            .I(N__35626));
    Span4Mux_h I__7647 (
            .O(N__35636),
            .I(N__35621));
    LocalMux I__7646 (
            .O(N__35633),
            .I(N__35621));
    InMux I__7645 (
            .O(N__35632),
            .I(N__35618));
    Span4Mux_h I__7644 (
            .O(N__35629),
            .I(N__35615));
    Odrv4 I__7643 (
            .O(N__35626),
            .I(rand_data_12));
    Odrv4 I__7642 (
            .O(N__35621),
            .I(rand_data_12));
    LocalMux I__7641 (
            .O(N__35618),
            .I(rand_data_12));
    Odrv4 I__7640 (
            .O(N__35615),
            .I(rand_data_12));
    InMux I__7639 (
            .O(N__35606),
            .I(n16423));
    InMux I__7638 (
            .O(N__35603),
            .I(N__35596));
    InMux I__7637 (
            .O(N__35602),
            .I(N__35596));
    InMux I__7636 (
            .O(N__35601),
            .I(N__35592));
    LocalMux I__7635 (
            .O(N__35596),
            .I(N__35589));
    InMux I__7634 (
            .O(N__35595),
            .I(N__35586));
    LocalMux I__7633 (
            .O(N__35592),
            .I(N__35582));
    Span4Mux_v I__7632 (
            .O(N__35589),
            .I(N__35579));
    LocalMux I__7631 (
            .O(N__35586),
            .I(N__35576));
    InMux I__7630 (
            .O(N__35585),
            .I(N__35573));
    Span4Mux_h I__7629 (
            .O(N__35582),
            .I(N__35570));
    Span4Mux_v I__7628 (
            .O(N__35579),
            .I(N__35567));
    Span4Mux_s1_h I__7627 (
            .O(N__35576),
            .I(N__35564));
    LocalMux I__7626 (
            .O(N__35573),
            .I(N__35560));
    Span4Mux_v I__7625 (
            .O(N__35570),
            .I(N__35557));
    Span4Mux_s1_h I__7624 (
            .O(N__35567),
            .I(N__35552));
    Span4Mux_v I__7623 (
            .O(N__35564),
            .I(N__35552));
    InMux I__7622 (
            .O(N__35563),
            .I(N__35549));
    Span4Mux_h I__7621 (
            .O(N__35560),
            .I(N__35546));
    Odrv4 I__7620 (
            .O(N__35557),
            .I(rand_data_13));
    Odrv4 I__7619 (
            .O(N__35552),
            .I(rand_data_13));
    LocalMux I__7618 (
            .O(N__35549),
            .I(rand_data_13));
    Odrv4 I__7617 (
            .O(N__35546),
            .I(rand_data_13));
    InMux I__7616 (
            .O(N__35537),
            .I(n16424));
    InMux I__7615 (
            .O(N__35534),
            .I(N__35529));
    InMux I__7614 (
            .O(N__35533),
            .I(N__35524));
    InMux I__7613 (
            .O(N__35532),
            .I(N__35524));
    LocalMux I__7612 (
            .O(N__35529),
            .I(N__35519));
    LocalMux I__7611 (
            .O(N__35524),
            .I(N__35516));
    InMux I__7610 (
            .O(N__35523),
            .I(N__35513));
    CascadeMux I__7609 (
            .O(N__35522),
            .I(N__35510));
    Span4Mux_v I__7608 (
            .O(N__35519),
            .I(N__35507));
    Span4Mux_h I__7607 (
            .O(N__35516),
            .I(N__35504));
    LocalMux I__7606 (
            .O(N__35513),
            .I(N__35500));
    InMux I__7605 (
            .O(N__35510),
            .I(N__35497));
    Span4Mux_v I__7604 (
            .O(N__35507),
            .I(N__35492));
    Span4Mux_v I__7603 (
            .O(N__35504),
            .I(N__35492));
    InMux I__7602 (
            .O(N__35503),
            .I(N__35489));
    Span12Mux_v I__7601 (
            .O(N__35500),
            .I(N__35484));
    LocalMux I__7600 (
            .O(N__35497),
            .I(N__35484));
    Odrv4 I__7599 (
            .O(N__35492),
            .I(rand_data_14));
    LocalMux I__7598 (
            .O(N__35489),
            .I(rand_data_14));
    Odrv12 I__7597 (
            .O(N__35484),
            .I(rand_data_14));
    InMux I__7596 (
            .O(N__35477),
            .I(n16425));
    InMux I__7595 (
            .O(N__35474),
            .I(N__35471));
    LocalMux I__7594 (
            .O(N__35471),
            .I(N__35468));
    Span4Mux_h I__7593 (
            .O(N__35468),
            .I(N__35464));
    InMux I__7592 (
            .O(N__35467),
            .I(N__35461));
    Span4Mux_v I__7591 (
            .O(N__35464),
            .I(N__35455));
    LocalMux I__7590 (
            .O(N__35461),
            .I(N__35452));
    InMux I__7589 (
            .O(N__35460),
            .I(N__35449));
    InMux I__7588 (
            .O(N__35459),
            .I(N__35446));
    InMux I__7587 (
            .O(N__35458),
            .I(N__35443));
    Span4Mux_h I__7586 (
            .O(N__35455),
            .I(N__35438));
    Span4Mux_h I__7585 (
            .O(N__35452),
            .I(N__35438));
    LocalMux I__7584 (
            .O(N__35449),
            .I(N__35432));
    LocalMux I__7583 (
            .O(N__35446),
            .I(N__35432));
    LocalMux I__7582 (
            .O(N__35443),
            .I(N__35429));
    Span4Mux_v I__7581 (
            .O(N__35438),
            .I(N__35426));
    InMux I__7580 (
            .O(N__35437),
            .I(N__35423));
    Span4Mux_v I__7579 (
            .O(N__35432),
            .I(N__35418));
    Span4Mux_h I__7578 (
            .O(N__35429),
            .I(N__35418));
    Odrv4 I__7577 (
            .O(N__35426),
            .I(rand_data_15));
    LocalMux I__7576 (
            .O(N__35423),
            .I(rand_data_15));
    Odrv4 I__7575 (
            .O(N__35418),
            .I(rand_data_15));
    InMux I__7574 (
            .O(N__35411),
            .I(n16426));
    InMux I__7573 (
            .O(N__35408),
            .I(N__35403));
    InMux I__7572 (
            .O(N__35407),
            .I(N__35400));
    InMux I__7571 (
            .O(N__35406),
            .I(N__35397));
    LocalMux I__7570 (
            .O(N__35403),
            .I(N__35393));
    LocalMux I__7569 (
            .O(N__35400),
            .I(N__35390));
    LocalMux I__7568 (
            .O(N__35397),
            .I(N__35387));
    InMux I__7567 (
            .O(N__35396),
            .I(N__35383));
    Span4Mux_h I__7566 (
            .O(N__35393),
            .I(N__35380));
    Span4Mux_h I__7565 (
            .O(N__35390),
            .I(N__35375));
    Span4Mux_v I__7564 (
            .O(N__35387),
            .I(N__35375));
    InMux I__7563 (
            .O(N__35386),
            .I(N__35372));
    LocalMux I__7562 (
            .O(N__35383),
            .I(N__35369));
    Odrv4 I__7561 (
            .O(N__35380),
            .I(rand_data_16));
    Odrv4 I__7560 (
            .O(N__35375),
            .I(rand_data_16));
    LocalMux I__7559 (
            .O(N__35372),
            .I(rand_data_16));
    Odrv12 I__7558 (
            .O(N__35369),
            .I(rand_data_16));
    InMux I__7557 (
            .O(N__35360),
            .I(bfn_9_31_0_));
    InMux I__7556 (
            .O(N__35357),
            .I(N__35352));
    InMux I__7555 (
            .O(N__35356),
            .I(N__35349));
    InMux I__7554 (
            .O(N__35355),
            .I(N__35346));
    LocalMux I__7553 (
            .O(N__35352),
            .I(N__35342));
    LocalMux I__7552 (
            .O(N__35349),
            .I(N__35339));
    LocalMux I__7551 (
            .O(N__35346),
            .I(N__35336));
    InMux I__7550 (
            .O(N__35345),
            .I(N__35332));
    Span4Mux_v I__7549 (
            .O(N__35342),
            .I(N__35329));
    Span4Mux_v I__7548 (
            .O(N__35339),
            .I(N__35324));
    Span4Mux_h I__7547 (
            .O(N__35336),
            .I(N__35324));
    InMux I__7546 (
            .O(N__35335),
            .I(N__35321));
    LocalMux I__7545 (
            .O(N__35332),
            .I(N__35318));
    Odrv4 I__7544 (
            .O(N__35329),
            .I(rand_data_17));
    Odrv4 I__7543 (
            .O(N__35324),
            .I(rand_data_17));
    LocalMux I__7542 (
            .O(N__35321),
            .I(rand_data_17));
    Odrv12 I__7541 (
            .O(N__35318),
            .I(rand_data_17));
    InMux I__7540 (
            .O(N__35309),
            .I(n16428));
    InMux I__7539 (
            .O(N__35306),
            .I(N__35302));
    InMux I__7538 (
            .O(N__35305),
            .I(N__35299));
    LocalMux I__7537 (
            .O(N__35302),
            .I(N__35293));
    LocalMux I__7536 (
            .O(N__35299),
            .I(N__35293));
    InMux I__7535 (
            .O(N__35298),
            .I(N__35290));
    Span4Mux_v I__7534 (
            .O(N__35293),
            .I(N__35284));
    LocalMux I__7533 (
            .O(N__35290),
            .I(N__35284));
    InMux I__7532 (
            .O(N__35289),
            .I(N__35280));
    Span4Mux_v I__7531 (
            .O(N__35284),
            .I(N__35277));
    InMux I__7530 (
            .O(N__35283),
            .I(N__35274));
    LocalMux I__7529 (
            .O(N__35280),
            .I(N__35271));
    Odrv4 I__7528 (
            .O(N__35277),
            .I(rand_data_18));
    LocalMux I__7527 (
            .O(N__35274),
            .I(rand_data_18));
    Odrv12 I__7526 (
            .O(N__35271),
            .I(rand_data_18));
    InMux I__7525 (
            .O(N__35264),
            .I(n16429));
    InMux I__7524 (
            .O(N__35261),
            .I(N__35257));
    InMux I__7523 (
            .O(N__35260),
            .I(N__35254));
    LocalMux I__7522 (
            .O(N__35257),
            .I(N__35251));
    LocalMux I__7521 (
            .O(N__35254),
            .I(N__35246));
    Span4Mux_v I__7520 (
            .O(N__35251),
            .I(N__35243));
    InMux I__7519 (
            .O(N__35250),
            .I(N__35240));
    InMux I__7518 (
            .O(N__35249),
            .I(N__35236));
    Span4Mux_h I__7517 (
            .O(N__35246),
            .I(N__35233));
    Sp12to4 I__7516 (
            .O(N__35243),
            .I(N__35228));
    LocalMux I__7515 (
            .O(N__35240),
            .I(N__35228));
    InMux I__7514 (
            .O(N__35239),
            .I(N__35225));
    LocalMux I__7513 (
            .O(N__35236),
            .I(N__35222));
    Odrv4 I__7512 (
            .O(N__35233),
            .I(rand_data_19));
    Odrv12 I__7511 (
            .O(N__35228),
            .I(rand_data_19));
    LocalMux I__7510 (
            .O(N__35225),
            .I(rand_data_19));
    Odrv12 I__7509 (
            .O(N__35222),
            .I(rand_data_19));
    InMux I__7508 (
            .O(N__35213),
            .I(n16430));
    InMux I__7507 (
            .O(N__35210),
            .I(N__35206));
    InMux I__7506 (
            .O(N__35209),
            .I(N__35201));
    LocalMux I__7505 (
            .O(N__35206),
            .I(N__35198));
    InMux I__7504 (
            .O(N__35205),
            .I(N__35195));
    InMux I__7503 (
            .O(N__35204),
            .I(N__35191));
    LocalMux I__7502 (
            .O(N__35201),
            .I(N__35187));
    Span4Mux_v I__7501 (
            .O(N__35198),
            .I(N__35184));
    LocalMux I__7500 (
            .O(N__35195),
            .I(N__35181));
    InMux I__7499 (
            .O(N__35194),
            .I(N__35178));
    LocalMux I__7498 (
            .O(N__35191),
            .I(N__35175));
    InMux I__7497 (
            .O(N__35190),
            .I(N__35172));
    Span4Mux_v I__7496 (
            .O(N__35187),
            .I(N__35165));
    Span4Mux_s3_h I__7495 (
            .O(N__35184),
            .I(N__35165));
    Span4Mux_h I__7494 (
            .O(N__35181),
            .I(N__35165));
    LocalMux I__7493 (
            .O(N__35178),
            .I(rand_data_3));
    Odrv4 I__7492 (
            .O(N__35175),
            .I(rand_data_3));
    LocalMux I__7491 (
            .O(N__35172),
            .I(rand_data_3));
    Odrv4 I__7490 (
            .O(N__35165),
            .I(rand_data_3));
    InMux I__7489 (
            .O(N__35156),
            .I(n16414));
    InMux I__7488 (
            .O(N__35153),
            .I(N__35150));
    LocalMux I__7487 (
            .O(N__35150),
            .I(N__35146));
    CascadeMux I__7486 (
            .O(N__35149),
            .I(N__35143));
    Span4Mux_v I__7485 (
            .O(N__35146),
            .I(N__35140));
    InMux I__7484 (
            .O(N__35143),
            .I(N__35134));
    Span4Mux_h I__7483 (
            .O(N__35140),
            .I(N__35130));
    InMux I__7482 (
            .O(N__35139),
            .I(N__35127));
    InMux I__7481 (
            .O(N__35138),
            .I(N__35122));
    InMux I__7480 (
            .O(N__35137),
            .I(N__35122));
    LocalMux I__7479 (
            .O(N__35134),
            .I(N__35119));
    InMux I__7478 (
            .O(N__35133),
            .I(N__35116));
    Sp12to4 I__7477 (
            .O(N__35130),
            .I(N__35111));
    LocalMux I__7476 (
            .O(N__35127),
            .I(N__35111));
    LocalMux I__7475 (
            .O(N__35122),
            .I(rand_data_4));
    Odrv4 I__7474 (
            .O(N__35119),
            .I(rand_data_4));
    LocalMux I__7473 (
            .O(N__35116),
            .I(rand_data_4));
    Odrv12 I__7472 (
            .O(N__35111),
            .I(rand_data_4));
    InMux I__7471 (
            .O(N__35102),
            .I(n16415));
    InMux I__7470 (
            .O(N__35099),
            .I(N__35094));
    InMux I__7469 (
            .O(N__35098),
            .I(N__35088));
    InMux I__7468 (
            .O(N__35097),
            .I(N__35088));
    LocalMux I__7467 (
            .O(N__35094),
            .I(N__35084));
    InMux I__7466 (
            .O(N__35093),
            .I(N__35081));
    LocalMux I__7465 (
            .O(N__35088),
            .I(N__35078));
    InMux I__7464 (
            .O(N__35087),
            .I(N__35075));
    Span4Mux_v I__7463 (
            .O(N__35084),
            .I(N__35072));
    LocalMux I__7462 (
            .O(N__35081),
            .I(N__35066));
    Span4Mux_v I__7461 (
            .O(N__35078),
            .I(N__35066));
    LocalMux I__7460 (
            .O(N__35075),
            .I(N__35063));
    Span4Mux_h I__7459 (
            .O(N__35072),
            .I(N__35060));
    InMux I__7458 (
            .O(N__35071),
            .I(N__35057));
    Span4Mux_h I__7457 (
            .O(N__35066),
            .I(N__35052));
    Span4Mux_h I__7456 (
            .O(N__35063),
            .I(N__35052));
    Odrv4 I__7455 (
            .O(N__35060),
            .I(rand_data_5));
    LocalMux I__7454 (
            .O(N__35057),
            .I(rand_data_5));
    Odrv4 I__7453 (
            .O(N__35052),
            .I(rand_data_5));
    InMux I__7452 (
            .O(N__35045),
            .I(n16416));
    InMux I__7451 (
            .O(N__35042),
            .I(N__35036));
    InMux I__7450 (
            .O(N__35041),
            .I(N__35033));
    InMux I__7449 (
            .O(N__35040),
            .I(N__35030));
    CascadeMux I__7448 (
            .O(N__35039),
            .I(N__35026));
    LocalMux I__7447 (
            .O(N__35036),
            .I(N__35023));
    LocalMux I__7446 (
            .O(N__35033),
            .I(N__35020));
    LocalMux I__7445 (
            .O(N__35030),
            .I(N__35017));
    InMux I__7444 (
            .O(N__35029),
            .I(N__35014));
    InMux I__7443 (
            .O(N__35026),
            .I(N__35010));
    Span4Mux_h I__7442 (
            .O(N__35023),
            .I(N__35007));
    Span4Mux_v I__7441 (
            .O(N__35020),
            .I(N__35002));
    Span4Mux_h I__7440 (
            .O(N__35017),
            .I(N__35002));
    LocalMux I__7439 (
            .O(N__35014),
            .I(N__34999));
    InMux I__7438 (
            .O(N__35013),
            .I(N__34996));
    LocalMux I__7437 (
            .O(N__35010),
            .I(N__34993));
    Odrv4 I__7436 (
            .O(N__35007),
            .I(rand_data_6));
    Odrv4 I__7435 (
            .O(N__35002),
            .I(rand_data_6));
    Odrv12 I__7434 (
            .O(N__34999),
            .I(rand_data_6));
    LocalMux I__7433 (
            .O(N__34996),
            .I(rand_data_6));
    Odrv12 I__7432 (
            .O(N__34993),
            .I(rand_data_6));
    InMux I__7431 (
            .O(N__34982),
            .I(N__34979));
    LocalMux I__7430 (
            .O(N__34979),
            .I(N__34975));
    InMux I__7429 (
            .O(N__34978),
            .I(N__34972));
    Odrv12 I__7428 (
            .O(N__34975),
            .I(rand_setpoint_6));
    LocalMux I__7427 (
            .O(N__34972),
            .I(rand_setpoint_6));
    InMux I__7426 (
            .O(N__34967),
            .I(n16417));
    InMux I__7425 (
            .O(N__34964),
            .I(N__34960));
    InMux I__7424 (
            .O(N__34963),
            .I(N__34957));
    LocalMux I__7423 (
            .O(N__34960),
            .I(N__34952));
    LocalMux I__7422 (
            .O(N__34957),
            .I(N__34948));
    InMux I__7421 (
            .O(N__34956),
            .I(N__34945));
    InMux I__7420 (
            .O(N__34955),
            .I(N__34942));
    Span4Mux_h I__7419 (
            .O(N__34952),
            .I(N__34939));
    InMux I__7418 (
            .O(N__34951),
            .I(N__34935));
    Span4Mux_h I__7417 (
            .O(N__34948),
            .I(N__34932));
    LocalMux I__7416 (
            .O(N__34945),
            .I(N__34927));
    LocalMux I__7415 (
            .O(N__34942),
            .I(N__34927));
    Span4Mux_v I__7414 (
            .O(N__34939),
            .I(N__34924));
    InMux I__7413 (
            .O(N__34938),
            .I(N__34921));
    LocalMux I__7412 (
            .O(N__34935),
            .I(N__34918));
    Odrv4 I__7411 (
            .O(N__34932),
            .I(rand_data_7));
    Odrv4 I__7410 (
            .O(N__34927),
            .I(rand_data_7));
    Odrv4 I__7409 (
            .O(N__34924),
            .I(rand_data_7));
    LocalMux I__7408 (
            .O(N__34921),
            .I(rand_data_7));
    Odrv12 I__7407 (
            .O(N__34918),
            .I(rand_data_7));
    InMux I__7406 (
            .O(N__34907),
            .I(N__34903));
    CascadeMux I__7405 (
            .O(N__34906),
            .I(N__34900));
    LocalMux I__7404 (
            .O(N__34903),
            .I(N__34897));
    InMux I__7403 (
            .O(N__34900),
            .I(N__34894));
    Odrv4 I__7402 (
            .O(N__34897),
            .I(rand_setpoint_7));
    LocalMux I__7401 (
            .O(N__34894),
            .I(rand_setpoint_7));
    InMux I__7400 (
            .O(N__34889),
            .I(n16418));
    InMux I__7399 (
            .O(N__34886),
            .I(N__34881));
    InMux I__7398 (
            .O(N__34885),
            .I(N__34877));
    InMux I__7397 (
            .O(N__34884),
            .I(N__34874));
    LocalMux I__7396 (
            .O(N__34881),
            .I(N__34871));
    InMux I__7395 (
            .O(N__34880),
            .I(N__34868));
    LocalMux I__7394 (
            .O(N__34877),
            .I(N__34862));
    LocalMux I__7393 (
            .O(N__34874),
            .I(N__34862));
    Span4Mux_v I__7392 (
            .O(N__34871),
            .I(N__34857));
    LocalMux I__7391 (
            .O(N__34868),
            .I(N__34857));
    InMux I__7390 (
            .O(N__34867),
            .I(N__34853));
    Span4Mux_h I__7389 (
            .O(N__34862),
            .I(N__34850));
    Span4Mux_h I__7388 (
            .O(N__34857),
            .I(N__34847));
    InMux I__7387 (
            .O(N__34856),
            .I(N__34844));
    LocalMux I__7386 (
            .O(N__34853),
            .I(N__34841));
    Odrv4 I__7385 (
            .O(N__34850),
            .I(rand_data_8));
    Odrv4 I__7384 (
            .O(N__34847),
            .I(rand_data_8));
    LocalMux I__7383 (
            .O(N__34844),
            .I(rand_data_8));
    Odrv12 I__7382 (
            .O(N__34841),
            .I(rand_data_8));
    InMux I__7381 (
            .O(N__34832),
            .I(bfn_9_30_0_));
    InMux I__7380 (
            .O(N__34829),
            .I(N__34826));
    LocalMux I__7379 (
            .O(N__34826),
            .I(N__34821));
    InMux I__7378 (
            .O(N__34825),
            .I(N__34818));
    InMux I__7377 (
            .O(N__34824),
            .I(N__34814));
    Span4Mux_v I__7376 (
            .O(N__34821),
            .I(N__34808));
    LocalMux I__7375 (
            .O(N__34818),
            .I(N__34808));
    InMux I__7374 (
            .O(N__34817),
            .I(N__34805));
    LocalMux I__7373 (
            .O(N__34814),
            .I(N__34802));
    InMux I__7372 (
            .O(N__34813),
            .I(N__34798));
    Span4Mux_h I__7371 (
            .O(N__34808),
            .I(N__34795));
    LocalMux I__7370 (
            .O(N__34805),
            .I(N__34792));
    Span4Mux_h I__7369 (
            .O(N__34802),
            .I(N__34789));
    InMux I__7368 (
            .O(N__34801),
            .I(N__34786));
    LocalMux I__7367 (
            .O(N__34798),
            .I(N__34783));
    Odrv4 I__7366 (
            .O(N__34795),
            .I(rand_data_9));
    Odrv4 I__7365 (
            .O(N__34792),
            .I(rand_data_9));
    Odrv4 I__7364 (
            .O(N__34789),
            .I(rand_data_9));
    LocalMux I__7363 (
            .O(N__34786),
            .I(rand_data_9));
    Odrv12 I__7362 (
            .O(N__34783),
            .I(rand_data_9));
    InMux I__7361 (
            .O(N__34772),
            .I(n16420));
    InMux I__7360 (
            .O(N__34769),
            .I(N__34766));
    LocalMux I__7359 (
            .O(N__34766),
            .I(N__34761));
    InMux I__7358 (
            .O(N__34765),
            .I(N__34758));
    InMux I__7357 (
            .O(N__34764),
            .I(N__34754));
    Span4Mux_v I__7356 (
            .O(N__34761),
            .I(N__34749));
    LocalMux I__7355 (
            .O(N__34758),
            .I(N__34749));
    InMux I__7354 (
            .O(N__34757),
            .I(N__34746));
    LocalMux I__7353 (
            .O(N__34754),
            .I(N__34742));
    Span4Mux_v I__7352 (
            .O(N__34749),
            .I(N__34737));
    LocalMux I__7351 (
            .O(N__34746),
            .I(N__34737));
    InMux I__7350 (
            .O(N__34745),
            .I(N__34733));
    Span4Mux_h I__7349 (
            .O(N__34742),
            .I(N__34730));
    Span4Mux_h I__7348 (
            .O(N__34737),
            .I(N__34727));
    InMux I__7347 (
            .O(N__34736),
            .I(N__34724));
    LocalMux I__7346 (
            .O(N__34733),
            .I(N__34721));
    Odrv4 I__7345 (
            .O(N__34730),
            .I(rand_data_10));
    Odrv4 I__7344 (
            .O(N__34727),
            .I(rand_data_10));
    LocalMux I__7343 (
            .O(N__34724),
            .I(rand_data_10));
    Odrv12 I__7342 (
            .O(N__34721),
            .I(rand_data_10));
    InMux I__7341 (
            .O(N__34712),
            .I(n16421));
    InMux I__7340 (
            .O(N__34709),
            .I(N__34706));
    LocalMux I__7339 (
            .O(N__34706),
            .I(N__34702));
    InMux I__7338 (
            .O(N__34705),
            .I(N__34699));
    Odrv12 I__7337 (
            .O(N__34702),
            .I(data_in_13_2));
    LocalMux I__7336 (
            .O(N__34699),
            .I(data_in_13_2));
    InMux I__7335 (
            .O(N__34694),
            .I(N__34688));
    InMux I__7334 (
            .O(N__34693),
            .I(N__34688));
    LocalMux I__7333 (
            .O(N__34688),
            .I(data_in_12_2));
    InMux I__7332 (
            .O(N__34685),
            .I(N__34680));
    InMux I__7331 (
            .O(N__34684),
            .I(N__34676));
    InMux I__7330 (
            .O(N__34683),
            .I(N__34669));
    LocalMux I__7329 (
            .O(N__34680),
            .I(N__34666));
    InMux I__7328 (
            .O(N__34679),
            .I(N__34663));
    LocalMux I__7327 (
            .O(N__34676),
            .I(N__34656));
    InMux I__7326 (
            .O(N__34675),
            .I(N__34653));
    InMux I__7325 (
            .O(N__34674),
            .I(N__34648));
    InMux I__7324 (
            .O(N__34673),
            .I(N__34648));
    InMux I__7323 (
            .O(N__34672),
            .I(N__34645));
    LocalMux I__7322 (
            .O(N__34669),
            .I(N__34637));
    Span4Mux_v I__7321 (
            .O(N__34666),
            .I(N__34632));
    LocalMux I__7320 (
            .O(N__34663),
            .I(N__34632));
    InMux I__7319 (
            .O(N__34662),
            .I(N__34629));
    CascadeMux I__7318 (
            .O(N__34661),
            .I(N__34623));
    InMux I__7317 (
            .O(N__34660),
            .I(N__34619));
    InMux I__7316 (
            .O(N__34659),
            .I(N__34616));
    Span4Mux_s2_h I__7315 (
            .O(N__34656),
            .I(N__34607));
    LocalMux I__7314 (
            .O(N__34653),
            .I(N__34607));
    LocalMux I__7313 (
            .O(N__34648),
            .I(N__34607));
    LocalMux I__7312 (
            .O(N__34645),
            .I(N__34607));
    CascadeMux I__7311 (
            .O(N__34644),
            .I(N__34602));
    InMux I__7310 (
            .O(N__34643),
            .I(N__34598));
    CascadeMux I__7309 (
            .O(N__34642),
            .I(N__34595));
    InMux I__7308 (
            .O(N__34641),
            .I(N__34589));
    InMux I__7307 (
            .O(N__34640),
            .I(N__34589));
    Span4Mux_v I__7306 (
            .O(N__34637),
            .I(N__34582));
    Span4Mux_v I__7305 (
            .O(N__34632),
            .I(N__34582));
    LocalMux I__7304 (
            .O(N__34629),
            .I(N__34582));
    InMux I__7303 (
            .O(N__34628),
            .I(N__34577));
    InMux I__7302 (
            .O(N__34627),
            .I(N__34577));
    InMux I__7301 (
            .O(N__34626),
            .I(N__34562));
    InMux I__7300 (
            .O(N__34623),
            .I(N__34562));
    InMux I__7299 (
            .O(N__34622),
            .I(N__34562));
    LocalMux I__7298 (
            .O(N__34619),
            .I(N__34555));
    LocalMux I__7297 (
            .O(N__34616),
            .I(N__34555));
    Span4Mux_v I__7296 (
            .O(N__34607),
            .I(N__34555));
    InMux I__7295 (
            .O(N__34606),
            .I(N__34545));
    InMux I__7294 (
            .O(N__34605),
            .I(N__34542));
    InMux I__7293 (
            .O(N__34602),
            .I(N__34537));
    InMux I__7292 (
            .O(N__34601),
            .I(N__34537));
    LocalMux I__7291 (
            .O(N__34598),
            .I(N__34534));
    InMux I__7290 (
            .O(N__34595),
            .I(N__34529));
    InMux I__7289 (
            .O(N__34594),
            .I(N__34529));
    LocalMux I__7288 (
            .O(N__34589),
            .I(N__34522));
    Span4Mux_h I__7287 (
            .O(N__34582),
            .I(N__34522));
    LocalMux I__7286 (
            .O(N__34577),
            .I(N__34522));
    InMux I__7285 (
            .O(N__34576),
            .I(N__34515));
    InMux I__7284 (
            .O(N__34575),
            .I(N__34515));
    InMux I__7283 (
            .O(N__34574),
            .I(N__34515));
    InMux I__7282 (
            .O(N__34573),
            .I(N__34510));
    InMux I__7281 (
            .O(N__34572),
            .I(N__34510));
    InMux I__7280 (
            .O(N__34571),
            .I(N__34503));
    InMux I__7279 (
            .O(N__34570),
            .I(N__34503));
    InMux I__7278 (
            .O(N__34569),
            .I(N__34503));
    LocalMux I__7277 (
            .O(N__34562),
            .I(N__34498));
    Span4Mux_h I__7276 (
            .O(N__34555),
            .I(N__34498));
    InMux I__7275 (
            .O(N__34554),
            .I(N__34491));
    InMux I__7274 (
            .O(N__34553),
            .I(N__34491));
    InMux I__7273 (
            .O(N__34552),
            .I(N__34491));
    InMux I__7272 (
            .O(N__34551),
            .I(N__34482));
    InMux I__7271 (
            .O(N__34550),
            .I(N__34482));
    InMux I__7270 (
            .O(N__34549),
            .I(N__34482));
    InMux I__7269 (
            .O(N__34548),
            .I(N__34482));
    LocalMux I__7268 (
            .O(N__34545),
            .I(FRAME_MATCHER_next_state_31_N_2026_1));
    LocalMux I__7267 (
            .O(N__34542),
            .I(FRAME_MATCHER_next_state_31_N_2026_1));
    LocalMux I__7266 (
            .O(N__34537),
            .I(FRAME_MATCHER_next_state_31_N_2026_1));
    Odrv4 I__7265 (
            .O(N__34534),
            .I(FRAME_MATCHER_next_state_31_N_2026_1));
    LocalMux I__7264 (
            .O(N__34529),
            .I(FRAME_MATCHER_next_state_31_N_2026_1));
    Odrv4 I__7263 (
            .O(N__34522),
            .I(FRAME_MATCHER_next_state_31_N_2026_1));
    LocalMux I__7262 (
            .O(N__34515),
            .I(FRAME_MATCHER_next_state_31_N_2026_1));
    LocalMux I__7261 (
            .O(N__34510),
            .I(FRAME_MATCHER_next_state_31_N_2026_1));
    LocalMux I__7260 (
            .O(N__34503),
            .I(FRAME_MATCHER_next_state_31_N_2026_1));
    Odrv4 I__7259 (
            .O(N__34498),
            .I(FRAME_MATCHER_next_state_31_N_2026_1));
    LocalMux I__7258 (
            .O(N__34491),
            .I(FRAME_MATCHER_next_state_31_N_2026_1));
    LocalMux I__7257 (
            .O(N__34482),
            .I(FRAME_MATCHER_next_state_31_N_2026_1));
    InMux I__7256 (
            .O(N__34457),
            .I(N__34449));
    InMux I__7255 (
            .O(N__34456),
            .I(N__34437));
    InMux I__7254 (
            .O(N__34455),
            .I(N__34437));
    InMux I__7253 (
            .O(N__34454),
            .I(N__34437));
    InMux I__7252 (
            .O(N__34453),
            .I(N__34430));
    InMux I__7251 (
            .O(N__34452),
            .I(N__34427));
    LocalMux I__7250 (
            .O(N__34449),
            .I(N__34423));
    InMux I__7249 (
            .O(N__34448),
            .I(N__34420));
    InMux I__7248 (
            .O(N__34447),
            .I(N__34417));
    InMux I__7247 (
            .O(N__34446),
            .I(N__34414));
    InMux I__7246 (
            .O(N__34445),
            .I(N__34409));
    InMux I__7245 (
            .O(N__34444),
            .I(N__34409));
    LocalMux I__7244 (
            .O(N__34437),
            .I(N__34405));
    InMux I__7243 (
            .O(N__34436),
            .I(N__34400));
    InMux I__7242 (
            .O(N__34435),
            .I(N__34400));
    InMux I__7241 (
            .O(N__34434),
            .I(N__34395));
    InMux I__7240 (
            .O(N__34433),
            .I(N__34395));
    LocalMux I__7239 (
            .O(N__34430),
            .I(N__34390));
    LocalMux I__7238 (
            .O(N__34427),
            .I(N__34387));
    InMux I__7237 (
            .O(N__34426),
            .I(N__34384));
    Span4Mux_v I__7236 (
            .O(N__34423),
            .I(N__34379));
    LocalMux I__7235 (
            .O(N__34420),
            .I(N__34379));
    LocalMux I__7234 (
            .O(N__34417),
            .I(N__34376));
    LocalMux I__7233 (
            .O(N__34414),
            .I(N__34371));
    LocalMux I__7232 (
            .O(N__34409),
            .I(N__34371));
    CascadeMux I__7231 (
            .O(N__34408),
            .I(N__34368));
    Span4Mux_v I__7230 (
            .O(N__34405),
            .I(N__34362));
    LocalMux I__7229 (
            .O(N__34400),
            .I(N__34362));
    LocalMux I__7228 (
            .O(N__34395),
            .I(N__34359));
    InMux I__7227 (
            .O(N__34394),
            .I(N__34354));
    InMux I__7226 (
            .O(N__34393),
            .I(N__34354));
    Span4Mux_v I__7225 (
            .O(N__34390),
            .I(N__34341));
    Span4Mux_h I__7224 (
            .O(N__34387),
            .I(N__34341));
    LocalMux I__7223 (
            .O(N__34384),
            .I(N__34341));
    Span4Mux_v I__7222 (
            .O(N__34379),
            .I(N__34341));
    Span4Mux_h I__7221 (
            .O(N__34376),
            .I(N__34341));
    Span4Mux_v I__7220 (
            .O(N__34371),
            .I(N__34341));
    InMux I__7219 (
            .O(N__34368),
            .I(N__34336));
    InMux I__7218 (
            .O(N__34367),
            .I(N__34336));
    Odrv4 I__7217 (
            .O(N__34362),
            .I(n63_adj_2642));
    Odrv12 I__7216 (
            .O(N__34359),
            .I(n63_adj_2642));
    LocalMux I__7215 (
            .O(N__34354),
            .I(n63_adj_2642));
    Odrv4 I__7214 (
            .O(N__34341),
            .I(n63_adj_2642));
    LocalMux I__7213 (
            .O(N__34336),
            .I(n63_adj_2642));
    InMux I__7212 (
            .O(N__34325),
            .I(N__34322));
    LocalMux I__7211 (
            .O(N__34322),
            .I(N__34319));
    Span4Mux_v I__7210 (
            .O(N__34319),
            .I(N__34315));
    InMux I__7209 (
            .O(N__34318),
            .I(N__34312));
    Span4Mux_v I__7208 (
            .O(N__34315),
            .I(N__34309));
    LocalMux I__7207 (
            .O(N__34312),
            .I(N__34304));
    Span4Mux_h I__7206 (
            .O(N__34309),
            .I(N__34301));
    InMux I__7205 (
            .O(N__34308),
            .I(N__34296));
    InMux I__7204 (
            .O(N__34307),
            .I(N__34296));
    Odrv4 I__7203 (
            .O(N__34304),
            .I(n63));
    Odrv4 I__7202 (
            .O(N__34301),
            .I(n63));
    LocalMux I__7201 (
            .O(N__34296),
            .I(n63));
    InMux I__7200 (
            .O(N__34289),
            .I(N__34285));
    CascadeMux I__7199 (
            .O(N__34288),
            .I(N__34282));
    LocalMux I__7198 (
            .O(N__34285),
            .I(N__34279));
    InMux I__7197 (
            .O(N__34282),
            .I(N__34276));
    Span4Mux_v I__7196 (
            .O(N__34279),
            .I(N__34273));
    LocalMux I__7195 (
            .O(N__34276),
            .I(FRAME_MATCHER_next_state_0));
    Odrv4 I__7194 (
            .O(N__34273),
            .I(FRAME_MATCHER_next_state_0));
    InMux I__7193 (
            .O(N__34268),
            .I(N__34265));
    LocalMux I__7192 (
            .O(N__34265),
            .I(N__34261));
    InMux I__7191 (
            .O(N__34264),
            .I(N__34258));
    Odrv4 I__7190 (
            .O(N__34261),
            .I(data_in_17_5));
    LocalMux I__7189 (
            .O(N__34258),
            .I(data_in_17_5));
    InMux I__7188 (
            .O(N__34253),
            .I(N__34250));
    LocalMux I__7187 (
            .O(N__34250),
            .I(N__34247));
    Span4Mux_h I__7186 (
            .O(N__34247),
            .I(N__34242));
    InMux I__7185 (
            .O(N__34246),
            .I(N__34237));
    InMux I__7184 (
            .O(N__34245),
            .I(N__34237));
    Odrv4 I__7183 (
            .O(N__34242),
            .I(\c0.rx.r_SM_Main_2_N_2386_0 ));
    LocalMux I__7182 (
            .O(N__34237),
            .I(\c0.rx.r_SM_Main_2_N_2386_0 ));
    InMux I__7181 (
            .O(N__34232),
            .I(N__34229));
    LocalMux I__7180 (
            .O(N__34229),
            .I(N__34226));
    Span4Mux_h I__7179 (
            .O(N__34226),
            .I(N__34223));
    Odrv4 I__7178 (
            .O(N__34223),
            .I(\c0.rx.n18066 ));
    InMux I__7177 (
            .O(N__34220),
            .I(N__34214));
    InMux I__7176 (
            .O(N__34219),
            .I(N__34214));
    LocalMux I__7175 (
            .O(N__34214),
            .I(N__34208));
    InMux I__7174 (
            .O(N__34213),
            .I(N__34205));
    InMux I__7173 (
            .O(N__34212),
            .I(N__34202));
    InMux I__7172 (
            .O(N__34211),
            .I(N__34198));
    Span4Mux_v I__7171 (
            .O(N__34208),
            .I(N__34195));
    LocalMux I__7170 (
            .O(N__34205),
            .I(N__34192));
    LocalMux I__7169 (
            .O(N__34202),
            .I(N__34189));
    InMux I__7168 (
            .O(N__34201),
            .I(N__34186));
    LocalMux I__7167 (
            .O(N__34198),
            .I(N__34183));
    Span4Mux_h I__7166 (
            .O(N__34195),
            .I(N__34180));
    Span4Mux_s3_h I__7165 (
            .O(N__34192),
            .I(N__34171));
    Span4Mux_v I__7164 (
            .O(N__34189),
            .I(N__34171));
    LocalMux I__7163 (
            .O(N__34186),
            .I(N__34171));
    Span4Mux_h I__7162 (
            .O(N__34183),
            .I(N__34171));
    Odrv4 I__7161 (
            .O(N__34180),
            .I(rand_data_0));
    Odrv4 I__7160 (
            .O(N__34171),
            .I(rand_data_0));
    InMux I__7159 (
            .O(N__34166),
            .I(N__34161));
    InMux I__7158 (
            .O(N__34165),
            .I(N__34155));
    InMux I__7157 (
            .O(N__34164),
            .I(N__34155));
    LocalMux I__7156 (
            .O(N__34161),
            .I(N__34152));
    InMux I__7155 (
            .O(N__34160),
            .I(N__34149));
    LocalMux I__7154 (
            .O(N__34155),
            .I(N__34145));
    Span4Mux_s3_h I__7153 (
            .O(N__34152),
            .I(N__34140));
    LocalMux I__7152 (
            .O(N__34149),
            .I(N__34140));
    InMux I__7151 (
            .O(N__34148),
            .I(N__34136));
    Span4Mux_h I__7150 (
            .O(N__34145),
            .I(N__34133));
    Span4Mux_v I__7149 (
            .O(N__34140),
            .I(N__34130));
    InMux I__7148 (
            .O(N__34139),
            .I(N__34127));
    LocalMux I__7147 (
            .O(N__34136),
            .I(N__34124));
    Odrv4 I__7146 (
            .O(N__34133),
            .I(rand_data_1));
    Odrv4 I__7145 (
            .O(N__34130),
            .I(rand_data_1));
    LocalMux I__7144 (
            .O(N__34127),
            .I(rand_data_1));
    Odrv12 I__7143 (
            .O(N__34124),
            .I(rand_data_1));
    InMux I__7142 (
            .O(N__34115),
            .I(n16412));
    InMux I__7141 (
            .O(N__34112),
            .I(N__34109));
    LocalMux I__7140 (
            .O(N__34109),
            .I(N__34105));
    InMux I__7139 (
            .O(N__34108),
            .I(N__34102));
    Span4Mux_v I__7138 (
            .O(N__34105),
            .I(N__34095));
    LocalMux I__7137 (
            .O(N__34102),
            .I(N__34095));
    InMux I__7136 (
            .O(N__34101),
            .I(N__34092));
    InMux I__7135 (
            .O(N__34100),
            .I(N__34089));
    Span4Mux_h I__7134 (
            .O(N__34095),
            .I(N__34085));
    LocalMux I__7133 (
            .O(N__34092),
            .I(N__34082));
    LocalMux I__7132 (
            .O(N__34089),
            .I(N__34079));
    InMux I__7131 (
            .O(N__34088),
            .I(N__34075));
    Sp12to4 I__7130 (
            .O(N__34085),
            .I(N__34070));
    Span12Mux_s4_h I__7129 (
            .O(N__34082),
            .I(N__34070));
    Span4Mux_h I__7128 (
            .O(N__34079),
            .I(N__34067));
    InMux I__7127 (
            .O(N__34078),
            .I(N__34064));
    LocalMux I__7126 (
            .O(N__34075),
            .I(N__34061));
    Odrv12 I__7125 (
            .O(N__34070),
            .I(rand_data_2));
    Odrv4 I__7124 (
            .O(N__34067),
            .I(rand_data_2));
    LocalMux I__7123 (
            .O(N__34064),
            .I(rand_data_2));
    Odrv12 I__7122 (
            .O(N__34061),
            .I(rand_data_2));
    InMux I__7121 (
            .O(N__34052),
            .I(n16413));
    InMux I__7120 (
            .O(N__34049),
            .I(N__34046));
    LocalMux I__7119 (
            .O(N__34046),
            .I(N__34042));
    InMux I__7118 (
            .O(N__34045),
            .I(N__34039));
    Odrv4 I__7117 (
            .O(N__34042),
            .I(data_in_16_2));
    LocalMux I__7116 (
            .O(N__34039),
            .I(data_in_16_2));
    InMux I__7115 (
            .O(N__34034),
            .I(N__34030));
    InMux I__7114 (
            .O(N__34033),
            .I(N__34027));
    LocalMux I__7113 (
            .O(N__34030),
            .I(N__34024));
    LocalMux I__7112 (
            .O(N__34027),
            .I(N__34021));
    Span4Mux_h I__7111 (
            .O(N__34024),
            .I(N__34018));
    Span4Mux_v I__7110 (
            .O(N__34021),
            .I(N__34015));
    Sp12to4 I__7109 (
            .O(N__34018),
            .I(N__34012));
    Span4Mux_v I__7108 (
            .O(N__34015),
            .I(N__34009));
    Span12Mux_v I__7107 (
            .O(N__34012),
            .I(N__34006));
    Span4Mux_h I__7106 (
            .O(N__34009),
            .I(N__34003));
    Odrv12 I__7105 (
            .O(N__34006),
            .I(n4));
    Odrv4 I__7104 (
            .O(N__34003),
            .I(n4));
    InMux I__7103 (
            .O(N__33998),
            .I(N__33994));
    CascadeMux I__7102 (
            .O(N__33997),
            .I(N__33991));
    LocalMux I__7101 (
            .O(N__33994),
            .I(N__33988));
    InMux I__7100 (
            .O(N__33991),
            .I(N__33985));
    Odrv12 I__7099 (
            .O(N__33988),
            .I(rx_data_3));
    LocalMux I__7098 (
            .O(N__33985),
            .I(rx_data_3));
    InMux I__7097 (
            .O(N__33980),
            .I(N__33977));
    LocalMux I__7096 (
            .O(N__33977),
            .I(N__33973));
    InMux I__7095 (
            .O(N__33976),
            .I(N__33970));
    Span4Mux_h I__7094 (
            .O(N__33973),
            .I(N__33965));
    LocalMux I__7093 (
            .O(N__33970),
            .I(N__33965));
    Span4Mux_v I__7092 (
            .O(N__33965),
            .I(N__33962));
    Span4Mux_v I__7091 (
            .O(N__33962),
            .I(N__33959));
    Span4Mux_h I__7090 (
            .O(N__33959),
            .I(N__33956));
    Odrv4 I__7089 (
            .O(N__33956),
            .I(n4_adj_2582));
    InMux I__7088 (
            .O(N__33953),
            .I(N__33949));
    InMux I__7087 (
            .O(N__33952),
            .I(N__33946));
    LocalMux I__7086 (
            .O(N__33949),
            .I(data_in_20_6));
    LocalMux I__7085 (
            .O(N__33946),
            .I(data_in_20_6));
    InMux I__7084 (
            .O(N__33941),
            .I(N__33938));
    LocalMux I__7083 (
            .O(N__33938),
            .I(N__33935));
    Span4Mux_h I__7082 (
            .O(N__33935),
            .I(N__33932));
    Span4Mux_h I__7081 (
            .O(N__33932),
            .I(N__33928));
    InMux I__7080 (
            .O(N__33931),
            .I(N__33925));
    Span4Mux_v I__7079 (
            .O(N__33928),
            .I(N__33919));
    LocalMux I__7078 (
            .O(N__33925),
            .I(N__33919));
    InMux I__7077 (
            .O(N__33924),
            .I(N__33916));
    Odrv4 I__7076 (
            .O(N__33919),
            .I(data_in_8_2));
    LocalMux I__7075 (
            .O(N__33916),
            .I(data_in_8_2));
    CascadeMux I__7074 (
            .O(N__33911),
            .I(N__33907));
    CascadeMux I__7073 (
            .O(N__33910),
            .I(N__33904));
    InMux I__7072 (
            .O(N__33907),
            .I(N__33895));
    InMux I__7071 (
            .O(N__33904),
            .I(N__33895));
    InMux I__7070 (
            .O(N__33903),
            .I(N__33895));
    InMux I__7069 (
            .O(N__33902),
            .I(N__33892));
    LocalMux I__7068 (
            .O(N__33895),
            .I(N__33887));
    LocalMux I__7067 (
            .O(N__33892),
            .I(N__33887));
    Span4Mux_v I__7066 (
            .O(N__33887),
            .I(N__33884));
    Odrv4 I__7065 (
            .O(N__33884),
            .I(n8567));
    InMux I__7064 (
            .O(N__33881),
            .I(N__33878));
    LocalMux I__7063 (
            .O(N__33878),
            .I(N__33874));
    InMux I__7062 (
            .O(N__33877),
            .I(N__33871));
    Odrv12 I__7061 (
            .O(N__33874),
            .I(data_in_11_2));
    LocalMux I__7060 (
            .O(N__33871),
            .I(data_in_11_2));
    CascadeMux I__7059 (
            .O(N__33866),
            .I(n9390_cascade_));
    CascadeMux I__7058 (
            .O(N__33863),
            .I(n17681_cascade_));
    InMux I__7057 (
            .O(N__33860),
            .I(N__33856));
    InMux I__7056 (
            .O(N__33859),
            .I(N__33853));
    LocalMux I__7055 (
            .O(N__33856),
            .I(N__33849));
    LocalMux I__7054 (
            .O(N__33853),
            .I(N__33846));
    InMux I__7053 (
            .O(N__33852),
            .I(N__33843));
    Span4Mux_h I__7052 (
            .O(N__33849),
            .I(N__33840));
    Odrv4 I__7051 (
            .O(N__33846),
            .I(n16466));
    LocalMux I__7050 (
            .O(N__33843),
            .I(n16466));
    Odrv4 I__7049 (
            .O(N__33840),
            .I(n16466));
    InMux I__7048 (
            .O(N__33833),
            .I(N__33828));
    InMux I__7047 (
            .O(N__33832),
            .I(N__33825));
    InMux I__7046 (
            .O(N__33831),
            .I(N__33822));
    LocalMux I__7045 (
            .O(N__33828),
            .I(N__33819));
    LocalMux I__7044 (
            .O(N__33825),
            .I(N__33814));
    LocalMux I__7043 (
            .O(N__33822),
            .I(N__33814));
    Span4Mux_h I__7042 (
            .O(N__33819),
            .I(N__33811));
    Span4Mux_h I__7041 (
            .O(N__33814),
            .I(N__33808));
    Odrv4 I__7040 (
            .O(N__33811),
            .I(n17356));
    Odrv4 I__7039 (
            .O(N__33808),
            .I(n17356));
    InMux I__7038 (
            .O(N__33803),
            .I(N__33800));
    LocalMux I__7037 (
            .O(N__33800),
            .I(N__33797));
    Odrv12 I__7036 (
            .O(N__33797),
            .I(n18102));
    InMux I__7035 (
            .O(N__33794),
            .I(N__33790));
    InMux I__7034 (
            .O(N__33793),
            .I(N__33786));
    LocalMux I__7033 (
            .O(N__33790),
            .I(N__33783));
    InMux I__7032 (
            .O(N__33789),
            .I(N__33780));
    LocalMux I__7031 (
            .O(N__33786),
            .I(N__33773));
    Span4Mux_h I__7030 (
            .O(N__33783),
            .I(N__33773));
    LocalMux I__7029 (
            .O(N__33780),
            .I(N__33773));
    Odrv4 I__7028 (
            .O(N__33773),
            .I(r_Clock_Count_2));
    InMux I__7027 (
            .O(N__33770),
            .I(N__33767));
    LocalMux I__7026 (
            .O(N__33767),
            .I(n13601));
    InMux I__7025 (
            .O(N__33764),
            .I(N__33760));
    InMux I__7024 (
            .O(N__33763),
            .I(N__33757));
    LocalMux I__7023 (
            .O(N__33760),
            .I(N__33754));
    LocalMux I__7022 (
            .O(N__33757),
            .I(N__33751));
    Span4Mux_h I__7021 (
            .O(N__33754),
            .I(N__33747));
    Span4Mux_h I__7020 (
            .O(N__33751),
            .I(N__33744));
    InMux I__7019 (
            .O(N__33750),
            .I(N__33741));
    Span4Mux_h I__7018 (
            .O(N__33747),
            .I(N__33738));
    Odrv4 I__7017 (
            .O(N__33744),
            .I(data_in_7_2));
    LocalMux I__7016 (
            .O(N__33741),
            .I(data_in_7_2));
    Odrv4 I__7015 (
            .O(N__33738),
            .I(data_in_7_2));
    InMux I__7014 (
            .O(N__33731),
            .I(N__33728));
    LocalMux I__7013 (
            .O(N__33728),
            .I(N__33725));
    Span4Mux_h I__7012 (
            .O(N__33725),
            .I(N__33721));
    InMux I__7011 (
            .O(N__33724),
            .I(N__33718));
    Odrv4 I__7010 (
            .O(N__33721),
            .I(n13597));
    LocalMux I__7009 (
            .O(N__33718),
            .I(n13597));
    InMux I__7008 (
            .O(N__33713),
            .I(N__33710));
    LocalMux I__7007 (
            .O(N__33710),
            .I(N__33706));
    InMux I__7006 (
            .O(N__33709),
            .I(N__33703));
    Odrv4 I__7005 (
            .O(N__33706),
            .I(rx_data_6));
    LocalMux I__7004 (
            .O(N__33703),
            .I(rx_data_6));
    CascadeMux I__7003 (
            .O(N__33698),
            .I(N__33694));
    CascadeMux I__7002 (
            .O(N__33697),
            .I(N__33689));
    InMux I__7001 (
            .O(N__33694),
            .I(N__33686));
    CascadeMux I__7000 (
            .O(N__33693),
            .I(N__33683));
    CascadeMux I__6999 (
            .O(N__33692),
            .I(N__33679));
    InMux I__6998 (
            .O(N__33689),
            .I(N__33674));
    LocalMux I__6997 (
            .O(N__33686),
            .I(N__33671));
    InMux I__6996 (
            .O(N__33683),
            .I(N__33668));
    InMux I__6995 (
            .O(N__33682),
            .I(N__33663));
    InMux I__6994 (
            .O(N__33679),
            .I(N__33660));
    CascadeMux I__6993 (
            .O(N__33678),
            .I(N__33657));
    CascadeMux I__6992 (
            .O(N__33677),
            .I(N__33654));
    LocalMux I__6991 (
            .O(N__33674),
            .I(N__33651));
    Span4Mux_h I__6990 (
            .O(N__33671),
            .I(N__33646));
    LocalMux I__6989 (
            .O(N__33668),
            .I(N__33646));
    InMux I__6988 (
            .O(N__33667),
            .I(N__33640));
    InMux I__6987 (
            .O(N__33666),
            .I(N__33640));
    LocalMux I__6986 (
            .O(N__33663),
            .I(N__33637));
    LocalMux I__6985 (
            .O(N__33660),
            .I(N__33634));
    InMux I__6984 (
            .O(N__33657),
            .I(N__33630));
    InMux I__6983 (
            .O(N__33654),
            .I(N__33627));
    Span4Mux_s2_h I__6982 (
            .O(N__33651),
            .I(N__33622));
    Span4Mux_v I__6981 (
            .O(N__33646),
            .I(N__33622));
    InMux I__6980 (
            .O(N__33645),
            .I(N__33619));
    LocalMux I__6979 (
            .O(N__33640),
            .I(N__33614));
    Span4Mux_v I__6978 (
            .O(N__33637),
            .I(N__33614));
    Span4Mux_s2_h I__6977 (
            .O(N__33634),
            .I(N__33611));
    SRMux I__6976 (
            .O(N__33633),
            .I(N__33608));
    LocalMux I__6975 (
            .O(N__33630),
            .I(N__33605));
    LocalMux I__6974 (
            .O(N__33627),
            .I(N__33600));
    Span4Mux_h I__6973 (
            .O(N__33622),
            .I(N__33600));
    LocalMux I__6972 (
            .O(N__33619),
            .I(N__33595));
    Sp12to4 I__6971 (
            .O(N__33614),
            .I(N__33595));
    Span4Mux_v I__6970 (
            .O(N__33611),
            .I(N__33592));
    LocalMux I__6969 (
            .O(N__33608),
            .I(N__33589));
    Span12Mux_s3_h I__6968 (
            .O(N__33605),
            .I(N__33586));
    Span4Mux_v I__6967 (
            .O(N__33600),
            .I(N__33583));
    Span12Mux_h I__6966 (
            .O(N__33595),
            .I(N__33580));
    Span4Mux_v I__6965 (
            .O(N__33592),
            .I(N__33577));
    Sp12to4 I__6964 (
            .O(N__33589),
            .I(N__33572));
    Span12Mux_v I__6963 (
            .O(N__33586),
            .I(N__33572));
    Span4Mux_v I__6962 (
            .O(N__33583),
            .I(N__33569));
    Odrv12 I__6961 (
            .O(N__33580),
            .I(\c0.n142 ));
    Odrv4 I__6960 (
            .O(N__33577),
            .I(\c0.n142 ));
    Odrv12 I__6959 (
            .O(N__33572),
            .I(\c0.n142 ));
    Odrv4 I__6958 (
            .O(N__33569),
            .I(\c0.n142 ));
    SRMux I__6957 (
            .O(N__33560),
            .I(N__33557));
    LocalMux I__6956 (
            .O(N__33557),
            .I(N__33554));
    Span4Mux_h I__6955 (
            .O(N__33554),
            .I(N__33551));
    Odrv4 I__6954 (
            .O(N__33551),
            .I(\c0.n1 ));
    CascadeMux I__6953 (
            .O(N__33548),
            .I(N__33544));
    InMux I__6952 (
            .O(N__33547),
            .I(N__33541));
    InMux I__6951 (
            .O(N__33544),
            .I(N__33538));
    LocalMux I__6950 (
            .O(N__33541),
            .I(N__33535));
    LocalMux I__6949 (
            .O(N__33538),
            .I(FRAME_MATCHER_next_state_1));
    Odrv12 I__6948 (
            .O(N__33535),
            .I(FRAME_MATCHER_next_state_1));
    CascadeMux I__6947 (
            .O(N__33530),
            .I(N__33526));
    CascadeMux I__6946 (
            .O(N__33529),
            .I(N__33523));
    InMux I__6945 (
            .O(N__33526),
            .I(N__33519));
    InMux I__6944 (
            .O(N__33523),
            .I(N__33509));
    InMux I__6943 (
            .O(N__33522),
            .I(N__33509));
    LocalMux I__6942 (
            .O(N__33519),
            .I(N__33505));
    InMux I__6941 (
            .O(N__33518),
            .I(N__33498));
    InMux I__6940 (
            .O(N__33517),
            .I(N__33498));
    InMux I__6939 (
            .O(N__33516),
            .I(N__33498));
    InMux I__6938 (
            .O(N__33515),
            .I(N__33495));
    InMux I__6937 (
            .O(N__33514),
            .I(N__33492));
    LocalMux I__6936 (
            .O(N__33509),
            .I(N__33488));
    InMux I__6935 (
            .O(N__33508),
            .I(N__33485));
    Span4Mux_v I__6934 (
            .O(N__33505),
            .I(N__33480));
    LocalMux I__6933 (
            .O(N__33498),
            .I(N__33480));
    LocalMux I__6932 (
            .O(N__33495),
            .I(N__33477));
    LocalMux I__6931 (
            .O(N__33492),
            .I(N__33474));
    InMux I__6930 (
            .O(N__33491),
            .I(N__33471));
    Span4Mux_s3_h I__6929 (
            .O(N__33488),
            .I(N__33468));
    LocalMux I__6928 (
            .O(N__33485),
            .I(N__33465));
    Span4Mux_v I__6927 (
            .O(N__33480),
            .I(N__33462));
    Sp12to4 I__6926 (
            .O(N__33477),
            .I(N__33456));
    Span4Mux_v I__6925 (
            .O(N__33474),
            .I(N__33453));
    LocalMux I__6924 (
            .O(N__33471),
            .I(N__33448));
    Sp12to4 I__6923 (
            .O(N__33468),
            .I(N__33448));
    Span4Mux_h I__6922 (
            .O(N__33465),
            .I(N__33445));
    Span4Mux_h I__6921 (
            .O(N__33462),
            .I(N__33442));
    InMux I__6920 (
            .O(N__33461),
            .I(N__33435));
    InMux I__6919 (
            .O(N__33460),
            .I(N__33435));
    InMux I__6918 (
            .O(N__33459),
            .I(N__33435));
    Span12Mux_v I__6917 (
            .O(N__33456),
            .I(N__33428));
    Sp12to4 I__6916 (
            .O(N__33453),
            .I(N__33428));
    Span12Mux_s8_v I__6915 (
            .O(N__33448),
            .I(N__33428));
    Span4Mux_h I__6914 (
            .O(N__33445),
            .I(N__33425));
    Span4Mux_v I__6913 (
            .O(N__33442),
            .I(N__33422));
    LocalMux I__6912 (
            .O(N__33435),
            .I(\c0.FRAME_MATCHER_state_0 ));
    Odrv12 I__6911 (
            .O(N__33428),
            .I(\c0.FRAME_MATCHER_state_0 ));
    Odrv4 I__6910 (
            .O(N__33425),
            .I(\c0.FRAME_MATCHER_state_0 ));
    Odrv4 I__6909 (
            .O(N__33422),
            .I(\c0.FRAME_MATCHER_state_0 ));
    SRMux I__6908 (
            .O(N__33413),
            .I(N__33410));
    LocalMux I__6907 (
            .O(N__33410),
            .I(N__33407));
    Span4Mux_h I__6906 (
            .O(N__33407),
            .I(N__33404));
    Span4Mux_h I__6905 (
            .O(N__33404),
            .I(N__33401));
    Span4Mux_v I__6904 (
            .O(N__33401),
            .I(N__33398));
    Odrv4 I__6903 (
            .O(N__33398),
            .I(\c0.n1_adj_2437 ));
    CascadeMux I__6902 (
            .O(N__33395),
            .I(r_SM_Main_2_N_2323_1_cascade_));
    CascadeMux I__6901 (
            .O(N__33392),
            .I(n17757_cascade_));
    CascadeMux I__6900 (
            .O(N__33389),
            .I(N__33384));
    CascadeMux I__6899 (
            .O(N__33388),
            .I(N__33381));
    InMux I__6898 (
            .O(N__33387),
            .I(N__33375));
    InMux I__6897 (
            .O(N__33384),
            .I(N__33368));
    InMux I__6896 (
            .O(N__33381),
            .I(N__33368));
    InMux I__6895 (
            .O(N__33380),
            .I(N__33368));
    CascadeMux I__6894 (
            .O(N__33379),
            .I(N__33364));
    InMux I__6893 (
            .O(N__33378),
            .I(N__33360));
    LocalMux I__6892 (
            .O(N__33375),
            .I(N__33357));
    LocalMux I__6891 (
            .O(N__33368),
            .I(N__33354));
    CascadeMux I__6890 (
            .O(N__33367),
            .I(N__33351));
    InMux I__6889 (
            .O(N__33364),
            .I(N__33346));
    InMux I__6888 (
            .O(N__33363),
            .I(N__33346));
    LocalMux I__6887 (
            .O(N__33360),
            .I(N__33342));
    Span4Mux_h I__6886 (
            .O(N__33357),
            .I(N__33339));
    Span4Mux_v I__6885 (
            .O(N__33354),
            .I(N__33336));
    InMux I__6884 (
            .O(N__33351),
            .I(N__33333));
    LocalMux I__6883 (
            .O(N__33346),
            .I(N__33330));
    InMux I__6882 (
            .O(N__33345),
            .I(N__33327));
    Sp12to4 I__6881 (
            .O(N__33342),
            .I(N__33323));
    Span4Mux_v I__6880 (
            .O(N__33339),
            .I(N__33317));
    Span4Mux_h I__6879 (
            .O(N__33336),
            .I(N__33312));
    LocalMux I__6878 (
            .O(N__33333),
            .I(N__33312));
    Span4Mux_s3_h I__6877 (
            .O(N__33330),
            .I(N__33307));
    LocalMux I__6876 (
            .O(N__33327),
            .I(N__33307));
    InMux I__6875 (
            .O(N__33326),
            .I(N__33304));
    Span12Mux_v I__6874 (
            .O(N__33323),
            .I(N__33301));
    InMux I__6873 (
            .O(N__33322),
            .I(N__33296));
    InMux I__6872 (
            .O(N__33321),
            .I(N__33296));
    InMux I__6871 (
            .O(N__33320),
            .I(N__33293));
    Span4Mux_v I__6870 (
            .O(N__33317),
            .I(N__33288));
    Span4Mux_v I__6869 (
            .O(N__33312),
            .I(N__33288));
    Span4Mux_v I__6868 (
            .O(N__33307),
            .I(N__33285));
    LocalMux I__6867 (
            .O(N__33304),
            .I(\c0.FRAME_MATCHER_state_2 ));
    Odrv12 I__6866 (
            .O(N__33301),
            .I(\c0.FRAME_MATCHER_state_2 ));
    LocalMux I__6865 (
            .O(N__33296),
            .I(\c0.FRAME_MATCHER_state_2 ));
    LocalMux I__6864 (
            .O(N__33293),
            .I(\c0.FRAME_MATCHER_state_2 ));
    Odrv4 I__6863 (
            .O(N__33288),
            .I(\c0.FRAME_MATCHER_state_2 ));
    Odrv4 I__6862 (
            .O(N__33285),
            .I(\c0.FRAME_MATCHER_state_2 ));
    InMux I__6861 (
            .O(N__33272),
            .I(N__33269));
    LocalMux I__6860 (
            .O(N__33269),
            .I(N__33262));
    InMux I__6859 (
            .O(N__33268),
            .I(N__33255));
    InMux I__6858 (
            .O(N__33267),
            .I(N__33255));
    InMux I__6857 (
            .O(N__33266),
            .I(N__33255));
    InMux I__6856 (
            .O(N__33265),
            .I(N__33252));
    Span4Mux_v I__6855 (
            .O(N__33262),
            .I(N__33246));
    LocalMux I__6854 (
            .O(N__33255),
            .I(N__33243));
    LocalMux I__6853 (
            .O(N__33252),
            .I(N__33238));
    InMux I__6852 (
            .O(N__33251),
            .I(N__33231));
    InMux I__6851 (
            .O(N__33250),
            .I(N__33231));
    InMux I__6850 (
            .O(N__33249),
            .I(N__33231));
    Span4Mux_h I__6849 (
            .O(N__33246),
            .I(N__33226));
    Span4Mux_v I__6848 (
            .O(N__33243),
            .I(N__33223));
    InMux I__6847 (
            .O(N__33242),
            .I(N__33218));
    InMux I__6846 (
            .O(N__33241),
            .I(N__33218));
    Span4Mux_h I__6845 (
            .O(N__33238),
            .I(N__33214));
    LocalMux I__6844 (
            .O(N__33231),
            .I(N__33211));
    InMux I__6843 (
            .O(N__33230),
            .I(N__33208));
    InMux I__6842 (
            .O(N__33229),
            .I(N__33205));
    Span4Mux_v I__6841 (
            .O(N__33226),
            .I(N__33200));
    Span4Mux_h I__6840 (
            .O(N__33223),
            .I(N__33200));
    LocalMux I__6839 (
            .O(N__33218),
            .I(N__33197));
    InMux I__6838 (
            .O(N__33217),
            .I(N__33194));
    Sp12to4 I__6837 (
            .O(N__33214),
            .I(N__33187));
    Sp12to4 I__6836 (
            .O(N__33211),
            .I(N__33187));
    LocalMux I__6835 (
            .O(N__33208),
            .I(N__33187));
    LocalMux I__6834 (
            .O(N__33205),
            .I(N__33182));
    Span4Mux_v I__6833 (
            .O(N__33200),
            .I(N__33182));
    Sp12to4 I__6832 (
            .O(N__33197),
            .I(N__33175));
    LocalMux I__6831 (
            .O(N__33194),
            .I(N__33175));
    Span12Mux_s7_v I__6830 (
            .O(N__33187),
            .I(N__33175));
    Odrv4 I__6829 (
            .O(N__33182),
            .I(\c0.FRAME_MATCHER_state_1 ));
    Odrv12 I__6828 (
            .O(N__33175),
            .I(\c0.FRAME_MATCHER_state_1 ));
    InMux I__6827 (
            .O(N__33170),
            .I(N__33167));
    LocalMux I__6826 (
            .O(N__33167),
            .I(N__33163));
    InMux I__6825 (
            .O(N__33166),
            .I(N__33160));
    Span4Mux_v I__6824 (
            .O(N__33163),
            .I(N__33153));
    LocalMux I__6823 (
            .O(N__33160),
            .I(N__33153));
    InMux I__6822 (
            .O(N__33159),
            .I(N__33150));
    InMux I__6821 (
            .O(N__33158),
            .I(N__33145));
    Span4Mux_h I__6820 (
            .O(N__33153),
            .I(N__33140));
    LocalMux I__6819 (
            .O(N__33150),
            .I(N__33140));
    InMux I__6818 (
            .O(N__33149),
            .I(N__33137));
    CascadeMux I__6817 (
            .O(N__33148),
            .I(N__33134));
    LocalMux I__6816 (
            .O(N__33145),
            .I(N__33131));
    Span4Mux_v I__6815 (
            .O(N__33140),
            .I(N__33126));
    LocalMux I__6814 (
            .O(N__33137),
            .I(N__33126));
    InMux I__6813 (
            .O(N__33134),
            .I(N__33123));
    Span4Mux_h I__6812 (
            .O(N__33131),
            .I(N__33120));
    Span4Mux_h I__6811 (
            .O(N__33126),
            .I(N__33117));
    LocalMux I__6810 (
            .O(N__33123),
            .I(N__33114));
    Span4Mux_v I__6809 (
            .O(N__33120),
            .I(N__33111));
    Span4Mux_h I__6808 (
            .O(N__33117),
            .I(N__33108));
    Span4Mux_h I__6807 (
            .O(N__33114),
            .I(N__33105));
    Odrv4 I__6806 (
            .O(N__33111),
            .I(\c0.n157 ));
    Odrv4 I__6805 (
            .O(N__33108),
            .I(\c0.n157 ));
    Odrv4 I__6804 (
            .O(N__33105),
            .I(\c0.n157 ));
    InMux I__6803 (
            .O(N__33098),
            .I(N__33095));
    LocalMux I__6802 (
            .O(N__33095),
            .I(N__33092));
    Span4Mux_h I__6801 (
            .O(N__33092),
            .I(N__33089));
    Odrv4 I__6800 (
            .O(N__33089),
            .I(n18010));
    InMux I__6799 (
            .O(N__33086),
            .I(N__33083));
    LocalMux I__6798 (
            .O(N__33083),
            .I(N__33080));
    Odrv4 I__6797 (
            .O(N__33080),
            .I(n9390));
    InMux I__6796 (
            .O(N__33077),
            .I(N__33074));
    LocalMux I__6795 (
            .O(N__33074),
            .I(n7364));
    CascadeMux I__6794 (
            .O(N__33071),
            .I(N__33068));
    InMux I__6793 (
            .O(N__33068),
            .I(N__33065));
    LocalMux I__6792 (
            .O(N__33065),
            .I(N__33062));
    Span4Mux_h I__6791 (
            .O(N__33062),
            .I(N__33057));
    InMux I__6790 (
            .O(N__33061),
            .I(N__33054));
    InMux I__6789 (
            .O(N__33060),
            .I(N__33051));
    Span4Mux_v I__6788 (
            .O(N__33057),
            .I(N__33048));
    LocalMux I__6787 (
            .O(N__33054),
            .I(N__33045));
    LocalMux I__6786 (
            .O(N__33051),
            .I(data_in_6_2));
    Odrv4 I__6785 (
            .O(N__33048),
            .I(data_in_6_2));
    Odrv12 I__6784 (
            .O(N__33045),
            .I(data_in_6_2));
    CascadeMux I__6783 (
            .O(N__33038),
            .I(N__33034));
    CascadeMux I__6782 (
            .O(N__33037),
            .I(N__33031));
    InMux I__6781 (
            .O(N__33034),
            .I(N__33028));
    InMux I__6780 (
            .O(N__33031),
            .I(N__33024));
    LocalMux I__6779 (
            .O(N__33028),
            .I(N__33021));
    InMux I__6778 (
            .O(N__33027),
            .I(N__33018));
    LocalMux I__6777 (
            .O(N__33024),
            .I(N__33015));
    Span4Mux_v I__6776 (
            .O(N__33021),
            .I(N__33011));
    LocalMux I__6775 (
            .O(N__33018),
            .I(N__33008));
    Span4Mux_h I__6774 (
            .O(N__33015),
            .I(N__33005));
    InMux I__6773 (
            .O(N__33014),
            .I(N__33002));
    Sp12to4 I__6772 (
            .O(N__33011),
            .I(N__32999));
    Span4Mux_h I__6771 (
            .O(N__33008),
            .I(N__32994));
    Span4Mux_h I__6770 (
            .O(N__33005),
            .I(N__32994));
    LocalMux I__6769 (
            .O(N__33002),
            .I(data_in_5_2));
    Odrv12 I__6768 (
            .O(N__32999),
            .I(data_in_5_2));
    Odrv4 I__6767 (
            .O(N__32994),
            .I(data_in_5_2));
    InMux I__6766 (
            .O(N__32987),
            .I(N__32980));
    CascadeMux I__6765 (
            .O(N__32986),
            .I(N__32977));
    InMux I__6764 (
            .O(N__32985),
            .I(N__32974));
    InMux I__6763 (
            .O(N__32984),
            .I(N__32971));
    InMux I__6762 (
            .O(N__32983),
            .I(N__32968));
    LocalMux I__6761 (
            .O(N__32980),
            .I(N__32965));
    InMux I__6760 (
            .O(N__32977),
            .I(N__32962));
    LocalMux I__6759 (
            .O(N__32974),
            .I(N__32957));
    LocalMux I__6758 (
            .O(N__32971),
            .I(N__32957));
    LocalMux I__6757 (
            .O(N__32968),
            .I(N__32952));
    Span4Mux_v I__6756 (
            .O(N__32965),
            .I(N__32952));
    LocalMux I__6755 (
            .O(N__32962),
            .I(N__32949));
    Span4Mux_v I__6754 (
            .O(N__32957),
            .I(N__32946));
    Span4Mux_v I__6753 (
            .O(N__32952),
            .I(N__32941));
    Span4Mux_h I__6752 (
            .O(N__32949),
            .I(N__32941));
    Odrv4 I__6751 (
            .O(N__32946),
            .I(\c0.data_in_frame_10_5 ));
    Odrv4 I__6750 (
            .O(N__32941),
            .I(\c0.data_in_frame_10_5 ));
    InMux I__6749 (
            .O(N__32936),
            .I(N__32932));
    InMux I__6748 (
            .O(N__32935),
            .I(N__32929));
    LocalMux I__6747 (
            .O(N__32932),
            .I(N__32924));
    LocalMux I__6746 (
            .O(N__32929),
            .I(N__32924));
    Odrv12 I__6745 (
            .O(N__32924),
            .I(n2562));
    InMux I__6744 (
            .O(N__32921),
            .I(N__32912));
    InMux I__6743 (
            .O(N__32920),
            .I(N__32912));
    InMux I__6742 (
            .O(N__32919),
            .I(N__32912));
    LocalMux I__6741 (
            .O(N__32912),
            .I(data_in_10_5));
    InMux I__6740 (
            .O(N__32909),
            .I(N__32905));
    InMux I__6739 (
            .O(N__32908),
            .I(N__32902));
    LocalMux I__6738 (
            .O(N__32905),
            .I(N__32899));
    LocalMux I__6737 (
            .O(N__32902),
            .I(N__32896));
    Span4Mux_h I__6736 (
            .O(N__32899),
            .I(N__32893));
    Span4Mux_v I__6735 (
            .O(N__32896),
            .I(N__32889));
    Span4Mux_h I__6734 (
            .O(N__32893),
            .I(N__32886));
    InMux I__6733 (
            .O(N__32892),
            .I(N__32883));
    Span4Mux_h I__6732 (
            .O(N__32889),
            .I(N__32880));
    Odrv4 I__6731 (
            .O(N__32886),
            .I(data_in_9_5));
    LocalMux I__6730 (
            .O(N__32883),
            .I(data_in_9_5));
    Odrv4 I__6729 (
            .O(N__32880),
            .I(data_in_9_5));
    InMux I__6728 (
            .O(N__32873),
            .I(N__32870));
    LocalMux I__6727 (
            .O(N__32870),
            .I(N__32866));
    InMux I__6726 (
            .O(N__32869),
            .I(N__32863));
    Odrv4 I__6725 (
            .O(N__32866),
            .I(data_in_12_5));
    LocalMux I__6724 (
            .O(N__32863),
            .I(data_in_12_5));
    InMux I__6723 (
            .O(N__32858),
            .I(N__32852));
    InMux I__6722 (
            .O(N__32857),
            .I(N__32852));
    LocalMux I__6721 (
            .O(N__32852),
            .I(data_in_11_5));
    InMux I__6720 (
            .O(N__32849),
            .I(N__32846));
    LocalMux I__6719 (
            .O(N__32846),
            .I(n18098));
    InMux I__6718 (
            .O(N__32843),
            .I(N__32838));
    CascadeMux I__6717 (
            .O(N__32842),
            .I(N__32835));
    CEMux I__6716 (
            .O(N__32841),
            .I(N__32829));
    LocalMux I__6715 (
            .O(N__32838),
            .I(N__32806));
    InMux I__6714 (
            .O(N__32835),
            .I(N__32801));
    InMux I__6713 (
            .O(N__32834),
            .I(N__32801));
    InMux I__6712 (
            .O(N__32833),
            .I(N__32793));
    InMux I__6711 (
            .O(N__32832),
            .I(N__32784));
    LocalMux I__6710 (
            .O(N__32829),
            .I(N__32781));
    CEMux I__6709 (
            .O(N__32828),
            .I(N__32778));
    InMux I__6708 (
            .O(N__32827),
            .I(N__32775));
    CascadeMux I__6707 (
            .O(N__32826),
            .I(N__32772));
    CascadeMux I__6706 (
            .O(N__32825),
            .I(N__32768));
    CascadeMux I__6705 (
            .O(N__32824),
            .I(N__32765));
    InMux I__6704 (
            .O(N__32823),
            .I(N__32738));
    InMux I__6703 (
            .O(N__32822),
            .I(N__32738));
    InMux I__6702 (
            .O(N__32821),
            .I(N__32729));
    InMux I__6701 (
            .O(N__32820),
            .I(N__32729));
    InMux I__6700 (
            .O(N__32819),
            .I(N__32729));
    InMux I__6699 (
            .O(N__32818),
            .I(N__32729));
    InMux I__6698 (
            .O(N__32817),
            .I(N__32724));
    InMux I__6697 (
            .O(N__32816),
            .I(N__32724));
    InMux I__6696 (
            .O(N__32815),
            .I(N__32712));
    CEMux I__6695 (
            .O(N__32814),
            .I(N__32709));
    InMux I__6694 (
            .O(N__32813),
            .I(N__32706));
    InMux I__6693 (
            .O(N__32812),
            .I(N__32699));
    InMux I__6692 (
            .O(N__32811),
            .I(N__32699));
    InMux I__6691 (
            .O(N__32810),
            .I(N__32699));
    InMux I__6690 (
            .O(N__32809),
            .I(N__32696));
    Span4Mux_h I__6689 (
            .O(N__32806),
            .I(N__32691));
    LocalMux I__6688 (
            .O(N__32801),
            .I(N__32691));
    InMux I__6687 (
            .O(N__32800),
            .I(N__32682));
    InMux I__6686 (
            .O(N__32799),
            .I(N__32682));
    InMux I__6685 (
            .O(N__32798),
            .I(N__32682));
    InMux I__6684 (
            .O(N__32797),
            .I(N__32682));
    InMux I__6683 (
            .O(N__32796),
            .I(N__32679));
    LocalMux I__6682 (
            .O(N__32793),
            .I(N__32675));
    CEMux I__6681 (
            .O(N__32792),
            .I(N__32672));
    InMux I__6680 (
            .O(N__32791),
            .I(N__32661));
    InMux I__6679 (
            .O(N__32790),
            .I(N__32661));
    InMux I__6678 (
            .O(N__32789),
            .I(N__32661));
    InMux I__6677 (
            .O(N__32788),
            .I(N__32661));
    InMux I__6676 (
            .O(N__32787),
            .I(N__32661));
    LocalMux I__6675 (
            .O(N__32784),
            .I(N__32656));
    Span4Mux_v I__6674 (
            .O(N__32781),
            .I(N__32656));
    LocalMux I__6673 (
            .O(N__32778),
            .I(N__32653));
    LocalMux I__6672 (
            .O(N__32775),
            .I(N__32644));
    InMux I__6671 (
            .O(N__32772),
            .I(N__32640));
    CEMux I__6670 (
            .O(N__32771),
            .I(N__32595));
    InMux I__6669 (
            .O(N__32768),
            .I(N__32588));
    InMux I__6668 (
            .O(N__32765),
            .I(N__32588));
    InMux I__6667 (
            .O(N__32764),
            .I(N__32588));
    InMux I__6666 (
            .O(N__32763),
            .I(N__32581));
    InMux I__6665 (
            .O(N__32762),
            .I(N__32581));
    InMux I__6664 (
            .O(N__32761),
            .I(N__32581));
    InMux I__6663 (
            .O(N__32760),
            .I(N__32566));
    InMux I__6662 (
            .O(N__32759),
            .I(N__32566));
    InMux I__6661 (
            .O(N__32758),
            .I(N__32566));
    InMux I__6660 (
            .O(N__32757),
            .I(N__32566));
    InMux I__6659 (
            .O(N__32756),
            .I(N__32566));
    InMux I__6658 (
            .O(N__32755),
            .I(N__32566));
    InMux I__6657 (
            .O(N__32754),
            .I(N__32566));
    InMux I__6656 (
            .O(N__32753),
            .I(N__32549));
    InMux I__6655 (
            .O(N__32752),
            .I(N__32549));
    InMux I__6654 (
            .O(N__32751),
            .I(N__32549));
    InMux I__6653 (
            .O(N__32750),
            .I(N__32549));
    InMux I__6652 (
            .O(N__32749),
            .I(N__32549));
    InMux I__6651 (
            .O(N__32748),
            .I(N__32549));
    InMux I__6650 (
            .O(N__32747),
            .I(N__32549));
    InMux I__6649 (
            .O(N__32746),
            .I(N__32549));
    InMux I__6648 (
            .O(N__32745),
            .I(N__32542));
    InMux I__6647 (
            .O(N__32744),
            .I(N__32542));
    InMux I__6646 (
            .O(N__32743),
            .I(N__32542));
    LocalMux I__6645 (
            .O(N__32738),
            .I(N__32539));
    LocalMux I__6644 (
            .O(N__32729),
            .I(N__32536));
    LocalMux I__6643 (
            .O(N__32724),
            .I(N__32533));
    InMux I__6642 (
            .O(N__32723),
            .I(N__32526));
    InMux I__6641 (
            .O(N__32722),
            .I(N__32526));
    InMux I__6640 (
            .O(N__32721),
            .I(N__32526));
    InMux I__6639 (
            .O(N__32720),
            .I(N__32513));
    InMux I__6638 (
            .O(N__32719),
            .I(N__32513));
    InMux I__6637 (
            .O(N__32718),
            .I(N__32513));
    InMux I__6636 (
            .O(N__32717),
            .I(N__32513));
    InMux I__6635 (
            .O(N__32716),
            .I(N__32513));
    InMux I__6634 (
            .O(N__32715),
            .I(N__32513));
    LocalMux I__6633 (
            .O(N__32712),
            .I(N__32508));
    LocalMux I__6632 (
            .O(N__32709),
            .I(N__32508));
    LocalMux I__6631 (
            .O(N__32706),
            .I(N__32497));
    LocalMux I__6630 (
            .O(N__32699),
            .I(N__32497));
    LocalMux I__6629 (
            .O(N__32696),
            .I(N__32497));
    Span4Mux_h I__6628 (
            .O(N__32691),
            .I(N__32497));
    LocalMux I__6627 (
            .O(N__32682),
            .I(N__32497));
    LocalMux I__6626 (
            .O(N__32679),
            .I(N__32494));
    InMux I__6625 (
            .O(N__32678),
            .I(N__32491));
    Span4Mux_h I__6624 (
            .O(N__32675),
            .I(N__32488));
    LocalMux I__6623 (
            .O(N__32672),
            .I(N__32485));
    LocalMux I__6622 (
            .O(N__32661),
            .I(N__32478));
    Span4Mux_h I__6621 (
            .O(N__32656),
            .I(N__32478));
    Span4Mux_v I__6620 (
            .O(N__32653),
            .I(N__32478));
    InMux I__6619 (
            .O(N__32652),
            .I(N__32475));
    InMux I__6618 (
            .O(N__32651),
            .I(N__32464));
    InMux I__6617 (
            .O(N__32650),
            .I(N__32464));
    InMux I__6616 (
            .O(N__32649),
            .I(N__32464));
    InMux I__6615 (
            .O(N__32648),
            .I(N__32464));
    InMux I__6614 (
            .O(N__32647),
            .I(N__32464));
    Sp12to4 I__6613 (
            .O(N__32644),
            .I(N__32461));
    InMux I__6612 (
            .O(N__32643),
            .I(N__32458));
    LocalMux I__6611 (
            .O(N__32640),
            .I(N__32455));
    InMux I__6610 (
            .O(N__32639),
            .I(N__32438));
    InMux I__6609 (
            .O(N__32638),
            .I(N__32438));
    InMux I__6608 (
            .O(N__32637),
            .I(N__32438));
    InMux I__6607 (
            .O(N__32636),
            .I(N__32438));
    InMux I__6606 (
            .O(N__32635),
            .I(N__32438));
    InMux I__6605 (
            .O(N__32634),
            .I(N__32438));
    InMux I__6604 (
            .O(N__32633),
            .I(N__32438));
    InMux I__6603 (
            .O(N__32632),
            .I(N__32438));
    InMux I__6602 (
            .O(N__32631),
            .I(N__32421));
    InMux I__6601 (
            .O(N__32630),
            .I(N__32421));
    InMux I__6600 (
            .O(N__32629),
            .I(N__32421));
    InMux I__6599 (
            .O(N__32628),
            .I(N__32421));
    InMux I__6598 (
            .O(N__32627),
            .I(N__32421));
    InMux I__6597 (
            .O(N__32626),
            .I(N__32421));
    InMux I__6596 (
            .O(N__32625),
            .I(N__32421));
    InMux I__6595 (
            .O(N__32624),
            .I(N__32421));
    InMux I__6594 (
            .O(N__32623),
            .I(N__32404));
    InMux I__6593 (
            .O(N__32622),
            .I(N__32404));
    InMux I__6592 (
            .O(N__32621),
            .I(N__32404));
    InMux I__6591 (
            .O(N__32620),
            .I(N__32404));
    InMux I__6590 (
            .O(N__32619),
            .I(N__32404));
    InMux I__6589 (
            .O(N__32618),
            .I(N__32404));
    InMux I__6588 (
            .O(N__32617),
            .I(N__32404));
    InMux I__6587 (
            .O(N__32616),
            .I(N__32404));
    InMux I__6586 (
            .O(N__32615),
            .I(N__32387));
    InMux I__6585 (
            .O(N__32614),
            .I(N__32387));
    InMux I__6584 (
            .O(N__32613),
            .I(N__32387));
    InMux I__6583 (
            .O(N__32612),
            .I(N__32387));
    InMux I__6582 (
            .O(N__32611),
            .I(N__32387));
    InMux I__6581 (
            .O(N__32610),
            .I(N__32387));
    InMux I__6580 (
            .O(N__32609),
            .I(N__32387));
    InMux I__6579 (
            .O(N__32608),
            .I(N__32387));
    InMux I__6578 (
            .O(N__32607),
            .I(N__32372));
    InMux I__6577 (
            .O(N__32606),
            .I(N__32372));
    InMux I__6576 (
            .O(N__32605),
            .I(N__32372));
    InMux I__6575 (
            .O(N__32604),
            .I(N__32372));
    InMux I__6574 (
            .O(N__32603),
            .I(N__32372));
    InMux I__6573 (
            .O(N__32602),
            .I(N__32372));
    InMux I__6572 (
            .O(N__32601),
            .I(N__32372));
    InMux I__6571 (
            .O(N__32600),
            .I(N__32365));
    InMux I__6570 (
            .O(N__32599),
            .I(N__32365));
    InMux I__6569 (
            .O(N__32598),
            .I(N__32365));
    LocalMux I__6568 (
            .O(N__32595),
            .I(N__32360));
    LocalMux I__6567 (
            .O(N__32588),
            .I(N__32360));
    LocalMux I__6566 (
            .O(N__32581),
            .I(N__32345));
    LocalMux I__6565 (
            .O(N__32566),
            .I(N__32345));
    LocalMux I__6564 (
            .O(N__32549),
            .I(N__32345));
    LocalMux I__6563 (
            .O(N__32542),
            .I(N__32345));
    Span4Mux_h I__6562 (
            .O(N__32539),
            .I(N__32345));
    Span4Mux_v I__6561 (
            .O(N__32536),
            .I(N__32345));
    Span4Mux_v I__6560 (
            .O(N__32533),
            .I(N__32345));
    LocalMux I__6559 (
            .O(N__32526),
            .I(N__32334));
    LocalMux I__6558 (
            .O(N__32513),
            .I(N__32334));
    Span4Mux_h I__6557 (
            .O(N__32508),
            .I(N__32334));
    Span4Mux_v I__6556 (
            .O(N__32497),
            .I(N__32334));
    Span4Mux_s2_h I__6555 (
            .O(N__32494),
            .I(N__32334));
    LocalMux I__6554 (
            .O(N__32491),
            .I(N__32329));
    Span4Mux_s3_h I__6553 (
            .O(N__32488),
            .I(N__32329));
    Span4Mux_v I__6552 (
            .O(N__32485),
            .I(N__32324));
    Span4Mux_v I__6551 (
            .O(N__32478),
            .I(N__32324));
    LocalMux I__6550 (
            .O(N__32475),
            .I(N__32317));
    LocalMux I__6549 (
            .O(N__32464),
            .I(N__32317));
    Span12Mux_v I__6548 (
            .O(N__32461),
            .I(N__32317));
    LocalMux I__6547 (
            .O(N__32458),
            .I(N__32312));
    Span12Mux_v I__6546 (
            .O(N__32455),
            .I(N__32312));
    LocalMux I__6545 (
            .O(N__32438),
            .I(n9606));
    LocalMux I__6544 (
            .O(N__32421),
            .I(n9606));
    LocalMux I__6543 (
            .O(N__32404),
            .I(n9606));
    LocalMux I__6542 (
            .O(N__32387),
            .I(n9606));
    LocalMux I__6541 (
            .O(N__32372),
            .I(n9606));
    LocalMux I__6540 (
            .O(N__32365),
            .I(n9606));
    Odrv4 I__6539 (
            .O(N__32360),
            .I(n9606));
    Odrv4 I__6538 (
            .O(N__32345),
            .I(n9606));
    Odrv4 I__6537 (
            .O(N__32334),
            .I(n9606));
    Odrv4 I__6536 (
            .O(N__32329),
            .I(n9606));
    Odrv4 I__6535 (
            .O(N__32324),
            .I(n9606));
    Odrv12 I__6534 (
            .O(N__32317),
            .I(n9606));
    Odrv12 I__6533 (
            .O(N__32312),
            .I(n9606));
    InMux I__6532 (
            .O(N__32285),
            .I(N__32282));
    LocalMux I__6531 (
            .O(N__32282),
            .I(N__32279));
    Span4Mux_h I__6530 (
            .O(N__32279),
            .I(N__32275));
    InMux I__6529 (
            .O(N__32278),
            .I(N__32272));
    Span4Mux_h I__6528 (
            .O(N__32275),
            .I(N__32269));
    LocalMux I__6527 (
            .O(N__32272),
            .I(data_out_frame2_7_7));
    Odrv4 I__6526 (
            .O(N__32269),
            .I(data_out_frame2_7_7));
    InMux I__6525 (
            .O(N__32264),
            .I(N__32260));
    CascadeMux I__6524 (
            .O(N__32263),
            .I(N__32257));
    LocalMux I__6523 (
            .O(N__32260),
            .I(N__32253));
    InMux I__6522 (
            .O(N__32257),
            .I(N__32250));
    InMux I__6521 (
            .O(N__32256),
            .I(N__32247));
    Span4Mux_v I__6520 (
            .O(N__32253),
            .I(N__32241));
    LocalMux I__6519 (
            .O(N__32250),
            .I(N__32241));
    LocalMux I__6518 (
            .O(N__32247),
            .I(N__32238));
    InMux I__6517 (
            .O(N__32246),
            .I(N__32235));
    Sp12to4 I__6516 (
            .O(N__32241),
            .I(N__32232));
    Span4Mux_s3_h I__6515 (
            .O(N__32238),
            .I(N__32229));
    LocalMux I__6514 (
            .O(N__32235),
            .I(N__32226));
    Span12Mux_s11_v I__6513 (
            .O(N__32232),
            .I(N__32223));
    Odrv4 I__6512 (
            .O(N__32229),
            .I(\c0.data_in_frame_9_7 ));
    Odrv12 I__6511 (
            .O(N__32226),
            .I(\c0.data_in_frame_9_7 ));
    Odrv12 I__6510 (
            .O(N__32223),
            .I(\c0.data_in_frame_9_7 ));
    InMux I__6509 (
            .O(N__32216),
            .I(N__32208));
    InMux I__6508 (
            .O(N__32215),
            .I(N__32208));
    InMux I__6507 (
            .O(N__32214),
            .I(N__32205));
    InMux I__6506 (
            .O(N__32213),
            .I(N__32202));
    LocalMux I__6505 (
            .O(N__32208),
            .I(N__32199));
    LocalMux I__6504 (
            .O(N__32205),
            .I(N__32196));
    LocalMux I__6503 (
            .O(N__32202),
            .I(N__32193));
    Span4Mux_h I__6502 (
            .O(N__32199),
            .I(N__32190));
    Span4Mux_v I__6501 (
            .O(N__32196),
            .I(N__32187));
    Span4Mux_h I__6500 (
            .O(N__32193),
            .I(N__32184));
    Span4Mux_h I__6499 (
            .O(N__32190),
            .I(N__32181));
    Span4Mux_h I__6498 (
            .O(N__32187),
            .I(N__32178));
    Span4Mux_h I__6497 (
            .O(N__32184),
            .I(N__32175));
    Sp12to4 I__6496 (
            .O(N__32181),
            .I(N__32172));
    Odrv4 I__6495 (
            .O(N__32178),
            .I(\c0.n17433 ));
    Odrv4 I__6494 (
            .O(N__32175),
            .I(\c0.n17433 ));
    Odrv12 I__6493 (
            .O(N__32172),
            .I(\c0.n17433 ));
    InMux I__6492 (
            .O(N__32165),
            .I(N__32162));
    LocalMux I__6491 (
            .O(N__32162),
            .I(N__32158));
    CascadeMux I__6490 (
            .O(N__32161),
            .I(N__32155));
    Span4Mux_v I__6489 (
            .O(N__32158),
            .I(N__32152));
    InMux I__6488 (
            .O(N__32155),
            .I(N__32149));
    Span4Mux_h I__6487 (
            .O(N__32152),
            .I(N__32144));
    LocalMux I__6486 (
            .O(N__32149),
            .I(N__32144));
    Span4Mux_h I__6485 (
            .O(N__32144),
            .I(N__32141));
    Span4Mux_s1_h I__6484 (
            .O(N__32141),
            .I(N__32137));
    InMux I__6483 (
            .O(N__32140),
            .I(N__32134));
    Span4Mux_v I__6482 (
            .O(N__32137),
            .I(N__32131));
    LocalMux I__6481 (
            .O(N__32134),
            .I(data_in_7_7));
    Odrv4 I__6480 (
            .O(N__32131),
            .I(data_in_7_7));
    InMux I__6479 (
            .O(N__32126),
            .I(N__32123));
    LocalMux I__6478 (
            .O(N__32123),
            .I(N__32120));
    Span4Mux_v I__6477 (
            .O(N__32120),
            .I(N__32117));
    Odrv4 I__6476 (
            .O(N__32117),
            .I(n2573));
    InMux I__6475 (
            .O(N__32114),
            .I(N__32111));
    LocalMux I__6474 (
            .O(N__32111),
            .I(N__32107));
    InMux I__6473 (
            .O(N__32110),
            .I(N__32103));
    Span4Mux_h I__6472 (
            .O(N__32107),
            .I(N__32100));
    InMux I__6471 (
            .O(N__32106),
            .I(N__32097));
    LocalMux I__6470 (
            .O(N__32103),
            .I(N__32094));
    Span4Mux_v I__6469 (
            .O(N__32100),
            .I(N__32089));
    LocalMux I__6468 (
            .O(N__32097),
            .I(N__32089));
    Span4Mux_v I__6467 (
            .O(N__32094),
            .I(N__32084));
    Span4Mux_v I__6466 (
            .O(N__32089),
            .I(N__32084));
    Sp12to4 I__6465 (
            .O(N__32084),
            .I(N__32081));
    Odrv12 I__6464 (
            .O(N__32081),
            .I(\c0.data_in_frame_9_2 ));
    InMux I__6463 (
            .O(N__32078),
            .I(N__32075));
    LocalMux I__6462 (
            .O(N__32075),
            .I(N__32072));
    Span4Mux_h I__6461 (
            .O(N__32072),
            .I(N__32069));
    Odrv4 I__6460 (
            .O(N__32069),
            .I(n2565));
    InMux I__6459 (
            .O(N__32066),
            .I(N__32061));
    InMux I__6458 (
            .O(N__32065),
            .I(N__32058));
    InMux I__6457 (
            .O(N__32064),
            .I(N__32054));
    LocalMux I__6456 (
            .O(N__32061),
            .I(N__32049));
    LocalMux I__6455 (
            .O(N__32058),
            .I(N__32049));
    CascadeMux I__6454 (
            .O(N__32057),
            .I(N__32046));
    LocalMux I__6453 (
            .O(N__32054),
            .I(N__32042));
    Span4Mux_h I__6452 (
            .O(N__32049),
            .I(N__32039));
    InMux I__6451 (
            .O(N__32046),
            .I(N__32036));
    InMux I__6450 (
            .O(N__32045),
            .I(N__32033));
    Span4Mux_h I__6449 (
            .O(N__32042),
            .I(N__32026));
    Span4Mux_v I__6448 (
            .O(N__32039),
            .I(N__32026));
    LocalMux I__6447 (
            .O(N__32036),
            .I(N__32026));
    LocalMux I__6446 (
            .O(N__32033),
            .I(N__32023));
    Span4Mux_v I__6445 (
            .O(N__32026),
            .I(N__32020));
    Span12Mux_s8_h I__6444 (
            .O(N__32023),
            .I(N__32017));
    Sp12to4 I__6443 (
            .O(N__32020),
            .I(N__32014));
    Odrv12 I__6442 (
            .O(N__32017),
            .I(\c0.data_in_frame_10_2 ));
    Odrv12 I__6441 (
            .O(N__32014),
            .I(\c0.data_in_frame_10_2 ));
    InMux I__6440 (
            .O(N__32009),
            .I(N__32006));
    LocalMux I__6439 (
            .O(N__32006),
            .I(N__32003));
    Span4Mux_v I__6438 (
            .O(N__32003),
            .I(N__32000));
    Odrv4 I__6437 (
            .O(N__32000),
            .I(n2566));
    CascadeMux I__6436 (
            .O(N__31997),
            .I(N__31989));
    CascadeMux I__6435 (
            .O(N__31996),
            .I(N__31985));
    CascadeMux I__6434 (
            .O(N__31995),
            .I(N__31982));
    InMux I__6433 (
            .O(N__31994),
            .I(N__31959));
    InMux I__6432 (
            .O(N__31993),
            .I(N__31959));
    InMux I__6431 (
            .O(N__31992),
            .I(N__31959));
    InMux I__6430 (
            .O(N__31989),
            .I(N__31959));
    InMux I__6429 (
            .O(N__31988),
            .I(N__31952));
    InMux I__6428 (
            .O(N__31985),
            .I(N__31952));
    InMux I__6427 (
            .O(N__31982),
            .I(N__31952));
    CascadeMux I__6426 (
            .O(N__31981),
            .I(N__31947));
    CascadeMux I__6425 (
            .O(N__31980),
            .I(N__31944));
    InMux I__6424 (
            .O(N__31979),
            .I(N__31938));
    CascadeMux I__6423 (
            .O(N__31978),
            .I(N__31934));
    InMux I__6422 (
            .O(N__31977),
            .I(N__31929));
    InMux I__6421 (
            .O(N__31976),
            .I(N__31929));
    InMux I__6420 (
            .O(N__31975),
            .I(N__31914));
    InMux I__6419 (
            .O(N__31974),
            .I(N__31911));
    InMux I__6418 (
            .O(N__31973),
            .I(N__31908));
    InMux I__6417 (
            .O(N__31972),
            .I(N__31903));
    InMux I__6416 (
            .O(N__31971),
            .I(N__31894));
    InMux I__6415 (
            .O(N__31970),
            .I(N__31894));
    InMux I__6414 (
            .O(N__31969),
            .I(N__31894));
    InMux I__6413 (
            .O(N__31968),
            .I(N__31894));
    LocalMux I__6412 (
            .O(N__31959),
            .I(N__31887));
    LocalMux I__6411 (
            .O(N__31952),
            .I(N__31887));
    InMux I__6410 (
            .O(N__31951),
            .I(N__31878));
    InMux I__6409 (
            .O(N__31950),
            .I(N__31878));
    InMux I__6408 (
            .O(N__31947),
            .I(N__31878));
    InMux I__6407 (
            .O(N__31944),
            .I(N__31878));
    CascadeMux I__6406 (
            .O(N__31943),
            .I(N__31872));
    CascadeMux I__6405 (
            .O(N__31942),
            .I(N__31867));
    CascadeMux I__6404 (
            .O(N__31941),
            .I(N__31864));
    LocalMux I__6403 (
            .O(N__31938),
            .I(N__31861));
    InMux I__6402 (
            .O(N__31937),
            .I(N__31856));
    InMux I__6401 (
            .O(N__31934),
            .I(N__31856));
    LocalMux I__6400 (
            .O(N__31929),
            .I(N__31853));
    CascadeMux I__6399 (
            .O(N__31928),
            .I(N__31844));
    CascadeMux I__6398 (
            .O(N__31927),
            .I(N__31841));
    CascadeMux I__6397 (
            .O(N__31926),
            .I(N__31835));
    CascadeMux I__6396 (
            .O(N__31925),
            .I(N__31832));
    CascadeMux I__6395 (
            .O(N__31924),
            .I(N__31825));
    CascadeMux I__6394 (
            .O(N__31923),
            .I(N__31813));
    CascadeMux I__6393 (
            .O(N__31922),
            .I(N__31810));
    CascadeMux I__6392 (
            .O(N__31921),
            .I(N__31800));
    CascadeMux I__6391 (
            .O(N__31920),
            .I(N__31792));
    InMux I__6390 (
            .O(N__31919),
            .I(N__31786));
    InMux I__6389 (
            .O(N__31918),
            .I(N__31783));
    InMux I__6388 (
            .O(N__31917),
            .I(N__31780));
    LocalMux I__6387 (
            .O(N__31914),
            .I(N__31777));
    LocalMux I__6386 (
            .O(N__31911),
            .I(N__31774));
    LocalMux I__6385 (
            .O(N__31908),
            .I(N__31771));
    InMux I__6384 (
            .O(N__31907),
            .I(N__31768));
    InMux I__6383 (
            .O(N__31906),
            .I(N__31765));
    LocalMux I__6382 (
            .O(N__31903),
            .I(N__31760));
    LocalMux I__6381 (
            .O(N__31894),
            .I(N__31760));
    InMux I__6380 (
            .O(N__31893),
            .I(N__31755));
    InMux I__6379 (
            .O(N__31892),
            .I(N__31755));
    Span4Mux_h I__6378 (
            .O(N__31887),
            .I(N__31750));
    LocalMux I__6377 (
            .O(N__31878),
            .I(N__31750));
    InMux I__6376 (
            .O(N__31877),
            .I(N__31747));
    InMux I__6375 (
            .O(N__31876),
            .I(N__31740));
    InMux I__6374 (
            .O(N__31875),
            .I(N__31740));
    InMux I__6373 (
            .O(N__31872),
            .I(N__31740));
    InMux I__6372 (
            .O(N__31871),
            .I(N__31731));
    InMux I__6371 (
            .O(N__31870),
            .I(N__31731));
    InMux I__6370 (
            .O(N__31867),
            .I(N__31731));
    InMux I__6369 (
            .O(N__31864),
            .I(N__31731));
    Span4Mux_s3_h I__6368 (
            .O(N__31861),
            .I(N__31724));
    LocalMux I__6367 (
            .O(N__31856),
            .I(N__31724));
    Span4Mux_s3_h I__6366 (
            .O(N__31853),
            .I(N__31724));
    CascadeMux I__6365 (
            .O(N__31852),
            .I(N__31720));
    CascadeMux I__6364 (
            .O(N__31851),
            .I(N__31717));
    CascadeMux I__6363 (
            .O(N__31850),
            .I(N__31714));
    InMux I__6362 (
            .O(N__31849),
            .I(N__31701));
    InMux I__6361 (
            .O(N__31848),
            .I(N__31701));
    InMux I__6360 (
            .O(N__31847),
            .I(N__31701));
    InMux I__6359 (
            .O(N__31844),
            .I(N__31701));
    InMux I__6358 (
            .O(N__31841),
            .I(N__31701));
    InMux I__6357 (
            .O(N__31840),
            .I(N__31686));
    InMux I__6356 (
            .O(N__31839),
            .I(N__31686));
    InMux I__6355 (
            .O(N__31838),
            .I(N__31686));
    InMux I__6354 (
            .O(N__31835),
            .I(N__31686));
    InMux I__6353 (
            .O(N__31832),
            .I(N__31686));
    InMux I__6352 (
            .O(N__31831),
            .I(N__31686));
    InMux I__6351 (
            .O(N__31830),
            .I(N__31686));
    InMux I__6350 (
            .O(N__31829),
            .I(N__31675));
    InMux I__6349 (
            .O(N__31828),
            .I(N__31675));
    InMux I__6348 (
            .O(N__31825),
            .I(N__31675));
    InMux I__6347 (
            .O(N__31824),
            .I(N__31675));
    InMux I__6346 (
            .O(N__31823),
            .I(N__31675));
    InMux I__6345 (
            .O(N__31822),
            .I(N__31664));
    InMux I__6344 (
            .O(N__31821),
            .I(N__31664));
    InMux I__6343 (
            .O(N__31820),
            .I(N__31664));
    InMux I__6342 (
            .O(N__31819),
            .I(N__31664));
    InMux I__6341 (
            .O(N__31818),
            .I(N__31664));
    InMux I__6340 (
            .O(N__31817),
            .I(N__31655));
    InMux I__6339 (
            .O(N__31816),
            .I(N__31655));
    InMux I__6338 (
            .O(N__31813),
            .I(N__31655));
    InMux I__6337 (
            .O(N__31810),
            .I(N__31655));
    InMux I__6336 (
            .O(N__31809),
            .I(N__31642));
    InMux I__6335 (
            .O(N__31808),
            .I(N__31642));
    InMux I__6334 (
            .O(N__31807),
            .I(N__31642));
    InMux I__6333 (
            .O(N__31806),
            .I(N__31642));
    InMux I__6332 (
            .O(N__31805),
            .I(N__31642));
    InMux I__6331 (
            .O(N__31804),
            .I(N__31642));
    InMux I__6330 (
            .O(N__31803),
            .I(N__31631));
    InMux I__6329 (
            .O(N__31800),
            .I(N__31631));
    InMux I__6328 (
            .O(N__31799),
            .I(N__31631));
    InMux I__6327 (
            .O(N__31798),
            .I(N__31631));
    InMux I__6326 (
            .O(N__31797),
            .I(N__31631));
    InMux I__6325 (
            .O(N__31796),
            .I(N__31618));
    InMux I__6324 (
            .O(N__31795),
            .I(N__31618));
    InMux I__6323 (
            .O(N__31792),
            .I(N__31618));
    InMux I__6322 (
            .O(N__31791),
            .I(N__31618));
    InMux I__6321 (
            .O(N__31790),
            .I(N__31618));
    InMux I__6320 (
            .O(N__31789),
            .I(N__31618));
    LocalMux I__6319 (
            .O(N__31786),
            .I(N__31615));
    LocalMux I__6318 (
            .O(N__31783),
            .I(N__31604));
    LocalMux I__6317 (
            .O(N__31780),
            .I(N__31604));
    Span4Mux_v I__6316 (
            .O(N__31777),
            .I(N__31604));
    Span4Mux_v I__6315 (
            .O(N__31774),
            .I(N__31604));
    Span4Mux_v I__6314 (
            .O(N__31771),
            .I(N__31604));
    LocalMux I__6313 (
            .O(N__31768),
            .I(N__31597));
    LocalMux I__6312 (
            .O(N__31765),
            .I(N__31597));
    Span4Mux_h I__6311 (
            .O(N__31760),
            .I(N__31597));
    LocalMux I__6310 (
            .O(N__31755),
            .I(N__31592));
    Span4Mux_s3_h I__6309 (
            .O(N__31750),
            .I(N__31592));
    LocalMux I__6308 (
            .O(N__31747),
            .I(N__31583));
    LocalMux I__6307 (
            .O(N__31740),
            .I(N__31583));
    LocalMux I__6306 (
            .O(N__31731),
            .I(N__31583));
    Span4Mux_h I__6305 (
            .O(N__31724),
            .I(N__31583));
    InMux I__6304 (
            .O(N__31723),
            .I(N__31570));
    InMux I__6303 (
            .O(N__31720),
            .I(N__31570));
    InMux I__6302 (
            .O(N__31717),
            .I(N__31570));
    InMux I__6301 (
            .O(N__31714),
            .I(N__31570));
    InMux I__6300 (
            .O(N__31713),
            .I(N__31570));
    InMux I__6299 (
            .O(N__31712),
            .I(N__31570));
    LocalMux I__6298 (
            .O(N__31701),
            .I(n1396));
    LocalMux I__6297 (
            .O(N__31686),
            .I(n1396));
    LocalMux I__6296 (
            .O(N__31675),
            .I(n1396));
    LocalMux I__6295 (
            .O(N__31664),
            .I(n1396));
    LocalMux I__6294 (
            .O(N__31655),
            .I(n1396));
    LocalMux I__6293 (
            .O(N__31642),
            .I(n1396));
    LocalMux I__6292 (
            .O(N__31631),
            .I(n1396));
    LocalMux I__6291 (
            .O(N__31618),
            .I(n1396));
    Odrv4 I__6290 (
            .O(N__31615),
            .I(n1396));
    Odrv4 I__6289 (
            .O(N__31604),
            .I(n1396));
    Odrv4 I__6288 (
            .O(N__31597),
            .I(n1396));
    Odrv4 I__6287 (
            .O(N__31592),
            .I(n1396));
    Odrv4 I__6286 (
            .O(N__31583),
            .I(n1396));
    LocalMux I__6285 (
            .O(N__31570),
            .I(n1396));
    InMux I__6284 (
            .O(N__31541),
            .I(N__31538));
    LocalMux I__6283 (
            .O(N__31538),
            .I(N__31534));
    InMux I__6282 (
            .O(N__31537),
            .I(N__31531));
    Span4Mux_h I__6281 (
            .O(N__31534),
            .I(N__31528));
    LocalMux I__6280 (
            .O(N__31531),
            .I(N__31525));
    Odrv4 I__6279 (
            .O(N__31528),
            .I(n2571));
    Odrv4 I__6278 (
            .O(N__31525),
            .I(n2571));
    CascadeMux I__6277 (
            .O(N__31520),
            .I(N__31517));
    InMux I__6276 (
            .O(N__31517),
            .I(N__31513));
    InMux I__6275 (
            .O(N__31516),
            .I(N__31509));
    LocalMux I__6274 (
            .O(N__31513),
            .I(N__31506));
    InMux I__6273 (
            .O(N__31512),
            .I(N__31502));
    LocalMux I__6272 (
            .O(N__31509),
            .I(N__31499));
    Span4Mux_h I__6271 (
            .O(N__31506),
            .I(N__31496));
    CascadeMux I__6270 (
            .O(N__31505),
            .I(N__31493));
    LocalMux I__6269 (
            .O(N__31502),
            .I(N__31486));
    Span4Mux_v I__6268 (
            .O(N__31499),
            .I(N__31486));
    Span4Mux_v I__6267 (
            .O(N__31496),
            .I(N__31486));
    InMux I__6266 (
            .O(N__31493),
            .I(N__31483));
    Span4Mux_v I__6265 (
            .O(N__31486),
            .I(N__31478));
    LocalMux I__6264 (
            .O(N__31483),
            .I(N__31478));
    Span4Mux_v I__6263 (
            .O(N__31478),
            .I(N__31475));
    Odrv4 I__6262 (
            .O(N__31475),
            .I(\c0.data_in_frame_9_4 ));
    InMux I__6261 (
            .O(N__31472),
            .I(N__31469));
    LocalMux I__6260 (
            .O(N__31469),
            .I(N__31466));
    Span4Mux_v I__6259 (
            .O(N__31466),
            .I(N__31463));
    Span4Mux_v I__6258 (
            .O(N__31463),
            .I(N__31459));
    InMux I__6257 (
            .O(N__31462),
            .I(N__31456));
    Odrv4 I__6256 (
            .O(N__31459),
            .I(data_in_17_7));
    LocalMux I__6255 (
            .O(N__31456),
            .I(data_in_17_7));
    InMux I__6254 (
            .O(N__31451),
            .I(N__31447));
    InMux I__6253 (
            .O(N__31450),
            .I(N__31444));
    LocalMux I__6252 (
            .O(N__31447),
            .I(N__31439));
    LocalMux I__6251 (
            .O(N__31444),
            .I(N__31439));
    Span4Mux_v I__6250 (
            .O(N__31439),
            .I(N__31436));
    Odrv4 I__6249 (
            .O(N__31436),
            .I(n2564));
    InMux I__6248 (
            .O(N__31433),
            .I(N__31430));
    LocalMux I__6247 (
            .O(N__31430),
            .I(N__31426));
    InMux I__6246 (
            .O(N__31429),
            .I(N__31423));
    Odrv4 I__6245 (
            .O(N__31426),
            .I(data_in_14_1));
    LocalMux I__6244 (
            .O(N__31423),
            .I(data_in_14_1));
    InMux I__6243 (
            .O(N__31418),
            .I(N__31415));
    LocalMux I__6242 (
            .O(N__31415),
            .I(N__31411));
    InMux I__6241 (
            .O(N__31414),
            .I(N__31406));
    Span4Mux_v I__6240 (
            .O(N__31411),
            .I(N__31403));
    CascadeMux I__6239 (
            .O(N__31410),
            .I(N__31400));
    InMux I__6238 (
            .O(N__31409),
            .I(N__31397));
    LocalMux I__6237 (
            .O(N__31406),
            .I(N__31392));
    Span4Mux_h I__6236 (
            .O(N__31403),
            .I(N__31392));
    InMux I__6235 (
            .O(N__31400),
            .I(N__31389));
    LocalMux I__6234 (
            .O(N__31397),
            .I(data_in_2_1));
    Odrv4 I__6233 (
            .O(N__31392),
            .I(data_in_2_1));
    LocalMux I__6232 (
            .O(N__31389),
            .I(data_in_2_1));
    InMux I__6231 (
            .O(N__31382),
            .I(N__31379));
    LocalMux I__6230 (
            .O(N__31379),
            .I(N__31373));
    InMux I__6229 (
            .O(N__31378),
            .I(N__31370));
    InMux I__6228 (
            .O(N__31377),
            .I(N__31367));
    InMux I__6227 (
            .O(N__31376),
            .I(N__31364));
    Span4Mux_v I__6226 (
            .O(N__31373),
            .I(N__31358));
    LocalMux I__6225 (
            .O(N__31370),
            .I(N__31358));
    LocalMux I__6224 (
            .O(N__31367),
            .I(N__31355));
    LocalMux I__6223 (
            .O(N__31364),
            .I(N__31352));
    InMux I__6222 (
            .O(N__31363),
            .I(N__31349));
    Span4Mux_h I__6221 (
            .O(N__31358),
            .I(N__31346));
    Span4Mux_h I__6220 (
            .O(N__31355),
            .I(N__31341));
    Span4Mux_h I__6219 (
            .O(N__31352),
            .I(N__31341));
    LocalMux I__6218 (
            .O(N__31349),
            .I(data_in_1_1));
    Odrv4 I__6217 (
            .O(N__31346),
            .I(data_in_1_1));
    Odrv4 I__6216 (
            .O(N__31341),
            .I(data_in_1_1));
    InMux I__6215 (
            .O(N__31334),
            .I(N__31328));
    InMux I__6214 (
            .O(N__31333),
            .I(N__31328));
    LocalMux I__6213 (
            .O(N__31328),
            .I(data_in_13_1));
    InMux I__6212 (
            .O(N__31325),
            .I(N__31319));
    InMux I__6211 (
            .O(N__31324),
            .I(N__31319));
    LocalMux I__6210 (
            .O(N__31319),
            .I(data_in_12_1));
    InMux I__6209 (
            .O(N__31316),
            .I(N__31313));
    LocalMux I__6208 (
            .O(N__31313),
            .I(N__31310));
    Span4Mux_h I__6207 (
            .O(N__31310),
            .I(N__31306));
    InMux I__6206 (
            .O(N__31309),
            .I(N__31303));
    Odrv4 I__6205 (
            .O(N__31306),
            .I(data_in_11_1));
    LocalMux I__6204 (
            .O(N__31303),
            .I(data_in_11_1));
    InMux I__6203 (
            .O(N__31298),
            .I(N__31295));
    LocalMux I__6202 (
            .O(N__31295),
            .I(N__31292));
    Span4Mux_h I__6201 (
            .O(N__31292),
            .I(N__31288));
    CascadeMux I__6200 (
            .O(N__31291),
            .I(N__31284));
    Span4Mux_h I__6199 (
            .O(N__31288),
            .I(N__31281));
    InMux I__6198 (
            .O(N__31287),
            .I(N__31276));
    InMux I__6197 (
            .O(N__31284),
            .I(N__31276));
    Odrv4 I__6196 (
            .O(N__31281),
            .I(data_in_6_6));
    LocalMux I__6195 (
            .O(N__31276),
            .I(data_in_6_6));
    InMux I__6194 (
            .O(N__31271),
            .I(N__31267));
    InMux I__6193 (
            .O(N__31270),
            .I(N__31264));
    LocalMux I__6192 (
            .O(N__31267),
            .I(N__31260));
    LocalMux I__6191 (
            .O(N__31264),
            .I(N__31257));
    InMux I__6190 (
            .O(N__31263),
            .I(N__31254));
    Span4Mux_v I__6189 (
            .O(N__31260),
            .I(N__31251));
    Sp12to4 I__6188 (
            .O(N__31257),
            .I(N__31248));
    LocalMux I__6187 (
            .O(N__31254),
            .I(N__31244));
    Sp12to4 I__6186 (
            .O(N__31251),
            .I(N__31239));
    Span12Mux_s11_v I__6185 (
            .O(N__31248),
            .I(N__31239));
    InMux I__6184 (
            .O(N__31247),
            .I(N__31236));
    Span4Mux_h I__6183 (
            .O(N__31244),
            .I(N__31233));
    Odrv12 I__6182 (
            .O(N__31239),
            .I(data_in_5_6));
    LocalMux I__6181 (
            .O(N__31236),
            .I(data_in_5_6));
    Odrv4 I__6180 (
            .O(N__31233),
            .I(data_in_5_6));
    InMux I__6179 (
            .O(N__31226),
            .I(N__31223));
    LocalMux I__6178 (
            .O(N__31223),
            .I(N__31220));
    Span4Mux_h I__6177 (
            .O(N__31220),
            .I(N__31216));
    InMux I__6176 (
            .O(N__31219),
            .I(N__31213));
    Sp12to4 I__6175 (
            .O(N__31216),
            .I(N__31210));
    LocalMux I__6174 (
            .O(N__31213),
            .I(data_out_frame2_9_4));
    Odrv12 I__6173 (
            .O(N__31210),
            .I(data_out_frame2_9_4));
    InMux I__6172 (
            .O(N__31205),
            .I(N__31201));
    InMux I__6171 (
            .O(N__31204),
            .I(N__31198));
    LocalMux I__6170 (
            .O(N__31201),
            .I(N__31195));
    LocalMux I__6169 (
            .O(N__31198),
            .I(data_out_frame2_8_4));
    Odrv12 I__6168 (
            .O(N__31195),
            .I(data_out_frame2_8_4));
    CascadeMux I__6167 (
            .O(N__31190),
            .I(N__31187));
    InMux I__6166 (
            .O(N__31187),
            .I(N__31184));
    LocalMux I__6165 (
            .O(N__31184),
            .I(\c0.n8 ));
    InMux I__6164 (
            .O(N__31181),
            .I(N__31178));
    LocalMux I__6163 (
            .O(N__31178),
            .I(N__31175));
    Span4Mux_v I__6162 (
            .O(N__31175),
            .I(N__31172));
    Span4Mux_v I__6161 (
            .O(N__31172),
            .I(N__31168));
    InMux I__6160 (
            .O(N__31171),
            .I(N__31165));
    Span4Mux_v I__6159 (
            .O(N__31168),
            .I(N__31162));
    LocalMux I__6158 (
            .O(N__31165),
            .I(\c0.data_out_frame2_0_1 ));
    Odrv4 I__6157 (
            .O(N__31162),
            .I(\c0.data_out_frame2_0_1 ));
    InMux I__6156 (
            .O(N__31157),
            .I(N__31147));
    InMux I__6155 (
            .O(N__31156),
            .I(N__31147));
    InMux I__6154 (
            .O(N__31155),
            .I(N__31147));
    InMux I__6153 (
            .O(N__31154),
            .I(N__31144));
    LocalMux I__6152 (
            .O(N__31147),
            .I(N__31135));
    LocalMux I__6151 (
            .O(N__31144),
            .I(N__31135));
    CascadeMux I__6150 (
            .O(N__31143),
            .I(N__31125));
    CascadeMux I__6149 (
            .O(N__31142),
            .I(N__31119));
    InMux I__6148 (
            .O(N__31141),
            .I(N__31113));
    InMux I__6147 (
            .O(N__31140),
            .I(N__31113));
    Span4Mux_h I__6146 (
            .O(N__31135),
            .I(N__31110));
    InMux I__6145 (
            .O(N__31134),
            .I(N__31101));
    InMux I__6144 (
            .O(N__31133),
            .I(N__31101));
    InMux I__6143 (
            .O(N__31132),
            .I(N__31101));
    InMux I__6142 (
            .O(N__31131),
            .I(N__31101));
    CascadeMux I__6141 (
            .O(N__31130),
            .I(N__31097));
    InMux I__6140 (
            .O(N__31129),
            .I(N__31091));
    InMux I__6139 (
            .O(N__31128),
            .I(N__31088));
    InMux I__6138 (
            .O(N__31125),
            .I(N__31085));
    InMux I__6137 (
            .O(N__31124),
            .I(N__31081));
    InMux I__6136 (
            .O(N__31123),
            .I(N__31078));
    InMux I__6135 (
            .O(N__31122),
            .I(N__31066));
    InMux I__6134 (
            .O(N__31119),
            .I(N__31066));
    InMux I__6133 (
            .O(N__31118),
            .I(N__31066));
    LocalMux I__6132 (
            .O(N__31113),
            .I(N__31059));
    Span4Mux_h I__6131 (
            .O(N__31110),
            .I(N__31059));
    LocalMux I__6130 (
            .O(N__31101),
            .I(N__31059));
    InMux I__6129 (
            .O(N__31100),
            .I(N__31054));
    InMux I__6128 (
            .O(N__31097),
            .I(N__31054));
    CascadeMux I__6127 (
            .O(N__31096),
            .I(N__31049));
    InMux I__6126 (
            .O(N__31095),
            .I(N__31044));
    InMux I__6125 (
            .O(N__31094),
            .I(N__31044));
    LocalMux I__6124 (
            .O(N__31091),
            .I(N__31036));
    LocalMux I__6123 (
            .O(N__31088),
            .I(N__31036));
    LocalMux I__6122 (
            .O(N__31085),
            .I(N__31036));
    CascadeMux I__6121 (
            .O(N__31084),
            .I(N__31027));
    LocalMux I__6120 (
            .O(N__31081),
            .I(N__31024));
    LocalMux I__6119 (
            .O(N__31078),
            .I(N__31021));
    InMux I__6118 (
            .O(N__31077),
            .I(N__31016));
    InMux I__6117 (
            .O(N__31076),
            .I(N__31016));
    InMux I__6116 (
            .O(N__31075),
            .I(N__31009));
    InMux I__6115 (
            .O(N__31074),
            .I(N__31009));
    InMux I__6114 (
            .O(N__31073),
            .I(N__31009));
    LocalMux I__6113 (
            .O(N__31066),
            .I(N__31002));
    Span4Mux_v I__6112 (
            .O(N__31059),
            .I(N__31002));
    LocalMux I__6111 (
            .O(N__31054),
            .I(N__31002));
    InMux I__6110 (
            .O(N__31053),
            .I(N__30995));
    InMux I__6109 (
            .O(N__31052),
            .I(N__30995));
    InMux I__6108 (
            .O(N__31049),
            .I(N__30995));
    LocalMux I__6107 (
            .O(N__31044),
            .I(N__30992));
    InMux I__6106 (
            .O(N__31043),
            .I(N__30975));
    Span4Mux_v I__6105 (
            .O(N__31036),
            .I(N__30972));
    InMux I__6104 (
            .O(N__31035),
            .I(N__30969));
    InMux I__6103 (
            .O(N__31034),
            .I(N__30957));
    InMux I__6102 (
            .O(N__31033),
            .I(N__30957));
    InMux I__6101 (
            .O(N__31032),
            .I(N__30954));
    InMux I__6100 (
            .O(N__31031),
            .I(N__30951));
    InMux I__6099 (
            .O(N__31030),
            .I(N__30948));
    InMux I__6098 (
            .O(N__31027),
            .I(N__30945));
    Span4Mux_v I__6097 (
            .O(N__31024),
            .I(N__30942));
    Span4Mux_v I__6096 (
            .O(N__31021),
            .I(N__30931));
    LocalMux I__6095 (
            .O(N__31016),
            .I(N__30931));
    LocalMux I__6094 (
            .O(N__31009),
            .I(N__30931));
    Span4Mux_h I__6093 (
            .O(N__31002),
            .I(N__30931));
    LocalMux I__6092 (
            .O(N__30995),
            .I(N__30931));
    Span4Mux_v I__6091 (
            .O(N__30992),
            .I(N__30927));
    InMux I__6090 (
            .O(N__30991),
            .I(N__30924));
    InMux I__6089 (
            .O(N__30990),
            .I(N__30921));
    InMux I__6088 (
            .O(N__30989),
            .I(N__30916));
    InMux I__6087 (
            .O(N__30988),
            .I(N__30916));
    InMux I__6086 (
            .O(N__30987),
            .I(N__30911));
    InMux I__6085 (
            .O(N__30986),
            .I(N__30911));
    InMux I__6084 (
            .O(N__30985),
            .I(N__30908));
    InMux I__6083 (
            .O(N__30984),
            .I(N__30899));
    InMux I__6082 (
            .O(N__30983),
            .I(N__30899));
    InMux I__6081 (
            .O(N__30982),
            .I(N__30899));
    InMux I__6080 (
            .O(N__30981),
            .I(N__30899));
    InMux I__6079 (
            .O(N__30980),
            .I(N__30892));
    InMux I__6078 (
            .O(N__30979),
            .I(N__30892));
    InMux I__6077 (
            .O(N__30978),
            .I(N__30892));
    LocalMux I__6076 (
            .O(N__30975),
            .I(N__30885));
    Sp12to4 I__6075 (
            .O(N__30972),
            .I(N__30885));
    LocalMux I__6074 (
            .O(N__30969),
            .I(N__30885));
    InMux I__6073 (
            .O(N__30968),
            .I(N__30876));
    InMux I__6072 (
            .O(N__30967),
            .I(N__30876));
    InMux I__6071 (
            .O(N__30966),
            .I(N__30876));
    InMux I__6070 (
            .O(N__30965),
            .I(N__30876));
    CascadeMux I__6069 (
            .O(N__30964),
            .I(N__30871));
    InMux I__6068 (
            .O(N__30963),
            .I(N__30866));
    InMux I__6067 (
            .O(N__30962),
            .I(N__30866));
    LocalMux I__6066 (
            .O(N__30957),
            .I(N__30861));
    LocalMux I__6065 (
            .O(N__30954),
            .I(N__30861));
    LocalMux I__6064 (
            .O(N__30951),
            .I(N__30854));
    LocalMux I__6063 (
            .O(N__30948),
            .I(N__30854));
    LocalMux I__6062 (
            .O(N__30945),
            .I(N__30854));
    Span4Mux_v I__6061 (
            .O(N__30942),
            .I(N__30849));
    Span4Mux_v I__6060 (
            .O(N__30931),
            .I(N__30849));
    InMux I__6059 (
            .O(N__30930),
            .I(N__30846));
    Span4Mux_v I__6058 (
            .O(N__30927),
            .I(N__30841));
    LocalMux I__6057 (
            .O(N__30924),
            .I(N__30841));
    LocalMux I__6056 (
            .O(N__30921),
            .I(N__30824));
    LocalMux I__6055 (
            .O(N__30916),
            .I(N__30824));
    LocalMux I__6054 (
            .O(N__30911),
            .I(N__30824));
    LocalMux I__6053 (
            .O(N__30908),
            .I(N__30824));
    LocalMux I__6052 (
            .O(N__30899),
            .I(N__30824));
    LocalMux I__6051 (
            .O(N__30892),
            .I(N__30824));
    Span12Mux_h I__6050 (
            .O(N__30885),
            .I(N__30824));
    LocalMux I__6049 (
            .O(N__30876),
            .I(N__30824));
    InMux I__6048 (
            .O(N__30875),
            .I(N__30817));
    InMux I__6047 (
            .O(N__30874),
            .I(N__30817));
    InMux I__6046 (
            .O(N__30871),
            .I(N__30817));
    LocalMux I__6045 (
            .O(N__30866),
            .I(N__30808));
    Span4Mux_v I__6044 (
            .O(N__30861),
            .I(N__30808));
    Span4Mux_v I__6043 (
            .O(N__30854),
            .I(N__30808));
    Span4Mux_h I__6042 (
            .O(N__30849),
            .I(N__30808));
    LocalMux I__6041 (
            .O(N__30846),
            .I(\c0.byte_transmit_counter2_1 ));
    Odrv4 I__6040 (
            .O(N__30841),
            .I(\c0.byte_transmit_counter2_1 ));
    Odrv12 I__6039 (
            .O(N__30824),
            .I(\c0.byte_transmit_counter2_1 ));
    LocalMux I__6038 (
            .O(N__30817),
            .I(\c0.byte_transmit_counter2_1 ));
    Odrv4 I__6037 (
            .O(N__30808),
            .I(\c0.byte_transmit_counter2_1 ));
    InMux I__6036 (
            .O(N__30797),
            .I(N__30782));
    InMux I__6035 (
            .O(N__30796),
            .I(N__30782));
    InMux I__6034 (
            .O(N__30795),
            .I(N__30782));
    InMux I__6033 (
            .O(N__30794),
            .I(N__30777));
    InMux I__6032 (
            .O(N__30793),
            .I(N__30777));
    InMux I__6031 (
            .O(N__30792),
            .I(N__30774));
    InMux I__6030 (
            .O(N__30791),
            .I(N__30755));
    InMux I__6029 (
            .O(N__30790),
            .I(N__30750));
    InMux I__6028 (
            .O(N__30789),
            .I(N__30747));
    LocalMux I__6027 (
            .O(N__30782),
            .I(N__30740));
    LocalMux I__6026 (
            .O(N__30777),
            .I(N__30740));
    LocalMux I__6025 (
            .O(N__30774),
            .I(N__30740));
    InMux I__6024 (
            .O(N__30773),
            .I(N__30726));
    InMux I__6023 (
            .O(N__30772),
            .I(N__30726));
    InMux I__6022 (
            .O(N__30771),
            .I(N__30726));
    InMux I__6021 (
            .O(N__30770),
            .I(N__30723));
    InMux I__6020 (
            .O(N__30769),
            .I(N__30719));
    InMux I__6019 (
            .O(N__30768),
            .I(N__30714));
    InMux I__6018 (
            .O(N__30767),
            .I(N__30714));
    InMux I__6017 (
            .O(N__30766),
            .I(N__30699));
    InMux I__6016 (
            .O(N__30765),
            .I(N__30699));
    InMux I__6015 (
            .O(N__30764),
            .I(N__30699));
    InMux I__6014 (
            .O(N__30763),
            .I(N__30699));
    InMux I__6013 (
            .O(N__30762),
            .I(N__30699));
    InMux I__6012 (
            .O(N__30761),
            .I(N__30699));
    InMux I__6011 (
            .O(N__30760),
            .I(N__30699));
    InMux I__6010 (
            .O(N__30759),
            .I(N__30696));
    InMux I__6009 (
            .O(N__30758),
            .I(N__30691));
    LocalMux I__6008 (
            .O(N__30755),
            .I(N__30688));
    InMux I__6007 (
            .O(N__30754),
            .I(N__30685));
    InMux I__6006 (
            .O(N__30753),
            .I(N__30682));
    LocalMux I__6005 (
            .O(N__30750),
            .I(N__30675));
    LocalMux I__6004 (
            .O(N__30747),
            .I(N__30675));
    Span4Mux_s2_v I__6003 (
            .O(N__30740),
            .I(N__30675));
    InMux I__6002 (
            .O(N__30739),
            .I(N__30664));
    InMux I__6001 (
            .O(N__30738),
            .I(N__30664));
    InMux I__6000 (
            .O(N__30737),
            .I(N__30655));
    InMux I__5999 (
            .O(N__30736),
            .I(N__30655));
    InMux I__5998 (
            .O(N__30735),
            .I(N__30655));
    InMux I__5997 (
            .O(N__30734),
            .I(N__30655));
    InMux I__5996 (
            .O(N__30733),
            .I(N__30652));
    LocalMux I__5995 (
            .O(N__30726),
            .I(N__30649));
    LocalMux I__5994 (
            .O(N__30723),
            .I(N__30646));
    InMux I__5993 (
            .O(N__30722),
            .I(N__30640));
    LocalMux I__5992 (
            .O(N__30719),
            .I(N__30631));
    LocalMux I__5991 (
            .O(N__30714),
            .I(N__30631));
    LocalMux I__5990 (
            .O(N__30699),
            .I(N__30631));
    LocalMux I__5989 (
            .O(N__30696),
            .I(N__30631));
    InMux I__5988 (
            .O(N__30695),
            .I(N__30626));
    InMux I__5987 (
            .O(N__30694),
            .I(N__30626));
    LocalMux I__5986 (
            .O(N__30691),
            .I(N__30622));
    Span4Mux_h I__5985 (
            .O(N__30688),
            .I(N__30617));
    LocalMux I__5984 (
            .O(N__30685),
            .I(N__30617));
    LocalMux I__5983 (
            .O(N__30682),
            .I(N__30612));
    Span4Mux_v I__5982 (
            .O(N__30675),
            .I(N__30612));
    InMux I__5981 (
            .O(N__30674),
            .I(N__30609));
    InMux I__5980 (
            .O(N__30673),
            .I(N__30604));
    InMux I__5979 (
            .O(N__30672),
            .I(N__30604));
    InMux I__5978 (
            .O(N__30671),
            .I(N__30601));
    InMux I__5977 (
            .O(N__30670),
            .I(N__30598));
    InMux I__5976 (
            .O(N__30669),
            .I(N__30595));
    LocalMux I__5975 (
            .O(N__30664),
            .I(N__30590));
    LocalMux I__5974 (
            .O(N__30655),
            .I(N__30590));
    LocalMux I__5973 (
            .O(N__30652),
            .I(N__30585));
    Span4Mux_h I__5972 (
            .O(N__30649),
            .I(N__30585));
    Span4Mux_v I__5971 (
            .O(N__30646),
            .I(N__30582));
    InMux I__5970 (
            .O(N__30645),
            .I(N__30575));
    InMux I__5969 (
            .O(N__30644),
            .I(N__30575));
    InMux I__5968 (
            .O(N__30643),
            .I(N__30575));
    LocalMux I__5967 (
            .O(N__30640),
            .I(N__30568));
    Span4Mux_h I__5966 (
            .O(N__30631),
            .I(N__30568));
    LocalMux I__5965 (
            .O(N__30626),
            .I(N__30568));
    CascadeMux I__5964 (
            .O(N__30625),
            .I(N__30565));
    Span4Mux_v I__5963 (
            .O(N__30622),
            .I(N__30555));
    Span4Mux_v I__5962 (
            .O(N__30617),
            .I(N__30555));
    Span4Mux_v I__5961 (
            .O(N__30612),
            .I(N__30550));
    LocalMux I__5960 (
            .O(N__30609),
            .I(N__30550));
    LocalMux I__5959 (
            .O(N__30604),
            .I(N__30537));
    LocalMux I__5958 (
            .O(N__30601),
            .I(N__30537));
    LocalMux I__5957 (
            .O(N__30598),
            .I(N__30537));
    LocalMux I__5956 (
            .O(N__30595),
            .I(N__30537));
    Span4Mux_v I__5955 (
            .O(N__30590),
            .I(N__30537));
    Span4Mux_v I__5954 (
            .O(N__30585),
            .I(N__30537));
    Span4Mux_h I__5953 (
            .O(N__30582),
            .I(N__30532));
    LocalMux I__5952 (
            .O(N__30575),
            .I(N__30532));
    Span4Mux_v I__5951 (
            .O(N__30568),
            .I(N__30529));
    InMux I__5950 (
            .O(N__30565),
            .I(N__30526));
    InMux I__5949 (
            .O(N__30564),
            .I(N__30523));
    InMux I__5948 (
            .O(N__30563),
            .I(N__30514));
    InMux I__5947 (
            .O(N__30562),
            .I(N__30514));
    InMux I__5946 (
            .O(N__30561),
            .I(N__30514));
    InMux I__5945 (
            .O(N__30560),
            .I(N__30514));
    Span4Mux_v I__5944 (
            .O(N__30555),
            .I(N__30509));
    Span4Mux_h I__5943 (
            .O(N__30550),
            .I(N__30509));
    Span4Mux_v I__5942 (
            .O(N__30537),
            .I(N__30504));
    Span4Mux_v I__5941 (
            .O(N__30532),
            .I(N__30504));
    Span4Mux_h I__5940 (
            .O(N__30529),
            .I(N__30501));
    LocalMux I__5939 (
            .O(N__30526),
            .I(\c0.byte_transmit_counter2_0 ));
    LocalMux I__5938 (
            .O(N__30523),
            .I(\c0.byte_transmit_counter2_0 ));
    LocalMux I__5937 (
            .O(N__30514),
            .I(\c0.byte_transmit_counter2_0 ));
    Odrv4 I__5936 (
            .O(N__30509),
            .I(\c0.byte_transmit_counter2_0 ));
    Odrv4 I__5935 (
            .O(N__30504),
            .I(\c0.byte_transmit_counter2_0 ));
    Odrv4 I__5934 (
            .O(N__30501),
            .I(\c0.byte_transmit_counter2_0 ));
    InMux I__5933 (
            .O(N__30488),
            .I(N__30485));
    LocalMux I__5932 (
            .O(N__30485),
            .I(N__30482));
    Span4Mux_s3_h I__5931 (
            .O(N__30482),
            .I(N__30479));
    Span4Mux_h I__5930 (
            .O(N__30479),
            .I(N__30476));
    Odrv4 I__5929 (
            .O(N__30476),
            .I(\c0.n18086 ));
    InMux I__5928 (
            .O(N__30473),
            .I(N__30469));
    InMux I__5927 (
            .O(N__30472),
            .I(N__30466));
    LocalMux I__5926 (
            .O(N__30469),
            .I(N__30463));
    LocalMux I__5925 (
            .O(N__30466),
            .I(N__30457));
    Span4Mux_h I__5924 (
            .O(N__30463),
            .I(N__30457));
    InMux I__5923 (
            .O(N__30462),
            .I(N__30454));
    Span4Mux_v I__5922 (
            .O(N__30457),
            .I(N__30451));
    LocalMux I__5921 (
            .O(N__30454),
            .I(data_in_10_7));
    Odrv4 I__5920 (
            .O(N__30451),
            .I(data_in_10_7));
    InMux I__5919 (
            .O(N__30446),
            .I(N__30440));
    InMux I__5918 (
            .O(N__30445),
            .I(N__30440));
    LocalMux I__5917 (
            .O(N__30440),
            .I(data_in_11_7));
    InMux I__5916 (
            .O(N__30437),
            .I(N__30431));
    InMux I__5915 (
            .O(N__30436),
            .I(N__30431));
    LocalMux I__5914 (
            .O(N__30431),
            .I(data_in_12_7));
    InMux I__5913 (
            .O(N__30428),
            .I(N__30422));
    InMux I__5912 (
            .O(N__30427),
            .I(N__30422));
    LocalMux I__5911 (
            .O(N__30422),
            .I(data_in_13_7));
    InMux I__5910 (
            .O(N__30419),
            .I(N__30413));
    InMux I__5909 (
            .O(N__30418),
            .I(N__30413));
    LocalMux I__5908 (
            .O(N__30413),
            .I(data_in_14_7));
    InMux I__5907 (
            .O(N__30410),
            .I(N__30407));
    LocalMux I__5906 (
            .O(N__30407),
            .I(N__30403));
    InMux I__5905 (
            .O(N__30406),
            .I(N__30400));
    Odrv12 I__5904 (
            .O(N__30403),
            .I(data_in_16_7));
    LocalMux I__5903 (
            .O(N__30400),
            .I(data_in_16_7));
    InMux I__5902 (
            .O(N__30395),
            .I(N__30389));
    InMux I__5901 (
            .O(N__30394),
            .I(N__30389));
    LocalMux I__5900 (
            .O(N__30389),
            .I(data_in_15_7));
    CascadeMux I__5899 (
            .O(N__30386),
            .I(\c0.rx.n97_cascade_ ));
    InMux I__5898 (
            .O(N__30383),
            .I(N__30380));
    LocalMux I__5897 (
            .O(N__30380),
            .I(\c0.rx.n17345 ));
    InMux I__5896 (
            .O(N__30377),
            .I(N__30367));
    InMux I__5895 (
            .O(N__30376),
            .I(N__30367));
    InMux I__5894 (
            .O(N__30375),
            .I(N__30364));
    InMux I__5893 (
            .O(N__30374),
            .I(N__30359));
    InMux I__5892 (
            .O(N__30373),
            .I(N__30359));
    InMux I__5891 (
            .O(N__30372),
            .I(N__30356));
    LocalMux I__5890 (
            .O(N__30367),
            .I(n13880));
    LocalMux I__5889 (
            .O(N__30364),
            .I(n13880));
    LocalMux I__5888 (
            .O(N__30359),
            .I(n13880));
    LocalMux I__5887 (
            .O(N__30356),
            .I(n13880));
    InMux I__5886 (
            .O(N__30347),
            .I(N__30344));
    LocalMux I__5885 (
            .O(N__30344),
            .I(n222));
    CascadeMux I__5884 (
            .O(N__30341),
            .I(N__30338));
    InMux I__5883 (
            .O(N__30338),
            .I(N__30335));
    LocalMux I__5882 (
            .O(N__30335),
            .I(N__30330));
    InMux I__5881 (
            .O(N__30334),
            .I(N__30327));
    InMux I__5880 (
            .O(N__30333),
            .I(N__30324));
    Odrv4 I__5879 (
            .O(N__30330),
            .I(r_Clock_Count_4_adj_2620));
    LocalMux I__5878 (
            .O(N__30327),
            .I(r_Clock_Count_4_adj_2620));
    LocalMux I__5877 (
            .O(N__30324),
            .I(r_Clock_Count_4_adj_2620));
    CascadeMux I__5876 (
            .O(N__30317),
            .I(N__30311));
    InMux I__5875 (
            .O(N__30316),
            .I(N__30306));
    InMux I__5874 (
            .O(N__30315),
            .I(N__30295));
    InMux I__5873 (
            .O(N__30314),
            .I(N__30295));
    InMux I__5872 (
            .O(N__30311),
            .I(N__30295));
    InMux I__5871 (
            .O(N__30310),
            .I(N__30295));
    InMux I__5870 (
            .O(N__30309),
            .I(N__30295));
    LocalMux I__5869 (
            .O(N__30306),
            .I(N__30288));
    LocalMux I__5868 (
            .O(N__30295),
            .I(N__30288));
    InMux I__5867 (
            .O(N__30294),
            .I(N__30283));
    InMux I__5866 (
            .O(N__30293),
            .I(N__30283));
    Odrv4 I__5865 (
            .O(N__30288),
            .I(n3));
    LocalMux I__5864 (
            .O(N__30283),
            .I(n3));
    InMux I__5863 (
            .O(N__30278),
            .I(N__30275));
    LocalMux I__5862 (
            .O(N__30275),
            .I(\c0.rx.n18001 ));
    CascadeMux I__5861 (
            .O(N__30272),
            .I(n17856_cascade_));
    InMux I__5860 (
            .O(N__30269),
            .I(N__30266));
    LocalMux I__5859 (
            .O(N__30266),
            .I(n17855));
    IoInMux I__5858 (
            .O(N__30263),
            .I(N__30260));
    LocalMux I__5857 (
            .O(N__30260),
            .I(N__30257));
    IoSpan4Mux I__5856 (
            .O(N__30257),
            .I(N__30254));
    Odrv4 I__5855 (
            .O(N__30254),
            .I(LED_c));
    InMux I__5854 (
            .O(N__30251),
            .I(N__30247));
    InMux I__5853 (
            .O(N__30250),
            .I(N__30244));
    LocalMux I__5852 (
            .O(N__30247),
            .I(\c0.rx.n112 ));
    LocalMux I__5851 (
            .O(N__30244),
            .I(\c0.rx.n112 ));
    InMux I__5850 (
            .O(N__30239),
            .I(N__30236));
    LocalMux I__5849 (
            .O(N__30236),
            .I(N__30232));
    InMux I__5848 (
            .O(N__30235),
            .I(N__30229));
    Span4Mux_v I__5847 (
            .O(N__30232),
            .I(N__30226));
    LocalMux I__5846 (
            .O(N__30229),
            .I(data_out_frame2_7_4));
    Odrv4 I__5845 (
            .O(N__30226),
            .I(data_out_frame2_7_4));
    InMux I__5844 (
            .O(N__30221),
            .I(N__30218));
    LocalMux I__5843 (
            .O(N__30218),
            .I(N__30215));
    Span4Mux_s2_v I__5842 (
            .O(N__30215),
            .I(N__30211));
    InMux I__5841 (
            .O(N__30214),
            .I(N__30208));
    Span4Mux_h I__5840 (
            .O(N__30211),
            .I(N__30205));
    LocalMux I__5839 (
            .O(N__30208),
            .I(data_out_frame2_6_4));
    Odrv4 I__5838 (
            .O(N__30205),
            .I(data_out_frame2_6_4));
    InMux I__5837 (
            .O(N__30200),
            .I(N__30197));
    LocalMux I__5836 (
            .O(N__30197),
            .I(\c0.n5_adj_2425 ));
    InMux I__5835 (
            .O(N__30194),
            .I(N__30191));
    LocalMux I__5834 (
            .O(N__30191),
            .I(N__30188));
    Span4Mux_h I__5833 (
            .O(N__30188),
            .I(N__30185));
    Odrv4 I__5832 (
            .O(N__30185),
            .I(\c0.rx.n79 ));
    InMux I__5831 (
            .O(N__30182),
            .I(N__30179));
    LocalMux I__5830 (
            .O(N__30179),
            .I(N__30176));
    Odrv12 I__5829 (
            .O(N__30176),
            .I(\c0.rx.n18597 ));
    InMux I__5828 (
            .O(N__30173),
            .I(N__30170));
    LocalMux I__5827 (
            .O(N__30170),
            .I(N__30167));
    Span4Mux_h I__5826 (
            .O(N__30167),
            .I(N__30164));
    Span4Mux_h I__5825 (
            .O(N__30164),
            .I(N__30161));
    Odrv4 I__5824 (
            .O(N__30161),
            .I(\c0.rx.r_Rx_Data_R ));
    InMux I__5823 (
            .O(N__30158),
            .I(N__30152));
    InMux I__5822 (
            .O(N__30157),
            .I(N__30152));
    LocalMux I__5821 (
            .O(N__30152),
            .I(\c0.rx.n13537 ));
    InMux I__5820 (
            .O(N__30149),
            .I(N__30143));
    InMux I__5819 (
            .O(N__30148),
            .I(N__30143));
    LocalMux I__5818 (
            .O(N__30143),
            .I(\c0.rx.n4_adj_2424 ));
    InMux I__5817 (
            .O(N__30140),
            .I(N__30133));
    InMux I__5816 (
            .O(N__30139),
            .I(N__30133));
    InMux I__5815 (
            .O(N__30138),
            .I(N__30130));
    LocalMux I__5814 (
            .O(N__30133),
            .I(\c0.rx.n17381 ));
    LocalMux I__5813 (
            .O(N__30130),
            .I(\c0.rx.n17381 ));
    CascadeMux I__5812 (
            .O(N__30125),
            .I(\c0.rx.n18003_cascade_ ));
    CascadeMux I__5811 (
            .O(N__30122),
            .I(n13880_cascade_));
    InMux I__5810 (
            .O(N__30119),
            .I(N__30113));
    InMux I__5809 (
            .O(N__30118),
            .I(N__30113));
    LocalMux I__5808 (
            .O(N__30113),
            .I(\c0.rx.n10193 ));
    InMux I__5807 (
            .O(N__30110),
            .I(N__30104));
    InMux I__5806 (
            .O(N__30109),
            .I(N__30101));
    InMux I__5805 (
            .O(N__30108),
            .I(N__30096));
    InMux I__5804 (
            .O(N__30107),
            .I(N__30096));
    LocalMux I__5803 (
            .O(N__30104),
            .I(r_Clock_Count_2_adj_2622));
    LocalMux I__5802 (
            .O(N__30101),
            .I(r_Clock_Count_2_adj_2622));
    LocalMux I__5801 (
            .O(N__30096),
            .I(r_Clock_Count_2_adj_2622));
    CascadeMux I__5800 (
            .O(N__30089),
            .I(N__30086));
    InMux I__5799 (
            .O(N__30086),
            .I(N__30077));
    InMux I__5798 (
            .O(N__30085),
            .I(N__30077));
    InMux I__5797 (
            .O(N__30084),
            .I(N__30077));
    LocalMux I__5796 (
            .O(N__30077),
            .I(\c0.rx.n124 ));
    CascadeMux I__5795 (
            .O(N__30074),
            .I(N__30071));
    InMux I__5794 (
            .O(N__30071),
            .I(N__30065));
    InMux I__5793 (
            .O(N__30070),
            .I(N__30062));
    InMux I__5792 (
            .O(N__30069),
            .I(N__30059));
    InMux I__5791 (
            .O(N__30068),
            .I(N__30056));
    LocalMux I__5790 (
            .O(N__30065),
            .I(r_Clock_Count_3_adj_2621));
    LocalMux I__5789 (
            .O(N__30062),
            .I(r_Clock_Count_3_adj_2621));
    LocalMux I__5788 (
            .O(N__30059),
            .I(r_Clock_Count_3_adj_2621));
    LocalMux I__5787 (
            .O(N__30056),
            .I(r_Clock_Count_3_adj_2621));
    InMux I__5786 (
            .O(N__30047),
            .I(N__30044));
    LocalMux I__5785 (
            .O(N__30044),
            .I(N__30041));
    Span4Mux_s2_h I__5784 (
            .O(N__30041),
            .I(N__30037));
    InMux I__5783 (
            .O(N__30040),
            .I(N__30034));
    Span4Mux_h I__5782 (
            .O(N__30037),
            .I(N__30031));
    LocalMux I__5781 (
            .O(N__30034),
            .I(data_out_frame2_13_0));
    Odrv4 I__5780 (
            .O(N__30031),
            .I(data_out_frame2_13_0));
    InMux I__5779 (
            .O(N__30026),
            .I(N__30020));
    InMux I__5778 (
            .O(N__30025),
            .I(N__30020));
    LocalMux I__5777 (
            .O(N__30020),
            .I(data_in_18_5));
    CascadeMux I__5776 (
            .O(N__30017),
            .I(n8562_cascade_));
    InMux I__5775 (
            .O(N__30014),
            .I(N__30010));
    InMux I__5774 (
            .O(N__30013),
            .I(N__30007));
    LocalMux I__5773 (
            .O(N__30010),
            .I(rx_data_2));
    LocalMux I__5772 (
            .O(N__30007),
            .I(rx_data_2));
    CascadeMux I__5771 (
            .O(N__30002),
            .I(\c0.rx.n2_cascade_ ));
    InMux I__5770 (
            .O(N__29999),
            .I(N__29996));
    LocalMux I__5769 (
            .O(N__29996),
            .I(\c0.rx.n2 ));
    CascadeMux I__5768 (
            .O(N__29993),
            .I(N__29989));
    InMux I__5767 (
            .O(N__29992),
            .I(N__29985));
    InMux I__5766 (
            .O(N__29989),
            .I(N__29982));
    InMux I__5765 (
            .O(N__29988),
            .I(N__29979));
    LocalMux I__5764 (
            .O(N__29985),
            .I(N__29976));
    LocalMux I__5763 (
            .O(N__29982),
            .I(r_Clock_Count_0_adj_2624));
    LocalMux I__5762 (
            .O(N__29979),
            .I(r_Clock_Count_0_adj_2624));
    Odrv4 I__5761 (
            .O(N__29976),
            .I(r_Clock_Count_0_adj_2624));
    CascadeMux I__5760 (
            .O(N__29969),
            .I(N__29966));
    InMux I__5759 (
            .O(N__29966),
            .I(N__29962));
    CascadeMux I__5758 (
            .O(N__29965),
            .I(N__29959));
    LocalMux I__5757 (
            .O(N__29962),
            .I(N__29955));
    InMux I__5756 (
            .O(N__29959),
            .I(N__29952));
    InMux I__5755 (
            .O(N__29958),
            .I(N__29949));
    Odrv4 I__5754 (
            .O(N__29955),
            .I(r_Clock_Count_1_adj_2623));
    LocalMux I__5753 (
            .O(N__29952),
            .I(r_Clock_Count_1_adj_2623));
    LocalMux I__5752 (
            .O(N__29949),
            .I(r_Clock_Count_1_adj_2623));
    InMux I__5751 (
            .O(N__29942),
            .I(N__29939));
    LocalMux I__5750 (
            .O(N__29939),
            .I(N__29935));
    InMux I__5749 (
            .O(N__29938),
            .I(N__29932));
    Odrv4 I__5748 (
            .O(N__29935),
            .I(data_in_19_0));
    LocalMux I__5747 (
            .O(N__29932),
            .I(data_in_19_0));
    InMux I__5746 (
            .O(N__29927),
            .I(N__29923));
    InMux I__5745 (
            .O(N__29926),
            .I(N__29920));
    LocalMux I__5744 (
            .O(N__29923),
            .I(N__29916));
    LocalMux I__5743 (
            .O(N__29920),
            .I(N__29913));
    InMux I__5742 (
            .O(N__29919),
            .I(N__29910));
    Span4Mux_v I__5741 (
            .O(N__29916),
            .I(N__29907));
    Span4Mux_v I__5740 (
            .O(N__29913),
            .I(N__29904));
    LocalMux I__5739 (
            .O(N__29910),
            .I(data_in_10_0));
    Odrv4 I__5738 (
            .O(N__29907),
            .I(data_in_10_0));
    Odrv4 I__5737 (
            .O(N__29904),
            .I(data_in_10_0));
    CascadeMux I__5736 (
            .O(N__29897),
            .I(N__29893));
    InMux I__5735 (
            .O(N__29896),
            .I(N__29890));
    InMux I__5734 (
            .O(N__29893),
            .I(N__29887));
    LocalMux I__5733 (
            .O(N__29890),
            .I(rx_data_4));
    LocalMux I__5732 (
            .O(N__29887),
            .I(rx_data_4));
    InMux I__5731 (
            .O(N__29882),
            .I(N__29878));
    InMux I__5730 (
            .O(N__29881),
            .I(N__29875));
    LocalMux I__5729 (
            .O(N__29878),
            .I(data_in_15_2));
    LocalMux I__5728 (
            .O(N__29875),
            .I(data_in_15_2));
    InMux I__5727 (
            .O(N__29870),
            .I(N__29866));
    InMux I__5726 (
            .O(N__29869),
            .I(N__29863));
    LocalMux I__5725 (
            .O(N__29866),
            .I(data_in_14_2));
    LocalMux I__5724 (
            .O(N__29863),
            .I(data_in_14_2));
    InMux I__5723 (
            .O(N__29858),
            .I(N__29855));
    LocalMux I__5722 (
            .O(N__29855),
            .I(N__29852));
    Span4Mux_h I__5721 (
            .O(N__29852),
            .I(N__29848));
    InMux I__5720 (
            .O(N__29851),
            .I(N__29845));
    Span4Mux_v I__5719 (
            .O(N__29848),
            .I(N__29841));
    LocalMux I__5718 (
            .O(N__29845),
            .I(N__29838));
    InMux I__5717 (
            .O(N__29844),
            .I(N__29835));
    Odrv4 I__5716 (
            .O(N__29841),
            .I(data_in_4_2));
    Odrv4 I__5715 (
            .O(N__29838),
            .I(data_in_4_2));
    LocalMux I__5714 (
            .O(N__29835),
            .I(data_in_4_2));
    InMux I__5713 (
            .O(N__29828),
            .I(N__29823));
    InMux I__5712 (
            .O(N__29827),
            .I(N__29820));
    InMux I__5711 (
            .O(N__29826),
            .I(N__29817));
    LocalMux I__5710 (
            .O(N__29823),
            .I(N__29814));
    LocalMux I__5709 (
            .O(N__29820),
            .I(data_in_9_7));
    LocalMux I__5708 (
            .O(N__29817),
            .I(data_in_9_7));
    Odrv4 I__5707 (
            .O(N__29814),
            .I(data_in_9_7));
    CascadeMux I__5706 (
            .O(N__29807),
            .I(N__29804));
    InMux I__5705 (
            .O(N__29804),
            .I(N__29801));
    LocalMux I__5704 (
            .O(N__29801),
            .I(N__29797));
    InMux I__5703 (
            .O(N__29800),
            .I(N__29794));
    Span4Mux_v I__5702 (
            .O(N__29797),
            .I(N__29791));
    LocalMux I__5701 (
            .O(N__29794),
            .I(N__29788));
    Span4Mux_v I__5700 (
            .O(N__29791),
            .I(N__29785));
    Span4Mux_v I__5699 (
            .O(N__29788),
            .I(N__29781));
    Span4Mux_h I__5698 (
            .O(N__29785),
            .I(N__29778));
    InMux I__5697 (
            .O(N__29784),
            .I(N__29775));
    Span4Mux_h I__5696 (
            .O(N__29781),
            .I(N__29772));
    Span4Mux_h I__5695 (
            .O(N__29778),
            .I(N__29769));
    LocalMux I__5694 (
            .O(N__29775),
            .I(data_in_8_7));
    Odrv4 I__5693 (
            .O(N__29772),
            .I(data_in_8_7));
    Odrv4 I__5692 (
            .O(N__29769),
            .I(data_in_8_7));
    InMux I__5691 (
            .O(N__29762),
            .I(N__29759));
    LocalMux I__5690 (
            .O(N__29759),
            .I(\c0.n10_adj_2536 ));
    InMux I__5689 (
            .O(N__29756),
            .I(N__29753));
    LocalMux I__5688 (
            .O(N__29753),
            .I(N__29750));
    Odrv4 I__5687 (
            .O(N__29750),
            .I(n18101));
    CascadeMux I__5686 (
            .O(N__29747),
            .I(N__29744));
    InMux I__5685 (
            .O(N__29744),
            .I(N__29741));
    LocalMux I__5684 (
            .O(N__29741),
            .I(N__29738));
    Span4Mux_v I__5683 (
            .O(N__29738),
            .I(N__29735));
    Span4Mux_h I__5682 (
            .O(N__29735),
            .I(N__29730));
    InMux I__5681 (
            .O(N__29734),
            .I(N__29727));
    InMux I__5680 (
            .O(N__29733),
            .I(N__29724));
    Odrv4 I__5679 (
            .O(N__29730),
            .I(data_in_8_3));
    LocalMux I__5678 (
            .O(N__29727),
            .I(data_in_8_3));
    LocalMux I__5677 (
            .O(N__29724),
            .I(data_in_8_3));
    CascadeMux I__5676 (
            .O(N__29717),
            .I(n8517_cascade_));
    InMux I__5675 (
            .O(N__29714),
            .I(N__29705));
    InMux I__5674 (
            .O(N__29713),
            .I(N__29705));
    InMux I__5673 (
            .O(N__29712),
            .I(N__29705));
    LocalMux I__5672 (
            .O(N__29705),
            .I(N__29702));
    Span4Mux_h I__5671 (
            .O(N__29702),
            .I(N__29696));
    InMux I__5670 (
            .O(N__29701),
            .I(N__29689));
    InMux I__5669 (
            .O(N__29700),
            .I(N__29689));
    InMux I__5668 (
            .O(N__29699),
            .I(N__29689));
    Span4Mux_h I__5667 (
            .O(N__29696),
            .I(N__29684));
    LocalMux I__5666 (
            .O(N__29689),
            .I(N__29684));
    Odrv4 I__5665 (
            .O(N__29684),
            .I(n17366));
    InMux I__5664 (
            .O(N__29681),
            .I(N__29678));
    LocalMux I__5663 (
            .O(N__29678),
            .I(N__29673));
    InMux I__5662 (
            .O(N__29677),
            .I(N__29668));
    InMux I__5661 (
            .O(N__29676),
            .I(N__29668));
    Span4Mux_h I__5660 (
            .O(N__29673),
            .I(N__29665));
    LocalMux I__5659 (
            .O(N__29668),
            .I(data_in_9_3));
    Odrv4 I__5658 (
            .O(N__29665),
            .I(data_in_9_3));
    InMux I__5657 (
            .O(N__29660),
            .I(N__29655));
    InMux I__5656 (
            .O(N__29659),
            .I(N__29652));
    InMux I__5655 (
            .O(N__29658),
            .I(N__29649));
    LocalMux I__5654 (
            .O(N__29655),
            .I(r_Clock_Count_0));
    LocalMux I__5653 (
            .O(N__29652),
            .I(r_Clock_Count_0));
    LocalMux I__5652 (
            .O(N__29649),
            .I(r_Clock_Count_0));
    CascadeMux I__5651 (
            .O(N__29642),
            .I(N__29637));
    InMux I__5650 (
            .O(N__29641),
            .I(N__29634));
    InMux I__5649 (
            .O(N__29640),
            .I(N__29631));
    InMux I__5648 (
            .O(N__29637),
            .I(N__29628));
    LocalMux I__5647 (
            .O(N__29634),
            .I(r_Clock_Count_5));
    LocalMux I__5646 (
            .O(N__29631),
            .I(r_Clock_Count_5));
    LocalMux I__5645 (
            .O(N__29628),
            .I(r_Clock_Count_5));
    InMux I__5644 (
            .O(N__29621),
            .I(N__29616));
    InMux I__5643 (
            .O(N__29620),
            .I(N__29613));
    InMux I__5642 (
            .O(N__29619),
            .I(N__29610));
    LocalMux I__5641 (
            .O(N__29616),
            .I(r_Clock_Count_3));
    LocalMux I__5640 (
            .O(N__29613),
            .I(r_Clock_Count_3));
    LocalMux I__5639 (
            .O(N__29610),
            .I(r_Clock_Count_3));
    InMux I__5638 (
            .O(N__29603),
            .I(N__29598));
    InMux I__5637 (
            .O(N__29602),
            .I(N__29595));
    InMux I__5636 (
            .O(N__29601),
            .I(N__29592));
    LocalMux I__5635 (
            .O(N__29598),
            .I(r_Clock_Count_4));
    LocalMux I__5634 (
            .O(N__29595),
            .I(r_Clock_Count_4));
    LocalMux I__5633 (
            .O(N__29592),
            .I(r_Clock_Count_4));
    CascadeMux I__5632 (
            .O(N__29585),
            .I(\c0.tx.n10_cascade_ ));
    InMux I__5631 (
            .O(N__29582),
            .I(N__29579));
    LocalMux I__5630 (
            .O(N__29579),
            .I(N__29574));
    InMux I__5629 (
            .O(N__29578),
            .I(N__29569));
    InMux I__5628 (
            .O(N__29577),
            .I(N__29569));
    Odrv12 I__5627 (
            .O(N__29574),
            .I(r_Clock_Count_1));
    LocalMux I__5626 (
            .O(N__29569),
            .I(r_Clock_Count_1));
    InMux I__5625 (
            .O(N__29564),
            .I(N__29558));
    InMux I__5624 (
            .O(N__29563),
            .I(N__29558));
    LocalMux I__5623 (
            .O(N__29558),
            .I(N__29554));
    InMux I__5622 (
            .O(N__29557),
            .I(N__29550));
    Span4Mux_v I__5621 (
            .O(N__29554),
            .I(N__29547));
    InMux I__5620 (
            .O(N__29553),
            .I(N__29544));
    LocalMux I__5619 (
            .O(N__29550),
            .I(N__29541));
    Span4Mux_h I__5618 (
            .O(N__29547),
            .I(N__29538));
    LocalMux I__5617 (
            .O(N__29544),
            .I(data_in_5_5));
    Odrv12 I__5616 (
            .O(N__29541),
            .I(data_in_5_5));
    Odrv4 I__5615 (
            .O(N__29538),
            .I(data_in_5_5));
    InMux I__5614 (
            .O(N__29531),
            .I(N__29527));
    InMux I__5613 (
            .O(N__29530),
            .I(N__29524));
    LocalMux I__5612 (
            .O(N__29527),
            .I(N__29518));
    LocalMux I__5611 (
            .O(N__29524),
            .I(N__29518));
    InMux I__5610 (
            .O(N__29523),
            .I(N__29515));
    Span4Mux_v I__5609 (
            .O(N__29518),
            .I(N__29512));
    LocalMux I__5608 (
            .O(N__29515),
            .I(data_in_10_1));
    Odrv4 I__5607 (
            .O(N__29512),
            .I(data_in_10_1));
    InMux I__5606 (
            .O(N__29507),
            .I(N__29503));
    InMux I__5605 (
            .O(N__29506),
            .I(N__29500));
    LocalMux I__5604 (
            .O(N__29503),
            .I(N__29497));
    LocalMux I__5603 (
            .O(N__29500),
            .I(N__29494));
    Span4Mux_v I__5602 (
            .O(N__29497),
            .I(N__29491));
    Span12Mux_v I__5601 (
            .O(N__29494),
            .I(N__29488));
    Span4Mux_h I__5600 (
            .O(N__29491),
            .I(N__29485));
    Odrv12 I__5599 (
            .O(N__29488),
            .I(\c0.n17544 ));
    Odrv4 I__5598 (
            .O(N__29485),
            .I(\c0.n17544 ));
    InMux I__5597 (
            .O(N__29480),
            .I(N__29476));
    InMux I__5596 (
            .O(N__29479),
            .I(N__29473));
    LocalMux I__5595 (
            .O(N__29476),
            .I(N__29470));
    LocalMux I__5594 (
            .O(N__29473),
            .I(N__29467));
    Span4Mux_h I__5593 (
            .O(N__29470),
            .I(N__29464));
    Span12Mux_h I__5592 (
            .O(N__29467),
            .I(N__29461));
    Span4Mux_v I__5591 (
            .O(N__29464),
            .I(N__29458));
    Odrv12 I__5590 (
            .O(N__29461),
            .I(\c0.n8056 ));
    Odrv4 I__5589 (
            .O(N__29458),
            .I(\c0.n8056 ));
    CascadeMux I__5588 (
            .O(N__29453),
            .I(n2566_cascade_));
    InMux I__5587 (
            .O(N__29450),
            .I(N__29447));
    LocalMux I__5586 (
            .O(N__29447),
            .I(N__29443));
    InMux I__5585 (
            .O(N__29446),
            .I(N__29440));
    Span4Mux_h I__5584 (
            .O(N__29443),
            .I(N__29437));
    LocalMux I__5583 (
            .O(N__29440),
            .I(N__29434));
    Odrv4 I__5582 (
            .O(N__29437),
            .I(n2561));
    Odrv4 I__5581 (
            .O(N__29434),
            .I(n2561));
    InMux I__5580 (
            .O(N__29429),
            .I(N__29426));
    LocalMux I__5579 (
            .O(N__29426),
            .I(\c0.n19 ));
    InMux I__5578 (
            .O(N__29423),
            .I(N__29420));
    LocalMux I__5577 (
            .O(N__29420),
            .I(N__29416));
    InMux I__5576 (
            .O(N__29419),
            .I(N__29413));
    Span4Mux_h I__5575 (
            .O(N__29416),
            .I(N__29409));
    LocalMux I__5574 (
            .O(N__29413),
            .I(N__29406));
    InMux I__5573 (
            .O(N__29412),
            .I(N__29403));
    Span4Mux_h I__5572 (
            .O(N__29409),
            .I(N__29400));
    Odrv4 I__5571 (
            .O(N__29406),
            .I(data_in_9_0));
    LocalMux I__5570 (
            .O(N__29403),
            .I(data_in_9_0));
    Odrv4 I__5569 (
            .O(N__29400),
            .I(data_in_9_0));
    InMux I__5568 (
            .O(N__29393),
            .I(N__29385));
    InMux I__5567 (
            .O(N__29392),
            .I(N__29382));
    InMux I__5566 (
            .O(N__29391),
            .I(N__29375));
    InMux I__5565 (
            .O(N__29390),
            .I(N__29375));
    InMux I__5564 (
            .O(N__29389),
            .I(N__29375));
    CascadeMux I__5563 (
            .O(N__29388),
            .I(N__29372));
    LocalMux I__5562 (
            .O(N__29385),
            .I(N__29365));
    LocalMux I__5561 (
            .O(N__29382),
            .I(N__29365));
    LocalMux I__5560 (
            .O(N__29375),
            .I(N__29365));
    InMux I__5559 (
            .O(N__29372),
            .I(N__29362));
    Span12Mux_s9_v I__5558 (
            .O(N__29365),
            .I(N__29357));
    LocalMux I__5557 (
            .O(N__29362),
            .I(N__29357));
    Span12Mux_h I__5556 (
            .O(N__29357),
            .I(N__29354));
    Odrv12 I__5555 (
            .O(N__29354),
            .I(\c0.data_in_frame_9_0 ));
    InMux I__5554 (
            .O(N__29351),
            .I(N__29348));
    LocalMux I__5553 (
            .O(N__29348),
            .I(N__29345));
    Span4Mux_h I__5552 (
            .O(N__29345),
            .I(N__29341));
    InMux I__5551 (
            .O(N__29344),
            .I(N__29338));
    Odrv4 I__5550 (
            .O(N__29341),
            .I(n2575));
    LocalMux I__5549 (
            .O(N__29338),
            .I(n2575));
    InMux I__5548 (
            .O(N__29333),
            .I(N__29330));
    LocalMux I__5547 (
            .O(N__29330),
            .I(N__29327));
    Span4Mux_h I__5546 (
            .O(N__29327),
            .I(N__29324));
    Span4Mux_v I__5545 (
            .O(N__29324),
            .I(N__29320));
    InMux I__5544 (
            .O(N__29323),
            .I(N__29317));
    Odrv4 I__5543 (
            .O(N__29320),
            .I(\c0.n17504 ));
    LocalMux I__5542 (
            .O(N__29317),
            .I(\c0.n17504 ));
    CascadeMux I__5541 (
            .O(N__29312),
            .I(\c0.n6_adj_2541_cascade_ ));
    InMux I__5540 (
            .O(N__29309),
            .I(N__29306));
    LocalMux I__5539 (
            .O(N__29306),
            .I(N__29303));
    Span4Mux_v I__5538 (
            .O(N__29303),
            .I(N__29300));
    Sp12to4 I__5537 (
            .O(N__29300),
            .I(N__29297));
    Odrv12 I__5536 (
            .O(N__29297),
            .I(\c0.n17591 ));
    InMux I__5535 (
            .O(N__29294),
            .I(N__29291));
    LocalMux I__5534 (
            .O(N__29291),
            .I(N__29288));
    Span4Mux_s2_v I__5533 (
            .O(N__29288),
            .I(N__29285));
    Span4Mux_v I__5532 (
            .O(N__29285),
            .I(N__29282));
    Odrv4 I__5531 (
            .O(N__29282),
            .I(\c0.data_out_frame2_20_4 ));
    InMux I__5530 (
            .O(N__29279),
            .I(N__29276));
    LocalMux I__5529 (
            .O(N__29276),
            .I(N__29273));
    Span4Mux_h I__5528 (
            .O(N__29273),
            .I(N__29270));
    Span4Mux_h I__5527 (
            .O(N__29270),
            .I(N__29266));
    InMux I__5526 (
            .O(N__29269),
            .I(N__29263));
    Odrv4 I__5525 (
            .O(N__29266),
            .I(\c0.n17488 ));
    LocalMux I__5524 (
            .O(N__29263),
            .I(\c0.n17488 ));
    InMux I__5523 (
            .O(N__29258),
            .I(N__29254));
    InMux I__5522 (
            .O(N__29257),
            .I(N__29251));
    LocalMux I__5521 (
            .O(N__29254),
            .I(N__29248));
    LocalMux I__5520 (
            .O(N__29251),
            .I(N__29240));
    Span4Mux_h I__5519 (
            .O(N__29248),
            .I(N__29240));
    InMux I__5518 (
            .O(N__29247),
            .I(N__29235));
    InMux I__5517 (
            .O(N__29246),
            .I(N__29235));
    CascadeMux I__5516 (
            .O(N__29245),
            .I(N__29232));
    Sp12to4 I__5515 (
            .O(N__29240),
            .I(N__29229));
    LocalMux I__5514 (
            .O(N__29235),
            .I(N__29226));
    InMux I__5513 (
            .O(N__29232),
            .I(N__29223));
    Span12Mux_s11_v I__5512 (
            .O(N__29229),
            .I(N__29220));
    Span4Mux_h I__5511 (
            .O(N__29226),
            .I(N__29215));
    LocalMux I__5510 (
            .O(N__29223),
            .I(N__29215));
    Odrv12 I__5509 (
            .O(N__29220),
            .I(data_in_frame_9_6));
    Odrv4 I__5508 (
            .O(N__29215),
            .I(data_in_frame_9_6));
    InMux I__5507 (
            .O(N__29210),
            .I(N__29207));
    LocalMux I__5506 (
            .O(N__29207),
            .I(N__29204));
    Odrv4 I__5505 (
            .O(N__29204),
            .I(n17479));
    CascadeMux I__5504 (
            .O(N__29201),
            .I(N__29198));
    InMux I__5503 (
            .O(N__29198),
            .I(N__29194));
    InMux I__5502 (
            .O(N__29197),
            .I(N__29191));
    LocalMux I__5501 (
            .O(N__29194),
            .I(N__29188));
    LocalMux I__5500 (
            .O(N__29191),
            .I(N__29185));
    Span4Mux_v I__5499 (
            .O(N__29188),
            .I(N__29180));
    Span4Mux_v I__5498 (
            .O(N__29185),
            .I(N__29180));
    Odrv4 I__5497 (
            .O(N__29180),
            .I(n9051));
    InMux I__5496 (
            .O(N__29177),
            .I(N__29174));
    LocalMux I__5495 (
            .O(N__29174),
            .I(N__29170));
    InMux I__5494 (
            .O(N__29173),
            .I(N__29167));
    Span4Mux_v I__5493 (
            .O(N__29170),
            .I(N__29162));
    LocalMux I__5492 (
            .O(N__29167),
            .I(N__29162));
    Span4Mux_v I__5491 (
            .O(N__29162),
            .I(N__29159));
    Odrv4 I__5490 (
            .O(N__29159),
            .I(n6_adj_2583));
    CascadeMux I__5489 (
            .O(N__29156),
            .I(N__29153));
    InMux I__5488 (
            .O(N__29153),
            .I(N__29150));
    LocalMux I__5487 (
            .O(N__29150),
            .I(N__29147));
    Span4Mux_s2_h I__5486 (
            .O(N__29147),
            .I(N__29144));
    Span4Mux_h I__5485 (
            .O(N__29144),
            .I(N__29141));
    Odrv4 I__5484 (
            .O(N__29141),
            .I(\c0.data_out_frame2_19_2 ));
    InMux I__5483 (
            .O(N__29138),
            .I(N__29135));
    LocalMux I__5482 (
            .O(N__29135),
            .I(N__29130));
    InMux I__5481 (
            .O(N__29134),
            .I(N__29127));
    CascadeMux I__5480 (
            .O(N__29133),
            .I(N__29123));
    Span4Mux_v I__5479 (
            .O(N__29130),
            .I(N__29119));
    LocalMux I__5478 (
            .O(N__29127),
            .I(N__29116));
    InMux I__5477 (
            .O(N__29126),
            .I(N__29113));
    InMux I__5476 (
            .O(N__29123),
            .I(N__29110));
    InMux I__5475 (
            .O(N__29122),
            .I(N__29107));
    Span4Mux_h I__5474 (
            .O(N__29119),
            .I(N__29102));
    Span4Mux_v I__5473 (
            .O(N__29116),
            .I(N__29102));
    LocalMux I__5472 (
            .O(N__29113),
            .I(\c0.data_in_frame_0_1 ));
    LocalMux I__5471 (
            .O(N__29110),
            .I(\c0.data_in_frame_0_1 ));
    LocalMux I__5470 (
            .O(N__29107),
            .I(\c0.data_in_frame_0_1 ));
    Odrv4 I__5469 (
            .O(N__29102),
            .I(\c0.data_in_frame_0_1 ));
    InMux I__5468 (
            .O(N__29093),
            .I(N__29090));
    LocalMux I__5467 (
            .O(N__29090),
            .I(N__29085));
    InMux I__5466 (
            .O(N__29089),
            .I(N__29081));
    InMux I__5465 (
            .O(N__29088),
            .I(N__29078));
    Span4Mux_h I__5464 (
            .O(N__29085),
            .I(N__29075));
    InMux I__5463 (
            .O(N__29084),
            .I(N__29072));
    LocalMux I__5462 (
            .O(N__29081),
            .I(N__29069));
    LocalMux I__5461 (
            .O(N__29078),
            .I(\c0.data_in_frame_3_6 ));
    Odrv4 I__5460 (
            .O(N__29075),
            .I(\c0.data_in_frame_3_6 ));
    LocalMux I__5459 (
            .O(N__29072),
            .I(\c0.data_in_frame_3_6 ));
    Odrv12 I__5458 (
            .O(N__29069),
            .I(\c0.data_in_frame_3_6 ));
    CascadeMux I__5457 (
            .O(N__29060),
            .I(N__29057));
    InMux I__5456 (
            .O(N__29057),
            .I(N__29053));
    InMux I__5455 (
            .O(N__29056),
            .I(N__29050));
    LocalMux I__5454 (
            .O(N__29053),
            .I(N__29047));
    LocalMux I__5453 (
            .O(N__29050),
            .I(N__29044));
    Span4Mux_h I__5452 (
            .O(N__29047),
            .I(N__29041));
    Span4Mux_h I__5451 (
            .O(N__29044),
            .I(N__29035));
    Span4Mux_h I__5450 (
            .O(N__29041),
            .I(N__29035));
    CascadeMux I__5449 (
            .O(N__29040),
            .I(N__29032));
    Span4Mux_v I__5448 (
            .O(N__29035),
            .I(N__29027));
    InMux I__5447 (
            .O(N__29032),
            .I(N__29022));
    InMux I__5446 (
            .O(N__29031),
            .I(N__29022));
    InMux I__5445 (
            .O(N__29030),
            .I(N__29019));
    Odrv4 I__5444 (
            .O(N__29027),
            .I(\c0.data_in_frame_2_1 ));
    LocalMux I__5443 (
            .O(N__29022),
            .I(\c0.data_in_frame_2_1 ));
    LocalMux I__5442 (
            .O(N__29019),
            .I(\c0.data_in_frame_2_1 ));
    InMux I__5441 (
            .O(N__29012),
            .I(N__29007));
    InMux I__5440 (
            .O(N__29011),
            .I(N__29002));
    InMux I__5439 (
            .O(N__29010),
            .I(N__29002));
    LocalMux I__5438 (
            .O(N__29007),
            .I(N__28998));
    LocalMux I__5437 (
            .O(N__29002),
            .I(N__28995));
    InMux I__5436 (
            .O(N__29001),
            .I(N__28992));
    Span12Mux_v I__5435 (
            .O(N__28998),
            .I(N__28989));
    Span4Mux_h I__5434 (
            .O(N__28995),
            .I(N__28986));
    LocalMux I__5433 (
            .O(N__28992),
            .I(\c0.data_in_frame_0_2 ));
    Odrv12 I__5432 (
            .O(N__28989),
            .I(\c0.data_in_frame_0_2 ));
    Odrv4 I__5431 (
            .O(N__28986),
            .I(\c0.data_in_frame_0_2 ));
    CascadeMux I__5430 (
            .O(N__28979),
            .I(N__28975));
    InMux I__5429 (
            .O(N__28978),
            .I(N__28971));
    InMux I__5428 (
            .O(N__28975),
            .I(N__28968));
    InMux I__5427 (
            .O(N__28974),
            .I(N__28965));
    LocalMux I__5426 (
            .O(N__28971),
            .I(N__28962));
    LocalMux I__5425 (
            .O(N__28968),
            .I(N__28959));
    LocalMux I__5424 (
            .O(N__28965),
            .I(N__28956));
    Span4Mux_h I__5423 (
            .O(N__28962),
            .I(N__28953));
    Span4Mux_h I__5422 (
            .O(N__28959),
            .I(N__28950));
    Span12Mux_s8_v I__5421 (
            .O(N__28956),
            .I(N__28947));
    Span4Mux_h I__5420 (
            .O(N__28953),
            .I(N__28942));
    Span4Mux_v I__5419 (
            .O(N__28950),
            .I(N__28942));
    Odrv12 I__5418 (
            .O(N__28947),
            .I(\c0.n9043 ));
    Odrv4 I__5417 (
            .O(N__28942),
            .I(\c0.n9043 ));
    InMux I__5416 (
            .O(N__28937),
            .I(N__28934));
    LocalMux I__5415 (
            .O(N__28934),
            .I(N__28930));
    InMux I__5414 (
            .O(N__28933),
            .I(N__28927));
    Span4Mux_h I__5413 (
            .O(N__28930),
            .I(N__28924));
    LocalMux I__5412 (
            .O(N__28927),
            .I(N__28921));
    Span4Mux_v I__5411 (
            .O(N__28924),
            .I(N__28917));
    Span4Mux_h I__5410 (
            .O(N__28921),
            .I(N__28914));
    InMux I__5409 (
            .O(N__28920),
            .I(N__28911));
    Span4Mux_v I__5408 (
            .O(N__28917),
            .I(N__28908));
    Span4Mux_h I__5407 (
            .O(N__28914),
            .I(N__28905));
    LocalMux I__5406 (
            .O(N__28911),
            .I(N__28902));
    Odrv4 I__5405 (
            .O(N__28908),
            .I(\c0.n8886 ));
    Odrv4 I__5404 (
            .O(N__28905),
            .I(\c0.n8886 ));
    Odrv12 I__5403 (
            .O(N__28902),
            .I(\c0.n8886 ));
    InMux I__5402 (
            .O(N__28895),
            .I(N__28891));
    InMux I__5401 (
            .O(N__28894),
            .I(N__28888));
    LocalMux I__5400 (
            .O(N__28891),
            .I(N__28885));
    LocalMux I__5399 (
            .O(N__28888),
            .I(\c0.n15927 ));
    Odrv4 I__5398 (
            .O(N__28885),
            .I(\c0.n15927 ));
    InMux I__5397 (
            .O(N__28880),
            .I(N__28877));
    LocalMux I__5396 (
            .O(N__28877),
            .I(N__28874));
    Span4Mux_v I__5395 (
            .O(N__28874),
            .I(N__28870));
    InMux I__5394 (
            .O(N__28873),
            .I(N__28867));
    Span4Mux_v I__5393 (
            .O(N__28870),
            .I(N__28864));
    LocalMux I__5392 (
            .O(N__28867),
            .I(N__28861));
    Span4Mux_v I__5391 (
            .O(N__28864),
            .I(N__28856));
    Span4Mux_v I__5390 (
            .O(N__28861),
            .I(N__28856));
    Sp12to4 I__5389 (
            .O(N__28856),
            .I(N__28853));
    Odrv12 I__5388 (
            .O(N__28853),
            .I(\c0.n17594 ));
    InMux I__5387 (
            .O(N__28850),
            .I(N__28846));
    InMux I__5386 (
            .O(N__28849),
            .I(N__28843));
    LocalMux I__5385 (
            .O(N__28846),
            .I(N__28840));
    LocalMux I__5384 (
            .O(N__28843),
            .I(N__28837));
    Span4Mux_v I__5383 (
            .O(N__28840),
            .I(N__28832));
    Span4Mux_h I__5382 (
            .O(N__28837),
            .I(N__28832));
    Odrv4 I__5381 (
            .O(N__28832),
            .I(\c0.n17412 ));
    CascadeMux I__5380 (
            .O(N__28829),
            .I(n2565_cascade_));
    InMux I__5379 (
            .O(N__28826),
            .I(N__28823));
    LocalMux I__5378 (
            .O(N__28823),
            .I(N__28820));
    Span4Mux_h I__5377 (
            .O(N__28820),
            .I(N__28816));
    InMux I__5376 (
            .O(N__28819),
            .I(N__28813));
    Odrv4 I__5375 (
            .O(N__28816),
            .I(n2574));
    LocalMux I__5374 (
            .O(N__28813),
            .I(n2574));
    InMux I__5373 (
            .O(N__28808),
            .I(N__28804));
    InMux I__5372 (
            .O(N__28807),
            .I(N__28801));
    LocalMux I__5371 (
            .O(N__28804),
            .I(N__28798));
    LocalMux I__5370 (
            .O(N__28801),
            .I(N__28795));
    Odrv4 I__5369 (
            .O(N__28798),
            .I(n17547));
    Odrv4 I__5368 (
            .O(N__28795),
            .I(n17547));
    CascadeMux I__5367 (
            .O(N__28790),
            .I(\c0.n23_cascade_ ));
    InMux I__5366 (
            .O(N__28787),
            .I(N__28784));
    LocalMux I__5365 (
            .O(N__28784),
            .I(\c0.n17536 ));
    InMux I__5364 (
            .O(N__28781),
            .I(N__28778));
    LocalMux I__5363 (
            .O(N__28778),
            .I(\c0.n28 ));
    InMux I__5362 (
            .O(N__28775),
            .I(N__28768));
    InMux I__5361 (
            .O(N__28774),
            .I(N__28768));
    InMux I__5360 (
            .O(N__28773),
            .I(N__28764));
    LocalMux I__5359 (
            .O(N__28768),
            .I(N__28761));
    InMux I__5358 (
            .O(N__28767),
            .I(N__28756));
    LocalMux I__5357 (
            .O(N__28764),
            .I(N__28753));
    Span12Mux_v I__5356 (
            .O(N__28761),
            .I(N__28750));
    InMux I__5355 (
            .O(N__28760),
            .I(N__28745));
    InMux I__5354 (
            .O(N__28759),
            .I(N__28745));
    LocalMux I__5353 (
            .O(N__28756),
            .I(N__28740));
    Span4Mux_v I__5352 (
            .O(N__28753),
            .I(N__28740));
    Odrv12 I__5351 (
            .O(N__28750),
            .I(data_in_frame_8_0));
    LocalMux I__5350 (
            .O(N__28745),
            .I(data_in_frame_8_0));
    Odrv4 I__5349 (
            .O(N__28740),
            .I(data_in_frame_8_0));
    InMux I__5348 (
            .O(N__28733),
            .I(N__28727));
    InMux I__5347 (
            .O(N__28732),
            .I(N__28727));
    LocalMux I__5346 (
            .O(N__28727),
            .I(N__28724));
    Span4Mux_v I__5345 (
            .O(N__28724),
            .I(N__28720));
    CascadeMux I__5344 (
            .O(N__28723),
            .I(N__28717));
    Span4Mux_h I__5343 (
            .O(N__28720),
            .I(N__28711));
    InMux I__5342 (
            .O(N__28717),
            .I(N__28706));
    InMux I__5341 (
            .O(N__28716),
            .I(N__28706));
    InMux I__5340 (
            .O(N__28715),
            .I(N__28701));
    InMux I__5339 (
            .O(N__28714),
            .I(N__28701));
    Odrv4 I__5338 (
            .O(N__28711),
            .I(data_in_frame_1_1));
    LocalMux I__5337 (
            .O(N__28706),
            .I(data_in_frame_1_1));
    LocalMux I__5336 (
            .O(N__28701),
            .I(data_in_frame_1_1));
    InMux I__5335 (
            .O(N__28694),
            .I(N__28689));
    InMux I__5334 (
            .O(N__28693),
            .I(N__28686));
    InMux I__5333 (
            .O(N__28692),
            .I(N__28683));
    LocalMux I__5332 (
            .O(N__28689),
            .I(N__28680));
    LocalMux I__5331 (
            .O(N__28686),
            .I(N__28672));
    LocalMux I__5330 (
            .O(N__28683),
            .I(N__28672));
    Span4Mux_v I__5329 (
            .O(N__28680),
            .I(N__28672));
    InMux I__5328 (
            .O(N__28679),
            .I(N__28669));
    Span4Mux_v I__5327 (
            .O(N__28672),
            .I(N__28664));
    LocalMux I__5326 (
            .O(N__28669),
            .I(N__28664));
    Span4Mux_h I__5325 (
            .O(N__28664),
            .I(N__28661));
    Odrv4 I__5324 (
            .O(N__28661),
            .I(\c0.data_in_frame_10_4 ));
    InMux I__5323 (
            .O(N__28658),
            .I(N__28655));
    LocalMux I__5322 (
            .O(N__28655),
            .I(N__28652));
    Span4Mux_h I__5321 (
            .O(N__28652),
            .I(N__28649));
    Odrv4 I__5320 (
            .O(N__28649),
            .I(n2563));
    CascadeMux I__5319 (
            .O(N__28646),
            .I(N__28642));
    InMux I__5318 (
            .O(N__28645),
            .I(N__28638));
    InMux I__5317 (
            .O(N__28642),
            .I(N__28635));
    InMux I__5316 (
            .O(N__28641),
            .I(N__28632));
    LocalMux I__5315 (
            .O(N__28638),
            .I(N__28628));
    LocalMux I__5314 (
            .O(N__28635),
            .I(N__28625));
    LocalMux I__5313 (
            .O(N__28632),
            .I(N__28622));
    CascadeMux I__5312 (
            .O(N__28631),
            .I(N__28618));
    Span4Mux_v I__5311 (
            .O(N__28628),
            .I(N__28615));
    Span4Mux_h I__5310 (
            .O(N__28625),
            .I(N__28610));
    Span4Mux_v I__5309 (
            .O(N__28622),
            .I(N__28610));
    InMux I__5308 (
            .O(N__28621),
            .I(N__28607));
    InMux I__5307 (
            .O(N__28618),
            .I(N__28604));
    Odrv4 I__5306 (
            .O(N__28615),
            .I(\c0.data_in_frame_7_2 ));
    Odrv4 I__5305 (
            .O(N__28610),
            .I(\c0.data_in_frame_7_2 ));
    LocalMux I__5304 (
            .O(N__28607),
            .I(\c0.data_in_frame_7_2 ));
    LocalMux I__5303 (
            .O(N__28604),
            .I(\c0.data_in_frame_7_2 ));
    InMux I__5302 (
            .O(N__28595),
            .I(N__28592));
    LocalMux I__5301 (
            .O(N__28592),
            .I(N__28588));
    InMux I__5300 (
            .O(N__28591),
            .I(N__28585));
    Span4Mux_h I__5299 (
            .O(N__28588),
            .I(N__28582));
    LocalMux I__5298 (
            .O(N__28585),
            .I(N__28579));
    Span4Mux_v I__5297 (
            .O(N__28582),
            .I(N__28576));
    Span4Mux_h I__5296 (
            .O(N__28579),
            .I(N__28573));
    Odrv4 I__5295 (
            .O(N__28576),
            .I(\c0.n8062 ));
    Odrv4 I__5294 (
            .O(N__28573),
            .I(\c0.n8062 ));
    CascadeMux I__5293 (
            .O(N__28568),
            .I(n2563_cascade_));
    InMux I__5292 (
            .O(N__28565),
            .I(N__28560));
    InMux I__5291 (
            .O(N__28564),
            .I(N__28557));
    InMux I__5290 (
            .O(N__28563),
            .I(N__28554));
    LocalMux I__5289 (
            .O(N__28560),
            .I(N__28551));
    LocalMux I__5288 (
            .O(N__28557),
            .I(N__28546));
    LocalMux I__5287 (
            .O(N__28554),
            .I(N__28546));
    Span4Mux_v I__5286 (
            .O(N__28551),
            .I(N__28541));
    Span4Mux_h I__5285 (
            .O(N__28546),
            .I(N__28541));
    Span4Mux_h I__5284 (
            .O(N__28541),
            .I(N__28538));
    Odrv4 I__5283 (
            .O(N__28538),
            .I(\c0.n9204 ));
    InMux I__5282 (
            .O(N__28535),
            .I(N__28531));
    InMux I__5281 (
            .O(N__28534),
            .I(N__28527));
    LocalMux I__5280 (
            .O(N__28531),
            .I(N__28524));
    InMux I__5279 (
            .O(N__28530),
            .I(N__28521));
    LocalMux I__5278 (
            .O(N__28527),
            .I(N__28518));
    Span4Mux_v I__5277 (
            .O(N__28524),
            .I(N__28513));
    LocalMux I__5276 (
            .O(N__28521),
            .I(N__28513));
    Span4Mux_h I__5275 (
            .O(N__28518),
            .I(N__28510));
    Span4Mux_h I__5274 (
            .O(N__28513),
            .I(N__28507));
    Odrv4 I__5273 (
            .O(N__28510),
            .I(\c0.n8890 ));
    Odrv4 I__5272 (
            .O(N__28507),
            .I(\c0.n8890 ));
    CascadeMux I__5271 (
            .O(N__28502),
            .I(\c0.n17592_cascade_ ));
    InMux I__5270 (
            .O(N__28499),
            .I(N__28496));
    LocalMux I__5269 (
            .O(N__28496),
            .I(\c0.n26 ));
    InMux I__5268 (
            .O(N__28493),
            .I(N__28488));
    InMux I__5267 (
            .O(N__28492),
            .I(N__28485));
    InMux I__5266 (
            .O(N__28491),
            .I(N__28482));
    LocalMux I__5265 (
            .O(N__28488),
            .I(N__28478));
    LocalMux I__5264 (
            .O(N__28485),
            .I(N__28473));
    LocalMux I__5263 (
            .O(N__28482),
            .I(N__28470));
    InMux I__5262 (
            .O(N__28481),
            .I(N__28467));
    Span4Mux_h I__5261 (
            .O(N__28478),
            .I(N__28464));
    InMux I__5260 (
            .O(N__28477),
            .I(N__28459));
    InMux I__5259 (
            .O(N__28476),
            .I(N__28459));
    Span4Mux_h I__5258 (
            .O(N__28473),
            .I(N__28454));
    Span4Mux_h I__5257 (
            .O(N__28470),
            .I(N__28454));
    LocalMux I__5256 (
            .O(N__28467),
            .I(N__28451));
    Span4Mux_h I__5255 (
            .O(N__28464),
            .I(N__28446));
    LocalMux I__5254 (
            .O(N__28459),
            .I(N__28446));
    Odrv4 I__5253 (
            .O(N__28454),
            .I(\c0.data_in_frame_7_5 ));
    Odrv12 I__5252 (
            .O(N__28451),
            .I(\c0.data_in_frame_7_5 ));
    Odrv4 I__5251 (
            .O(N__28446),
            .I(\c0.data_in_frame_7_5 ));
    InMux I__5250 (
            .O(N__28439),
            .I(N__28435));
    InMux I__5249 (
            .O(N__28438),
            .I(N__28429));
    LocalMux I__5248 (
            .O(N__28435),
            .I(N__28426));
    InMux I__5247 (
            .O(N__28434),
            .I(N__28423));
    InMux I__5246 (
            .O(N__28433),
            .I(N__28420));
    InMux I__5245 (
            .O(N__28432),
            .I(N__28417));
    LocalMux I__5244 (
            .O(N__28429),
            .I(N__28412));
    Span4Mux_v I__5243 (
            .O(N__28426),
            .I(N__28412));
    LocalMux I__5242 (
            .O(N__28423),
            .I(N__28409));
    LocalMux I__5241 (
            .O(N__28420),
            .I(N__28404));
    LocalMux I__5240 (
            .O(N__28417),
            .I(N__28404));
    Odrv4 I__5239 (
            .O(N__28412),
            .I(data_in_frame_8_6));
    Odrv12 I__5238 (
            .O(N__28409),
            .I(data_in_frame_8_6));
    Odrv12 I__5237 (
            .O(N__28404),
            .I(data_in_frame_8_6));
    InMux I__5236 (
            .O(N__28397),
            .I(N__28394));
    LocalMux I__5235 (
            .O(N__28394),
            .I(N__28391));
    Span4Mux_v I__5234 (
            .O(N__28391),
            .I(N__28388));
    Odrv4 I__5233 (
            .O(N__28388),
            .I(\c0.n17473 ));
    CascadeMux I__5232 (
            .O(N__28385),
            .I(N__28381));
    InMux I__5231 (
            .O(N__28384),
            .I(N__28378));
    InMux I__5230 (
            .O(N__28381),
            .I(N__28375));
    LocalMux I__5229 (
            .O(N__28378),
            .I(N__28372));
    LocalMux I__5228 (
            .O(N__28375),
            .I(N__28369));
    Span4Mux_h I__5227 (
            .O(N__28372),
            .I(N__28366));
    Span4Mux_v I__5226 (
            .O(N__28369),
            .I(N__28362));
    Span4Mux_v I__5225 (
            .O(N__28366),
            .I(N__28359));
    InMux I__5224 (
            .O(N__28365),
            .I(N__28356));
    Span4Mux_v I__5223 (
            .O(N__28362),
            .I(N__28353));
    Span4Mux_v I__5222 (
            .O(N__28359),
            .I(N__28350));
    LocalMux I__5221 (
            .O(N__28356),
            .I(\c0.data_in_4_6 ));
    Odrv4 I__5220 (
            .O(N__28353),
            .I(\c0.data_in_4_6 ));
    Odrv4 I__5219 (
            .O(N__28350),
            .I(\c0.data_in_4_6 ));
    InMux I__5218 (
            .O(N__28343),
            .I(N__28336));
    InMux I__5217 (
            .O(N__28342),
            .I(N__28332));
    InMux I__5216 (
            .O(N__28341),
            .I(N__28329));
    InMux I__5215 (
            .O(N__28340),
            .I(N__28326));
    InMux I__5214 (
            .O(N__28339),
            .I(N__28323));
    LocalMux I__5213 (
            .O(N__28336),
            .I(N__28320));
    InMux I__5212 (
            .O(N__28335),
            .I(N__28317));
    LocalMux I__5211 (
            .O(N__28332),
            .I(N__28312));
    LocalMux I__5210 (
            .O(N__28329),
            .I(N__28305));
    LocalMux I__5209 (
            .O(N__28326),
            .I(N__28305));
    LocalMux I__5208 (
            .O(N__28323),
            .I(N__28305));
    Span4Mux_v I__5207 (
            .O(N__28320),
            .I(N__28300));
    LocalMux I__5206 (
            .O(N__28317),
            .I(N__28300));
    InMux I__5205 (
            .O(N__28316),
            .I(N__28297));
    InMux I__5204 (
            .O(N__28315),
            .I(N__28294));
    Span12Mux_h I__5203 (
            .O(N__28312),
            .I(N__28291));
    Span4Mux_h I__5202 (
            .O(N__28305),
            .I(N__28286));
    Span4Mux_h I__5201 (
            .O(N__28300),
            .I(N__28286));
    LocalMux I__5200 (
            .O(N__28297),
            .I(N__28283));
    LocalMux I__5199 (
            .O(N__28294),
            .I(data_in_frame_5_7));
    Odrv12 I__5198 (
            .O(N__28291),
            .I(data_in_frame_5_7));
    Odrv4 I__5197 (
            .O(N__28286),
            .I(data_in_frame_5_7));
    Odrv4 I__5196 (
            .O(N__28283),
            .I(data_in_frame_5_7));
    InMux I__5195 (
            .O(N__28274),
            .I(N__28271));
    LocalMux I__5194 (
            .O(N__28271),
            .I(N__28268));
    Span4Mux_v I__5193 (
            .O(N__28268),
            .I(N__28265));
    Odrv4 I__5192 (
            .O(N__28265),
            .I(\c0.n9368 ));
    InMux I__5191 (
            .O(N__28262),
            .I(N__28258));
    CascadeMux I__5190 (
            .O(N__28261),
            .I(N__28255));
    LocalMux I__5189 (
            .O(N__28258),
            .I(N__28251));
    InMux I__5188 (
            .O(N__28255),
            .I(N__28248));
    InMux I__5187 (
            .O(N__28254),
            .I(N__28245));
    Span4Mux_v I__5186 (
            .O(N__28251),
            .I(N__28242));
    LocalMux I__5185 (
            .O(N__28248),
            .I(N__28239));
    LocalMux I__5184 (
            .O(N__28245),
            .I(N__28236));
    Span4Mux_h I__5183 (
            .O(N__28242),
            .I(N__28233));
    Span4Mux_h I__5182 (
            .O(N__28239),
            .I(N__28230));
    Span4Mux_h I__5181 (
            .O(N__28236),
            .I(N__28227));
    Odrv4 I__5180 (
            .O(N__28233),
            .I(\c0.n9365 ));
    Odrv4 I__5179 (
            .O(N__28230),
            .I(\c0.n9365 ));
    Odrv4 I__5178 (
            .O(N__28227),
            .I(\c0.n9365 ));
    CascadeMux I__5177 (
            .O(N__28220),
            .I(\c0.n2600_cascade_ ));
    InMux I__5176 (
            .O(N__28217),
            .I(N__28213));
    InMux I__5175 (
            .O(N__28216),
            .I(N__28210));
    LocalMux I__5174 (
            .O(N__28213),
            .I(N__28207));
    LocalMux I__5173 (
            .O(N__28210),
            .I(N__28204));
    Span4Mux_s2_h I__5172 (
            .O(N__28207),
            .I(N__28199));
    Span4Mux_v I__5171 (
            .O(N__28204),
            .I(N__28199));
    Odrv4 I__5170 (
            .O(N__28199),
            .I(\c0.n9334 ));
    InMux I__5169 (
            .O(N__28196),
            .I(N__28193));
    LocalMux I__5168 (
            .O(N__28193),
            .I(\c0.n10_adj_2493 ));
    InMux I__5167 (
            .O(N__28190),
            .I(N__28187));
    LocalMux I__5166 (
            .O(N__28187),
            .I(N__28184));
    Span4Mux_h I__5165 (
            .O(N__28184),
            .I(N__28178));
    InMux I__5164 (
            .O(N__28183),
            .I(N__28175));
    InMux I__5163 (
            .O(N__28182),
            .I(N__28171));
    InMux I__5162 (
            .O(N__28181),
            .I(N__28168));
    Span4Mux_h I__5161 (
            .O(N__28178),
            .I(N__28165));
    LocalMux I__5160 (
            .O(N__28175),
            .I(N__28162));
    InMux I__5159 (
            .O(N__28174),
            .I(N__28159));
    LocalMux I__5158 (
            .O(N__28171),
            .I(data_in_3_6));
    LocalMux I__5157 (
            .O(N__28168),
            .I(data_in_3_6));
    Odrv4 I__5156 (
            .O(N__28165),
            .I(data_in_3_6));
    Odrv4 I__5155 (
            .O(N__28162),
            .I(data_in_3_6));
    LocalMux I__5154 (
            .O(N__28159),
            .I(data_in_3_6));
    InMux I__5153 (
            .O(N__28148),
            .I(N__28145));
    LocalMux I__5152 (
            .O(N__28145),
            .I(N__28138));
    InMux I__5151 (
            .O(N__28144),
            .I(N__28131));
    InMux I__5150 (
            .O(N__28143),
            .I(N__28131));
    InMux I__5149 (
            .O(N__28142),
            .I(N__28131));
    InMux I__5148 (
            .O(N__28141),
            .I(N__28128));
    Span4Mux_v I__5147 (
            .O(N__28138),
            .I(N__28125));
    LocalMux I__5146 (
            .O(N__28131),
            .I(data_in_1_2));
    LocalMux I__5145 (
            .O(N__28128),
            .I(data_in_1_2));
    Odrv4 I__5144 (
            .O(N__28125),
            .I(data_in_1_2));
    CascadeMux I__5143 (
            .O(N__28118),
            .I(N__28114));
    CascadeMux I__5142 (
            .O(N__28117),
            .I(N__28111));
    InMux I__5141 (
            .O(N__28114),
            .I(N__28108));
    InMux I__5140 (
            .O(N__28111),
            .I(N__28105));
    LocalMux I__5139 (
            .O(N__28108),
            .I(\c0.n8572 ));
    LocalMux I__5138 (
            .O(N__28105),
            .I(\c0.n8572 ));
    InMux I__5137 (
            .O(N__28100),
            .I(N__28095));
    InMux I__5136 (
            .O(N__28099),
            .I(N__28089));
    InMux I__5135 (
            .O(N__28098),
            .I(N__28089));
    LocalMux I__5134 (
            .O(N__28095),
            .I(N__28086));
    InMux I__5133 (
            .O(N__28094),
            .I(N__28083));
    LocalMux I__5132 (
            .O(N__28089),
            .I(N__28080));
    Span4Mux_h I__5131 (
            .O(N__28086),
            .I(N__28077));
    LocalMux I__5130 (
            .O(N__28083),
            .I(N__28072));
    Span4Mux_v I__5129 (
            .O(N__28080),
            .I(N__28072));
    Odrv4 I__5128 (
            .O(N__28077),
            .I(data_in_frame_6_5));
    Odrv4 I__5127 (
            .O(N__28072),
            .I(data_in_frame_6_5));
    CascadeMux I__5126 (
            .O(N__28067),
            .I(N__28063));
    InMux I__5125 (
            .O(N__28066),
            .I(N__28059));
    InMux I__5124 (
            .O(N__28063),
            .I(N__28053));
    InMux I__5123 (
            .O(N__28062),
            .I(N__28053));
    LocalMux I__5122 (
            .O(N__28059),
            .I(N__28049));
    InMux I__5121 (
            .O(N__28058),
            .I(N__28046));
    LocalMux I__5120 (
            .O(N__28053),
            .I(N__28039));
    InMux I__5119 (
            .O(N__28052),
            .I(N__28036));
    Span4Mux_s3_h I__5118 (
            .O(N__28049),
            .I(N__28028));
    LocalMux I__5117 (
            .O(N__28046),
            .I(N__28028));
    InMux I__5116 (
            .O(N__28045),
            .I(N__28025));
    InMux I__5115 (
            .O(N__28044),
            .I(N__28016));
    InMux I__5114 (
            .O(N__28043),
            .I(N__28016));
    InMux I__5113 (
            .O(N__28042),
            .I(N__28016));
    Span4Mux_v I__5112 (
            .O(N__28039),
            .I(N__28013));
    LocalMux I__5111 (
            .O(N__28036),
            .I(N__28010));
    InMux I__5110 (
            .O(N__28035),
            .I(N__28001));
    InMux I__5109 (
            .O(N__28034),
            .I(N__27998));
    InMux I__5108 (
            .O(N__28033),
            .I(N__27995));
    Span4Mux_v I__5107 (
            .O(N__28028),
            .I(N__27990));
    LocalMux I__5106 (
            .O(N__28025),
            .I(N__27990));
    InMux I__5105 (
            .O(N__28024),
            .I(N__27985));
    InMux I__5104 (
            .O(N__28023),
            .I(N__27985));
    LocalMux I__5103 (
            .O(N__28016),
            .I(N__27978));
    Span4Mux_h I__5102 (
            .O(N__28013),
            .I(N__27978));
    Span4Mux_h I__5101 (
            .O(N__28010),
            .I(N__27978));
    InMux I__5100 (
            .O(N__28009),
            .I(N__27971));
    InMux I__5099 (
            .O(N__28008),
            .I(N__27971));
    InMux I__5098 (
            .O(N__28007),
            .I(N__27971));
    InMux I__5097 (
            .O(N__28006),
            .I(N__27964));
    InMux I__5096 (
            .O(N__28005),
            .I(N__27964));
    InMux I__5095 (
            .O(N__28004),
            .I(N__27964));
    LocalMux I__5094 (
            .O(N__28001),
            .I(\c0.n4_adj_2512 ));
    LocalMux I__5093 (
            .O(N__27998),
            .I(\c0.n4_adj_2512 ));
    LocalMux I__5092 (
            .O(N__27995),
            .I(\c0.n4_adj_2512 ));
    Odrv4 I__5091 (
            .O(N__27990),
            .I(\c0.n4_adj_2512 ));
    LocalMux I__5090 (
            .O(N__27985),
            .I(\c0.n4_adj_2512 ));
    Odrv4 I__5089 (
            .O(N__27978),
            .I(\c0.n4_adj_2512 ));
    LocalMux I__5088 (
            .O(N__27971),
            .I(\c0.n4_adj_2512 ));
    LocalMux I__5087 (
            .O(N__27964),
            .I(\c0.n4_adj_2512 ));
    InMux I__5086 (
            .O(N__27947),
            .I(N__27943));
    InMux I__5085 (
            .O(N__27946),
            .I(N__27939));
    LocalMux I__5084 (
            .O(N__27943),
            .I(N__27936));
    InMux I__5083 (
            .O(N__27942),
            .I(N__27933));
    LocalMux I__5082 (
            .O(N__27939),
            .I(N__27930));
    Span4Mux_v I__5081 (
            .O(N__27936),
            .I(N__27925));
    LocalMux I__5080 (
            .O(N__27933),
            .I(N__27925));
    Span4Mux_h I__5079 (
            .O(N__27930),
            .I(N__27922));
    Odrv4 I__5078 (
            .O(N__27925),
            .I(n2594));
    Odrv4 I__5077 (
            .O(N__27922),
            .I(n2594));
    CascadeMux I__5076 (
            .O(N__27917),
            .I(n2573_cascade_));
    InMux I__5075 (
            .O(N__27914),
            .I(N__27911));
    LocalMux I__5074 (
            .O(N__27911),
            .I(n17481));
    InMux I__5073 (
            .O(N__27908),
            .I(N__27905));
    LocalMux I__5072 (
            .O(N__27905),
            .I(N__27901));
    InMux I__5071 (
            .O(N__27904),
            .I(N__27898));
    Span4Mux_h I__5070 (
            .O(N__27901),
            .I(N__27890));
    LocalMux I__5069 (
            .O(N__27898),
            .I(N__27890));
    InMux I__5068 (
            .O(N__27897),
            .I(N__27885));
    InMux I__5067 (
            .O(N__27896),
            .I(N__27885));
    InMux I__5066 (
            .O(N__27895),
            .I(N__27882));
    Span4Mux_v I__5065 (
            .O(N__27890),
            .I(N__27877));
    LocalMux I__5064 (
            .O(N__27885),
            .I(N__27877));
    LocalMux I__5063 (
            .O(N__27882),
            .I(\c0.data_in_3_4 ));
    Odrv4 I__5062 (
            .O(N__27877),
            .I(\c0.data_in_3_4 ));
    InMux I__5061 (
            .O(N__27872),
            .I(N__27869));
    LocalMux I__5060 (
            .O(N__27869),
            .I(\c0.n17743 ));
    InMux I__5059 (
            .O(N__27866),
            .I(N__27862));
    InMux I__5058 (
            .O(N__27865),
            .I(N__27859));
    LocalMux I__5057 (
            .O(N__27862),
            .I(N__27856));
    LocalMux I__5056 (
            .O(N__27859),
            .I(N__27851));
    Span4Mux_v I__5055 (
            .O(N__27856),
            .I(N__27851));
    Span4Mux_h I__5054 (
            .O(N__27851),
            .I(N__27847));
    InMux I__5053 (
            .O(N__27850),
            .I(N__27844));
    Odrv4 I__5052 (
            .O(N__27847),
            .I(data_in_4_0));
    LocalMux I__5051 (
            .O(N__27844),
            .I(data_in_4_0));
    InMux I__5050 (
            .O(N__27839),
            .I(N__27836));
    LocalMux I__5049 (
            .O(N__27836),
            .I(N__27832));
    InMux I__5048 (
            .O(N__27835),
            .I(N__27828));
    Span4Mux_s3_h I__5047 (
            .O(N__27832),
            .I(N__27825));
    InMux I__5046 (
            .O(N__27831),
            .I(N__27820));
    LocalMux I__5045 (
            .O(N__27828),
            .I(N__27817));
    Span4Mux_h I__5044 (
            .O(N__27825),
            .I(N__27814));
    InMux I__5043 (
            .O(N__27824),
            .I(N__27811));
    InMux I__5042 (
            .O(N__27823),
            .I(N__27808));
    LocalMux I__5041 (
            .O(N__27820),
            .I(\c0.data_in_3_0 ));
    Odrv4 I__5040 (
            .O(N__27817),
            .I(\c0.data_in_3_0 ));
    Odrv4 I__5039 (
            .O(N__27814),
            .I(\c0.data_in_3_0 ));
    LocalMux I__5038 (
            .O(N__27811),
            .I(\c0.data_in_3_0 ));
    LocalMux I__5037 (
            .O(N__27808),
            .I(\c0.data_in_3_0 ));
    InMux I__5036 (
            .O(N__27797),
            .I(N__27793));
    InMux I__5035 (
            .O(N__27796),
            .I(N__27790));
    LocalMux I__5034 (
            .O(N__27793),
            .I(N__27786));
    LocalMux I__5033 (
            .O(N__27790),
            .I(N__27783));
    InMux I__5032 (
            .O(N__27789),
            .I(N__27779));
    Span4Mux_v I__5031 (
            .O(N__27786),
            .I(N__27773));
    Span4Mux_v I__5030 (
            .O(N__27783),
            .I(N__27773));
    InMux I__5029 (
            .O(N__27782),
            .I(N__27770));
    LocalMux I__5028 (
            .O(N__27779),
            .I(N__27767));
    InMux I__5027 (
            .O(N__27778),
            .I(N__27764));
    Span4Mux_h I__5026 (
            .O(N__27773),
            .I(N__27761));
    LocalMux I__5025 (
            .O(N__27770),
            .I(N__27756));
    Span12Mux_v I__5024 (
            .O(N__27767),
            .I(N__27756));
    LocalMux I__5023 (
            .O(N__27764),
            .I(data_in_1_6));
    Odrv4 I__5022 (
            .O(N__27761),
            .I(data_in_1_6));
    Odrv12 I__5021 (
            .O(N__27756),
            .I(data_in_1_6));
    InMux I__5020 (
            .O(N__27749),
            .I(N__27746));
    LocalMux I__5019 (
            .O(N__27746),
            .I(N__27743));
    Span4Mux_v I__5018 (
            .O(N__27743),
            .I(N__27737));
    InMux I__5017 (
            .O(N__27742),
            .I(N__27734));
    InMux I__5016 (
            .O(N__27741),
            .I(N__27731));
    InMux I__5015 (
            .O(N__27740),
            .I(N__27728));
    Odrv4 I__5014 (
            .O(N__27737),
            .I(data_in_0_6));
    LocalMux I__5013 (
            .O(N__27734),
            .I(data_in_0_6));
    LocalMux I__5012 (
            .O(N__27731),
            .I(data_in_0_6));
    LocalMux I__5011 (
            .O(N__27728),
            .I(data_in_0_6));
    InMux I__5010 (
            .O(N__27719),
            .I(N__27715));
    InMux I__5009 (
            .O(N__27718),
            .I(N__27711));
    LocalMux I__5008 (
            .O(N__27715),
            .I(N__27708));
    InMux I__5007 (
            .O(N__27714),
            .I(N__27704));
    LocalMux I__5006 (
            .O(N__27711),
            .I(N__27699));
    Span12Mux_v I__5005 (
            .O(N__27708),
            .I(N__27699));
    InMux I__5004 (
            .O(N__27707),
            .I(N__27696));
    LocalMux I__5003 (
            .O(N__27704),
            .I(data_in_2_6));
    Odrv12 I__5002 (
            .O(N__27699),
            .I(data_in_2_6));
    LocalMux I__5001 (
            .O(N__27696),
            .I(data_in_2_6));
    InMux I__5000 (
            .O(N__27689),
            .I(N__27686));
    LocalMux I__4999 (
            .O(N__27686),
            .I(N__27683));
    Span4Mux_h I__4998 (
            .O(N__27683),
            .I(N__27677));
    InMux I__4997 (
            .O(N__27682),
            .I(N__27672));
    InMux I__4996 (
            .O(N__27681),
            .I(N__27672));
    InMux I__4995 (
            .O(N__27680),
            .I(N__27669));
    Odrv4 I__4994 (
            .O(N__27677),
            .I(data_in_3_1));
    LocalMux I__4993 (
            .O(N__27672),
            .I(data_in_3_1));
    LocalMux I__4992 (
            .O(N__27669),
            .I(data_in_3_1));
    InMux I__4991 (
            .O(N__27662),
            .I(N__27659));
    LocalMux I__4990 (
            .O(N__27659),
            .I(N__27654));
    InMux I__4989 (
            .O(N__27658),
            .I(N__27649));
    InMux I__4988 (
            .O(N__27657),
            .I(N__27649));
    Odrv4 I__4987 (
            .O(N__27654),
            .I(data_in_9_1));
    LocalMux I__4986 (
            .O(N__27649),
            .I(data_in_9_1));
    InMux I__4985 (
            .O(N__27644),
            .I(N__27640));
    InMux I__4984 (
            .O(N__27643),
            .I(N__27637));
    LocalMux I__4983 (
            .O(N__27640),
            .I(N__27634));
    LocalMux I__4982 (
            .O(N__27637),
            .I(N__27631));
    Span4Mux_h I__4981 (
            .O(N__27634),
            .I(N__27626));
    Span4Mux_h I__4980 (
            .O(N__27631),
            .I(N__27623));
    InMux I__4979 (
            .O(N__27630),
            .I(N__27618));
    InMux I__4978 (
            .O(N__27629),
            .I(N__27618));
    Odrv4 I__4977 (
            .O(N__27626),
            .I(\c0.data_in_1_3 ));
    Odrv4 I__4976 (
            .O(N__27623),
            .I(\c0.data_in_1_3 ));
    LocalMux I__4975 (
            .O(N__27618),
            .I(\c0.data_in_1_3 ));
    InMux I__4974 (
            .O(N__27611),
            .I(N__27608));
    LocalMux I__4973 (
            .O(N__27608),
            .I(N__27605));
    Span4Mux_s2_h I__4972 (
            .O(N__27605),
            .I(N__27601));
    InMux I__4971 (
            .O(N__27604),
            .I(N__27598));
    Span4Mux_h I__4970 (
            .O(N__27601),
            .I(N__27593));
    LocalMux I__4969 (
            .O(N__27598),
            .I(N__27590));
    InMux I__4968 (
            .O(N__27597),
            .I(N__27585));
    InMux I__4967 (
            .O(N__27596),
            .I(N__27585));
    Odrv4 I__4966 (
            .O(N__27593),
            .I(\c0.data_in_0_3 ));
    Odrv4 I__4965 (
            .O(N__27590),
            .I(\c0.data_in_0_3 ));
    LocalMux I__4964 (
            .O(N__27585),
            .I(\c0.data_in_0_3 ));
    CascadeMux I__4963 (
            .O(N__27578),
            .I(N__27575));
    InMux I__4962 (
            .O(N__27575),
            .I(N__27572));
    LocalMux I__4961 (
            .O(N__27572),
            .I(N__27568));
    InMux I__4960 (
            .O(N__27571),
            .I(N__27565));
    Span4Mux_h I__4959 (
            .O(N__27568),
            .I(N__27561));
    LocalMux I__4958 (
            .O(N__27565),
            .I(N__27558));
    InMux I__4957 (
            .O(N__27564),
            .I(N__27555));
    Odrv4 I__4956 (
            .O(N__27561),
            .I(data_in_4_3));
    Odrv4 I__4955 (
            .O(N__27558),
            .I(data_in_4_3));
    LocalMux I__4954 (
            .O(N__27555),
            .I(data_in_4_3));
    InMux I__4953 (
            .O(N__27548),
            .I(N__27545));
    LocalMux I__4952 (
            .O(N__27545),
            .I(N__27542));
    Span4Mux_s2_h I__4951 (
            .O(N__27542),
            .I(N__27539));
    Span4Mux_h I__4950 (
            .O(N__27539),
            .I(N__27533));
    InMux I__4949 (
            .O(N__27538),
            .I(N__27528));
    InMux I__4948 (
            .O(N__27537),
            .I(N__27528));
    InMux I__4947 (
            .O(N__27536),
            .I(N__27525));
    Odrv4 I__4946 (
            .O(N__27533),
            .I(data_in_3_3));
    LocalMux I__4945 (
            .O(N__27528),
            .I(data_in_3_3));
    LocalMux I__4944 (
            .O(N__27525),
            .I(data_in_3_3));
    CascadeMux I__4943 (
            .O(N__27518),
            .I(N__27513));
    InMux I__4942 (
            .O(N__27517),
            .I(N__27510));
    InMux I__4941 (
            .O(N__27516),
            .I(N__27506));
    InMux I__4940 (
            .O(N__27513),
            .I(N__27503));
    LocalMux I__4939 (
            .O(N__27510),
            .I(N__27500));
    InMux I__4938 (
            .O(N__27509),
            .I(N__27497));
    LocalMux I__4937 (
            .O(N__27506),
            .I(N__27494));
    LocalMux I__4936 (
            .O(N__27503),
            .I(N__27491));
    Span4Mux_v I__4935 (
            .O(N__27500),
            .I(N__27486));
    LocalMux I__4934 (
            .O(N__27497),
            .I(N__27486));
    Span4Mux_v I__4933 (
            .O(N__27494),
            .I(N__27481));
    Span4Mux_v I__4932 (
            .O(N__27491),
            .I(N__27481));
    Span4Mux_h I__4931 (
            .O(N__27486),
            .I(N__27478));
    Odrv4 I__4930 (
            .O(N__27481),
            .I(\c0.data_in_frame_7_4 ));
    Odrv4 I__4929 (
            .O(N__27478),
            .I(\c0.data_in_frame_7_4 ));
    InMux I__4928 (
            .O(N__27473),
            .I(N__27470));
    LocalMux I__4927 (
            .O(N__27470),
            .I(N__27467));
    Span4Mux_h I__4926 (
            .O(N__27467),
            .I(N__27463));
    InMux I__4925 (
            .O(N__27466),
            .I(N__27460));
    Odrv4 I__4924 (
            .O(N__27463),
            .I(n2587));
    LocalMux I__4923 (
            .O(N__27460),
            .I(n2587));
    CascadeMux I__4922 (
            .O(N__27455),
            .I(N__27450));
    InMux I__4921 (
            .O(N__27454),
            .I(N__27447));
    InMux I__4920 (
            .O(N__27453),
            .I(N__27442));
    InMux I__4919 (
            .O(N__27450),
            .I(N__27442));
    LocalMux I__4918 (
            .O(N__27447),
            .I(\c0.data_in_7_4 ));
    LocalMux I__4917 (
            .O(N__27442),
            .I(\c0.data_in_7_4 ));
    CascadeMux I__4916 (
            .O(N__27437),
            .I(N__27434));
    InMux I__4915 (
            .O(N__27434),
            .I(N__27431));
    LocalMux I__4914 (
            .O(N__27431),
            .I(N__27428));
    Span4Mux_v I__4913 (
            .O(N__27428),
            .I(N__27423));
    InMux I__4912 (
            .O(N__27427),
            .I(N__27420));
    InMux I__4911 (
            .O(N__27426),
            .I(N__27417));
    Span4Mux_h I__4910 (
            .O(N__27423),
            .I(N__27414));
    LocalMux I__4909 (
            .O(N__27420),
            .I(\c0.data_in_6_4 ));
    LocalMux I__4908 (
            .O(N__27417),
            .I(\c0.data_in_6_4 ));
    Odrv4 I__4907 (
            .O(N__27414),
            .I(\c0.data_in_6_4 ));
    CascadeMux I__4906 (
            .O(N__27407),
            .I(N__27404));
    InMux I__4905 (
            .O(N__27404),
            .I(N__27400));
    CascadeMux I__4904 (
            .O(N__27403),
            .I(N__27397));
    LocalMux I__4903 (
            .O(N__27400),
            .I(N__27394));
    InMux I__4902 (
            .O(N__27397),
            .I(N__27391));
    Span4Mux_v I__4901 (
            .O(N__27394),
            .I(N__27384));
    LocalMux I__4900 (
            .O(N__27391),
            .I(N__27384));
    InMux I__4899 (
            .O(N__27390),
            .I(N__27379));
    InMux I__4898 (
            .O(N__27389),
            .I(N__27379));
    Span4Mux_h I__4897 (
            .O(N__27384),
            .I(N__27376));
    LocalMux I__4896 (
            .O(N__27379),
            .I(data_in_5_4));
    Odrv4 I__4895 (
            .O(N__27376),
            .I(data_in_5_4));
    InMux I__4894 (
            .O(N__27371),
            .I(N__27368));
    LocalMux I__4893 (
            .O(N__27368),
            .I(N__27365));
    Span4Mux_v I__4892 (
            .O(N__27365),
            .I(N__27361));
    InMux I__4891 (
            .O(N__27364),
            .I(N__27358));
    Span4Mux_s3_h I__4890 (
            .O(N__27361),
            .I(N__27354));
    LocalMux I__4889 (
            .O(N__27358),
            .I(N__27351));
    InMux I__4888 (
            .O(N__27357),
            .I(N__27348));
    Odrv4 I__4887 (
            .O(N__27354),
            .I(\c0.data_in_4_4 ));
    Odrv4 I__4886 (
            .O(N__27351),
            .I(\c0.data_in_4_4 ));
    LocalMux I__4885 (
            .O(N__27348),
            .I(\c0.data_in_4_4 ));
    InMux I__4884 (
            .O(N__27341),
            .I(N__27338));
    LocalMux I__4883 (
            .O(N__27338),
            .I(N__27335));
    Span4Mux_v I__4882 (
            .O(N__27335),
            .I(N__27332));
    Span4Mux_v I__4881 (
            .O(N__27332),
            .I(N__27329));
    Odrv4 I__4880 (
            .O(N__27329),
            .I(n17952));
    InMux I__4879 (
            .O(N__27326),
            .I(N__27322));
    InMux I__4878 (
            .O(N__27325),
            .I(N__27319));
    LocalMux I__4877 (
            .O(N__27322),
            .I(N__27316));
    LocalMux I__4876 (
            .O(N__27319),
            .I(N__27311));
    Span4Mux_v I__4875 (
            .O(N__27316),
            .I(N__27308));
    InMux I__4874 (
            .O(N__27315),
            .I(N__27305));
    InMux I__4873 (
            .O(N__27314),
            .I(N__27302));
    Sp12to4 I__4872 (
            .O(N__27311),
            .I(N__27299));
    Span4Mux_h I__4871 (
            .O(N__27308),
            .I(N__27296));
    LocalMux I__4870 (
            .O(N__27305),
            .I(N__27293));
    LocalMux I__4869 (
            .O(N__27302),
            .I(data_in_2_4));
    Odrv12 I__4868 (
            .O(N__27299),
            .I(data_in_2_4));
    Odrv4 I__4867 (
            .O(N__27296),
            .I(data_in_2_4));
    Odrv12 I__4866 (
            .O(N__27293),
            .I(data_in_2_4));
    InMux I__4865 (
            .O(N__27284),
            .I(N__27281));
    LocalMux I__4864 (
            .O(N__27281),
            .I(N__27277));
    InMux I__4863 (
            .O(N__27280),
            .I(N__27272));
    Span4Mux_v I__4862 (
            .O(N__27277),
            .I(N__27268));
    InMux I__4861 (
            .O(N__27276),
            .I(N__27265));
    InMux I__4860 (
            .O(N__27275),
            .I(N__27262));
    LocalMux I__4859 (
            .O(N__27272),
            .I(N__27259));
    InMux I__4858 (
            .O(N__27271),
            .I(N__27256));
    Odrv4 I__4857 (
            .O(N__27268),
            .I(data_in_2_7));
    LocalMux I__4856 (
            .O(N__27265),
            .I(data_in_2_7));
    LocalMux I__4855 (
            .O(N__27262),
            .I(data_in_2_7));
    Odrv12 I__4854 (
            .O(N__27259),
            .I(data_in_2_7));
    LocalMux I__4853 (
            .O(N__27256),
            .I(data_in_2_7));
    CascadeMux I__4852 (
            .O(N__27245),
            .I(N__27242));
    InMux I__4851 (
            .O(N__27242),
            .I(N__27239));
    LocalMux I__4850 (
            .O(N__27239),
            .I(N__27236));
    Span4Mux_v I__4849 (
            .O(N__27236),
            .I(N__27233));
    Span4Mux_h I__4848 (
            .O(N__27233),
            .I(N__27228));
    InMux I__4847 (
            .O(N__27232),
            .I(N__27225));
    InMux I__4846 (
            .O(N__27231),
            .I(N__27222));
    Odrv4 I__4845 (
            .O(N__27228),
            .I(data_in_4_7));
    LocalMux I__4844 (
            .O(N__27225),
            .I(data_in_4_7));
    LocalMux I__4843 (
            .O(N__27222),
            .I(data_in_4_7));
    CascadeMux I__4842 (
            .O(N__27215),
            .I(N__27212));
    InMux I__4841 (
            .O(N__27212),
            .I(N__27209));
    LocalMux I__4840 (
            .O(N__27209),
            .I(N__27206));
    Span4Mux_s3_h I__4839 (
            .O(N__27206),
            .I(N__27203));
    Span4Mux_v I__4838 (
            .O(N__27203),
            .I(N__27200));
    Span4Mux_h I__4837 (
            .O(N__27200),
            .I(N__27195));
    InMux I__4836 (
            .O(N__27199),
            .I(N__27192));
    InMux I__4835 (
            .O(N__27198),
            .I(N__27189));
    Odrv4 I__4834 (
            .O(N__27195),
            .I(data_in_4_5));
    LocalMux I__4833 (
            .O(N__27192),
            .I(data_in_4_5));
    LocalMux I__4832 (
            .O(N__27189),
            .I(data_in_4_5));
    InMux I__4831 (
            .O(N__27182),
            .I(N__27179));
    LocalMux I__4830 (
            .O(N__27179),
            .I(N__27176));
    Span4Mux_v I__4829 (
            .O(N__27176),
            .I(N__27169));
    InMux I__4828 (
            .O(N__27175),
            .I(N__27166));
    InMux I__4827 (
            .O(N__27174),
            .I(N__27161));
    InMux I__4826 (
            .O(N__27173),
            .I(N__27161));
    InMux I__4825 (
            .O(N__27172),
            .I(N__27158));
    Odrv4 I__4824 (
            .O(N__27169),
            .I(data_in_3_5));
    LocalMux I__4823 (
            .O(N__27166),
            .I(data_in_3_5));
    LocalMux I__4822 (
            .O(N__27161),
            .I(data_in_3_5));
    LocalMux I__4821 (
            .O(N__27158),
            .I(data_in_3_5));
    CascadeMux I__4820 (
            .O(N__27149),
            .I(\c0.n28_adj_2475_cascade_ ));
    InMux I__4819 (
            .O(N__27146),
            .I(N__27143));
    LocalMux I__4818 (
            .O(N__27143),
            .I(\c0.n8_adj_2474 ));
    InMux I__4817 (
            .O(N__27140),
            .I(N__27137));
    LocalMux I__4816 (
            .O(N__27137),
            .I(N__27134));
    Span4Mux_v I__4815 (
            .O(N__27134),
            .I(N__27130));
    InMux I__4814 (
            .O(N__27133),
            .I(N__27127));
    Odrv4 I__4813 (
            .O(N__27130),
            .I(\c0.n8559 ));
    LocalMux I__4812 (
            .O(N__27127),
            .I(\c0.n8559 ));
    InMux I__4811 (
            .O(N__27122),
            .I(N__27119));
    LocalMux I__4810 (
            .O(N__27119),
            .I(N__27116));
    Span4Mux_v I__4809 (
            .O(N__27116),
            .I(N__27112));
    InMux I__4808 (
            .O(N__27115),
            .I(N__27108));
    Span4Mux_h I__4807 (
            .O(N__27112),
            .I(N__27105));
    InMux I__4806 (
            .O(N__27111),
            .I(N__27100));
    LocalMux I__4805 (
            .O(N__27108),
            .I(N__27097));
    Sp12to4 I__4804 (
            .O(N__27105),
            .I(N__27094));
    InMux I__4803 (
            .O(N__27104),
            .I(N__27091));
    InMux I__4802 (
            .O(N__27103),
            .I(N__27088));
    LocalMux I__4801 (
            .O(N__27100),
            .I(\c0.data_in_2_0 ));
    Odrv4 I__4800 (
            .O(N__27097),
            .I(\c0.data_in_2_0 ));
    Odrv12 I__4799 (
            .O(N__27094),
            .I(\c0.data_in_2_0 ));
    LocalMux I__4798 (
            .O(N__27091),
            .I(\c0.data_in_2_0 ));
    LocalMux I__4797 (
            .O(N__27088),
            .I(\c0.data_in_2_0 ));
    InMux I__4796 (
            .O(N__27077),
            .I(N__27074));
    LocalMux I__4795 (
            .O(N__27074),
            .I(N__27070));
    InMux I__4794 (
            .O(N__27073),
            .I(N__27067));
    Span4Mux_s3_h I__4793 (
            .O(N__27070),
            .I(N__27064));
    LocalMux I__4792 (
            .O(N__27067),
            .I(N__27059));
    Span4Mux_h I__4791 (
            .O(N__27064),
            .I(N__27056));
    InMux I__4790 (
            .O(N__27063),
            .I(N__27053));
    InMux I__4789 (
            .O(N__27062),
            .I(N__27050));
    Odrv4 I__4788 (
            .O(N__27059),
            .I(data_in_0_1));
    Odrv4 I__4787 (
            .O(N__27056),
            .I(data_in_0_1));
    LocalMux I__4786 (
            .O(N__27053),
            .I(data_in_0_1));
    LocalMux I__4785 (
            .O(N__27050),
            .I(data_in_0_1));
    InMux I__4784 (
            .O(N__27041),
            .I(N__27038));
    LocalMux I__4783 (
            .O(N__27038),
            .I(N__27034));
    InMux I__4782 (
            .O(N__27037),
            .I(N__27029));
    Span4Mux_h I__4781 (
            .O(N__27034),
            .I(N__27026));
    CascadeMux I__4780 (
            .O(N__27033),
            .I(N__27023));
    InMux I__4779 (
            .O(N__27032),
            .I(N__27019));
    LocalMux I__4778 (
            .O(N__27029),
            .I(N__27016));
    Span4Mux_h I__4777 (
            .O(N__27026),
            .I(N__27013));
    InMux I__4776 (
            .O(N__27023),
            .I(N__27010));
    InMux I__4775 (
            .O(N__27022),
            .I(N__27007));
    LocalMux I__4774 (
            .O(N__27019),
            .I(data_in_1_7));
    Odrv4 I__4773 (
            .O(N__27016),
            .I(data_in_1_7));
    Odrv4 I__4772 (
            .O(N__27013),
            .I(data_in_1_7));
    LocalMux I__4771 (
            .O(N__27010),
            .I(data_in_1_7));
    LocalMux I__4770 (
            .O(N__27007),
            .I(data_in_1_7));
    InMux I__4769 (
            .O(N__26996),
            .I(N__26993));
    LocalMux I__4768 (
            .O(N__26993),
            .I(N__26990));
    Span4Mux_v I__4767 (
            .O(N__26990),
            .I(N__26986));
    InMux I__4766 (
            .O(N__26989),
            .I(N__26982));
    Span4Mux_s2_h I__4765 (
            .O(N__26986),
            .I(N__26979));
    InMux I__4764 (
            .O(N__26985),
            .I(N__26974));
    LocalMux I__4763 (
            .O(N__26982),
            .I(N__26971));
    Span4Mux_h I__4762 (
            .O(N__26979),
            .I(N__26968));
    InMux I__4761 (
            .O(N__26978),
            .I(N__26965));
    InMux I__4760 (
            .O(N__26977),
            .I(N__26962));
    LocalMux I__4759 (
            .O(N__26974),
            .I(data_in_2_5));
    Odrv4 I__4758 (
            .O(N__26971),
            .I(data_in_2_5));
    Odrv4 I__4757 (
            .O(N__26968),
            .I(data_in_2_5));
    LocalMux I__4756 (
            .O(N__26965),
            .I(data_in_2_5));
    LocalMux I__4755 (
            .O(N__26962),
            .I(data_in_2_5));
    InMux I__4754 (
            .O(N__26951),
            .I(N__26948));
    LocalMux I__4753 (
            .O(N__26948),
            .I(N__26945));
    Odrv4 I__4752 (
            .O(N__26945),
            .I(\c0.n17_adj_2486 ));
    InMux I__4751 (
            .O(N__26942),
            .I(N__26938));
    InMux I__4750 (
            .O(N__26941),
            .I(N__26935));
    LocalMux I__4749 (
            .O(N__26938),
            .I(N__26930));
    LocalMux I__4748 (
            .O(N__26935),
            .I(N__26926));
    InMux I__4747 (
            .O(N__26934),
            .I(N__26922));
    InMux I__4746 (
            .O(N__26933),
            .I(N__26919));
    Span4Mux_v I__4745 (
            .O(N__26930),
            .I(N__26916));
    InMux I__4744 (
            .O(N__26929),
            .I(N__26913));
    Span4Mux_v I__4743 (
            .O(N__26926),
            .I(N__26910));
    InMux I__4742 (
            .O(N__26925),
            .I(N__26907));
    LocalMux I__4741 (
            .O(N__26922),
            .I(N__26902));
    LocalMux I__4740 (
            .O(N__26919),
            .I(N__26895));
    Span4Mux_s1_h I__4739 (
            .O(N__26916),
            .I(N__26895));
    LocalMux I__4738 (
            .O(N__26913),
            .I(N__26895));
    Sp12to4 I__4737 (
            .O(N__26910),
            .I(N__26890));
    LocalMux I__4736 (
            .O(N__26907),
            .I(N__26890));
    InMux I__4735 (
            .O(N__26906),
            .I(N__26887));
    InMux I__4734 (
            .O(N__26905),
            .I(N__26884));
    Span4Mux_v I__4733 (
            .O(N__26902),
            .I(N__26879));
    Span4Mux_v I__4732 (
            .O(N__26895),
            .I(N__26879));
    Odrv12 I__4731 (
            .O(N__26890),
            .I(\c0.n134 ));
    LocalMux I__4730 (
            .O(N__26887),
            .I(\c0.n134 ));
    LocalMux I__4729 (
            .O(N__26884),
            .I(\c0.n134 ));
    Odrv4 I__4728 (
            .O(N__26879),
            .I(\c0.n134 ));
    CascadeMux I__4727 (
            .O(N__26870),
            .I(\c0.n18531_cascade_ ));
    InMux I__4726 (
            .O(N__26867),
            .I(N__26864));
    LocalMux I__4725 (
            .O(N__26864),
            .I(N__26860));
    InMux I__4724 (
            .O(N__26863),
            .I(N__26857));
    Span4Mux_s2_v I__4723 (
            .O(N__26860),
            .I(N__26854));
    LocalMux I__4722 (
            .O(N__26857),
            .I(data_out_frame2_5_4));
    Odrv4 I__4721 (
            .O(N__26854),
            .I(data_out_frame2_5_4));
    CascadeMux I__4720 (
            .O(N__26849),
            .I(\c0.n17955_cascade_ ));
    InMux I__4719 (
            .O(N__26846),
            .I(N__26835));
    InMux I__4718 (
            .O(N__26845),
            .I(N__26835));
    InMux I__4717 (
            .O(N__26844),
            .I(N__26828));
    InMux I__4716 (
            .O(N__26843),
            .I(N__26828));
    InMux I__4715 (
            .O(N__26842),
            .I(N__26823));
    InMux I__4714 (
            .O(N__26841),
            .I(N__26818));
    InMux I__4713 (
            .O(N__26840),
            .I(N__26818));
    LocalMux I__4712 (
            .O(N__26835),
            .I(N__26815));
    InMux I__4711 (
            .O(N__26834),
            .I(N__26812));
    InMux I__4710 (
            .O(N__26833),
            .I(N__26809));
    LocalMux I__4709 (
            .O(N__26828),
            .I(N__26806));
    InMux I__4708 (
            .O(N__26827),
            .I(N__26801));
    InMux I__4707 (
            .O(N__26826),
            .I(N__26801));
    LocalMux I__4706 (
            .O(N__26823),
            .I(N__26795));
    LocalMux I__4705 (
            .O(N__26818),
            .I(N__26786));
    Span4Mux_h I__4704 (
            .O(N__26815),
            .I(N__26786));
    LocalMux I__4703 (
            .O(N__26812),
            .I(N__26786));
    LocalMux I__4702 (
            .O(N__26809),
            .I(N__26786));
    Span4Mux_v I__4701 (
            .O(N__26806),
            .I(N__26775));
    LocalMux I__4700 (
            .O(N__26801),
            .I(N__26775));
    InMux I__4699 (
            .O(N__26800),
            .I(N__26768));
    InMux I__4698 (
            .O(N__26799),
            .I(N__26768));
    InMux I__4697 (
            .O(N__26798),
            .I(N__26768));
    Span4Mux_v I__4696 (
            .O(N__26795),
            .I(N__26765));
    Span4Mux_v I__4695 (
            .O(N__26786),
            .I(N__26762));
    InMux I__4694 (
            .O(N__26785),
            .I(N__26759));
    InMux I__4693 (
            .O(N__26784),
            .I(N__26755));
    InMux I__4692 (
            .O(N__26783),
            .I(N__26750));
    InMux I__4691 (
            .O(N__26782),
            .I(N__26750));
    InMux I__4690 (
            .O(N__26781),
            .I(N__26745));
    InMux I__4689 (
            .O(N__26780),
            .I(N__26745));
    Span4Mux_h I__4688 (
            .O(N__26775),
            .I(N__26742));
    LocalMux I__4687 (
            .O(N__26768),
            .I(N__26733));
    Sp12to4 I__4686 (
            .O(N__26765),
            .I(N__26733));
    Sp12to4 I__4685 (
            .O(N__26762),
            .I(N__26733));
    LocalMux I__4684 (
            .O(N__26759),
            .I(N__26733));
    InMux I__4683 (
            .O(N__26758),
            .I(N__26730));
    LocalMux I__4682 (
            .O(N__26755),
            .I(N__26719));
    LocalMux I__4681 (
            .O(N__26750),
            .I(N__26719));
    LocalMux I__4680 (
            .O(N__26745),
            .I(N__26719));
    Sp12to4 I__4679 (
            .O(N__26742),
            .I(N__26719));
    Span12Mux_h I__4678 (
            .O(N__26733),
            .I(N__26719));
    LocalMux I__4677 (
            .O(N__26730),
            .I(\c0.byte_transmit_counter2_2 ));
    Odrv12 I__4676 (
            .O(N__26719),
            .I(\c0.byte_transmit_counter2_2 ));
    InMux I__4675 (
            .O(N__26714),
            .I(N__26711));
    LocalMux I__4674 (
            .O(N__26711),
            .I(N__26707));
    InMux I__4673 (
            .O(N__26710),
            .I(N__26704));
    Span4Mux_s2_v I__4672 (
            .O(N__26707),
            .I(N__26701));
    LocalMux I__4671 (
            .O(N__26704),
            .I(\c0.data_out_frame2_0_4 ));
    Odrv4 I__4670 (
            .O(N__26701),
            .I(\c0.data_out_frame2_0_4 ));
    CascadeMux I__4669 (
            .O(N__26696),
            .I(\c0.n18456_cascade_ ));
    InMux I__4668 (
            .O(N__26693),
            .I(N__26690));
    LocalMux I__4667 (
            .O(N__26690),
            .I(\c0.n18447 ));
    CascadeMux I__4666 (
            .O(N__26687),
            .I(\c0.n18459_cascade_ ));
    InMux I__4665 (
            .O(N__26684),
            .I(N__26681));
    LocalMux I__4664 (
            .O(N__26681),
            .I(\c0.n22_adj_2525 ));
    InMux I__4663 (
            .O(N__26678),
            .I(N__26669));
    InMux I__4662 (
            .O(N__26677),
            .I(N__26654));
    InMux I__4661 (
            .O(N__26676),
            .I(N__26654));
    InMux I__4660 (
            .O(N__26675),
            .I(N__26654));
    InMux I__4659 (
            .O(N__26674),
            .I(N__26647));
    InMux I__4658 (
            .O(N__26673),
            .I(N__26647));
    InMux I__4657 (
            .O(N__26672),
            .I(N__26647));
    LocalMux I__4656 (
            .O(N__26669),
            .I(N__26644));
    InMux I__4655 (
            .O(N__26668),
            .I(N__26641));
    CascadeMux I__4654 (
            .O(N__26667),
            .I(N__26638));
    InMux I__4653 (
            .O(N__26666),
            .I(N__26635));
    InMux I__4652 (
            .O(N__26665),
            .I(N__26628));
    InMux I__4651 (
            .O(N__26664),
            .I(N__26628));
    InMux I__4650 (
            .O(N__26663),
            .I(N__26628));
    CascadeMux I__4649 (
            .O(N__26662),
            .I(N__26621));
    InMux I__4648 (
            .O(N__26661),
            .I(N__26613));
    LocalMux I__4647 (
            .O(N__26654),
            .I(N__26608));
    LocalMux I__4646 (
            .O(N__26647),
            .I(N__26608));
    Span4Mux_h I__4645 (
            .O(N__26644),
            .I(N__26603));
    LocalMux I__4644 (
            .O(N__26641),
            .I(N__26603));
    InMux I__4643 (
            .O(N__26638),
            .I(N__26599));
    LocalMux I__4642 (
            .O(N__26635),
            .I(N__26594));
    LocalMux I__4641 (
            .O(N__26628),
            .I(N__26594));
    InMux I__4640 (
            .O(N__26627),
            .I(N__26589));
    InMux I__4639 (
            .O(N__26626),
            .I(N__26589));
    InMux I__4638 (
            .O(N__26625),
            .I(N__26584));
    InMux I__4637 (
            .O(N__26624),
            .I(N__26584));
    InMux I__4636 (
            .O(N__26621),
            .I(N__26581));
    InMux I__4635 (
            .O(N__26620),
            .I(N__26576));
    InMux I__4634 (
            .O(N__26619),
            .I(N__26576));
    InMux I__4633 (
            .O(N__26618),
            .I(N__26569));
    InMux I__4632 (
            .O(N__26617),
            .I(N__26569));
    InMux I__4631 (
            .O(N__26616),
            .I(N__26569));
    LocalMux I__4630 (
            .O(N__26613),
            .I(N__26564));
    Span4Mux_h I__4629 (
            .O(N__26608),
            .I(N__26564));
    Span4Mux_h I__4628 (
            .O(N__26603),
            .I(N__26561));
    InMux I__4627 (
            .O(N__26602),
            .I(N__26558));
    LocalMux I__4626 (
            .O(N__26599),
            .I(N__26555));
    Span12Mux_s10_v I__4625 (
            .O(N__26594),
            .I(N__26552));
    LocalMux I__4624 (
            .O(N__26589),
            .I(N__26537));
    LocalMux I__4623 (
            .O(N__26584),
            .I(N__26537));
    LocalMux I__4622 (
            .O(N__26581),
            .I(N__26537));
    LocalMux I__4621 (
            .O(N__26576),
            .I(N__26537));
    LocalMux I__4620 (
            .O(N__26569),
            .I(N__26537));
    Sp12to4 I__4619 (
            .O(N__26564),
            .I(N__26537));
    Sp12to4 I__4618 (
            .O(N__26561),
            .I(N__26537));
    LocalMux I__4617 (
            .O(N__26558),
            .I(\c0.byte_transmit_counter2_3 ));
    Odrv4 I__4616 (
            .O(N__26555),
            .I(\c0.byte_transmit_counter2_3 ));
    Odrv12 I__4615 (
            .O(N__26552),
            .I(\c0.byte_transmit_counter2_3 ));
    Odrv12 I__4614 (
            .O(N__26537),
            .I(\c0.byte_transmit_counter2_3 ));
    CascadeMux I__4613 (
            .O(N__26528),
            .I(\c0.n15_cascade_ ));
    InMux I__4612 (
            .O(N__26525),
            .I(N__26522));
    LocalMux I__4611 (
            .O(N__26522),
            .I(N__26515));
    InMux I__4610 (
            .O(N__26521),
            .I(N__26512));
    InMux I__4609 (
            .O(N__26520),
            .I(N__26509));
    InMux I__4608 (
            .O(N__26519),
            .I(N__26505));
    InMux I__4607 (
            .O(N__26518),
            .I(N__26502));
    Span4Mux_s2_v I__4606 (
            .O(N__26515),
            .I(N__26495));
    LocalMux I__4605 (
            .O(N__26512),
            .I(N__26495));
    LocalMux I__4604 (
            .O(N__26509),
            .I(N__26492));
    InMux I__4603 (
            .O(N__26508),
            .I(N__26489));
    LocalMux I__4602 (
            .O(N__26505),
            .I(N__26486));
    LocalMux I__4601 (
            .O(N__26502),
            .I(N__26483));
    InMux I__4600 (
            .O(N__26501),
            .I(N__26480));
    InMux I__4599 (
            .O(N__26500),
            .I(N__26477));
    Span4Mux_v I__4598 (
            .O(N__26495),
            .I(N__26473));
    Span4Mux_h I__4597 (
            .O(N__26492),
            .I(N__26466));
    LocalMux I__4596 (
            .O(N__26489),
            .I(N__26466));
    Span4Mux_s2_v I__4595 (
            .O(N__26486),
            .I(N__26466));
    Span4Mux_s3_v I__4594 (
            .O(N__26483),
            .I(N__26459));
    LocalMux I__4593 (
            .O(N__26480),
            .I(N__26459));
    LocalMux I__4592 (
            .O(N__26477),
            .I(N__26459));
    InMux I__4591 (
            .O(N__26476),
            .I(N__26456));
    Span4Mux_h I__4590 (
            .O(N__26473),
            .I(N__26450));
    Span4Mux_v I__4589 (
            .O(N__26466),
            .I(N__26450));
    Span4Mux_v I__4588 (
            .O(N__26459),
            .I(N__26445));
    LocalMux I__4587 (
            .O(N__26456),
            .I(N__26445));
    InMux I__4586 (
            .O(N__26455),
            .I(N__26442));
    Span4Mux_v I__4585 (
            .O(N__26450),
            .I(N__26439));
    Odrv4 I__4584 (
            .O(N__26445),
            .I(\c0.byte_transmit_counter2_4 ));
    LocalMux I__4583 (
            .O(N__26442),
            .I(\c0.byte_transmit_counter2_4 ));
    Odrv4 I__4582 (
            .O(N__26439),
            .I(\c0.byte_transmit_counter2_4 ));
    CascadeMux I__4581 (
            .O(N__26432),
            .I(N__26429));
    InMux I__4580 (
            .O(N__26429),
            .I(N__26426));
    LocalMux I__4579 (
            .O(N__26426),
            .I(N__26423));
    Span4Mux_h I__4578 (
            .O(N__26423),
            .I(N__26420));
    Odrv4 I__4577 (
            .O(N__26420),
            .I(\c0.tx2.r_Tx_Data_4 ));
    CEMux I__4576 (
            .O(N__26417),
            .I(N__26413));
    CEMux I__4575 (
            .O(N__26416),
            .I(N__26410));
    LocalMux I__4574 (
            .O(N__26413),
            .I(N__26406));
    LocalMux I__4573 (
            .O(N__26410),
            .I(N__26401));
    CEMux I__4572 (
            .O(N__26409),
            .I(N__26397));
    Span4Mux_v I__4571 (
            .O(N__26406),
            .I(N__26394));
    CEMux I__4570 (
            .O(N__26405),
            .I(N__26391));
    CEMux I__4569 (
            .O(N__26404),
            .I(N__26388));
    Span4Mux_h I__4568 (
            .O(N__26401),
            .I(N__26385));
    CEMux I__4567 (
            .O(N__26400),
            .I(N__26382));
    LocalMux I__4566 (
            .O(N__26397),
            .I(N__26379));
    Sp12to4 I__4565 (
            .O(N__26394),
            .I(N__26374));
    LocalMux I__4564 (
            .O(N__26391),
            .I(N__26371));
    LocalMux I__4563 (
            .O(N__26388),
            .I(N__26368));
    Span4Mux_h I__4562 (
            .O(N__26385),
            .I(N__26365));
    LocalMux I__4561 (
            .O(N__26382),
            .I(N__26362));
    Span4Mux_s2_h I__4560 (
            .O(N__26379),
            .I(N__26359));
    CEMux I__4559 (
            .O(N__26378),
            .I(N__26356));
    CEMux I__4558 (
            .O(N__26377),
            .I(N__26353));
    Span12Mux_s1_h I__4557 (
            .O(N__26374),
            .I(N__26350));
    Span4Mux_v I__4556 (
            .O(N__26371),
            .I(N__26347));
    Span4Mux_s1_v I__4555 (
            .O(N__26368),
            .I(N__26344));
    Span4Mux_s1_h I__4554 (
            .O(N__26365),
            .I(N__26341));
    Sp12to4 I__4553 (
            .O(N__26362),
            .I(N__26338));
    Span4Mux_v I__4552 (
            .O(N__26359),
            .I(N__26335));
    LocalMux I__4551 (
            .O(N__26356),
            .I(\c0.tx2.n7727 ));
    LocalMux I__4550 (
            .O(N__26353),
            .I(\c0.tx2.n7727 ));
    Odrv12 I__4549 (
            .O(N__26350),
            .I(\c0.tx2.n7727 ));
    Odrv4 I__4548 (
            .O(N__26347),
            .I(\c0.tx2.n7727 ));
    Odrv4 I__4547 (
            .O(N__26344),
            .I(\c0.tx2.n7727 ));
    Odrv4 I__4546 (
            .O(N__26341),
            .I(\c0.tx2.n7727 ));
    Odrv12 I__4545 (
            .O(N__26338),
            .I(\c0.tx2.n7727 ));
    Odrv4 I__4544 (
            .O(N__26335),
            .I(\c0.tx2.n7727 ));
    InMux I__4543 (
            .O(N__26318),
            .I(N__26315));
    LocalMux I__4542 (
            .O(N__26315),
            .I(N__26312));
    Span4Mux_s2_v I__4541 (
            .O(N__26312),
            .I(N__26309));
    Odrv4 I__4540 (
            .O(N__26309),
            .I(n224));
    InMux I__4539 (
            .O(N__26306),
            .I(N__26303));
    LocalMux I__4538 (
            .O(N__26303),
            .I(n226));
    InMux I__4537 (
            .O(N__26300),
            .I(N__26297));
    LocalMux I__4536 (
            .O(N__26297),
            .I(n221));
    InMux I__4535 (
            .O(N__26294),
            .I(N__26291));
    LocalMux I__4534 (
            .O(N__26291),
            .I(n223));
    InMux I__4533 (
            .O(N__26288),
            .I(N__26285));
    LocalMux I__4532 (
            .O(N__26285),
            .I(\c0.rx.n17999 ));
    InMux I__4531 (
            .O(N__26282),
            .I(N__26279));
    LocalMux I__4530 (
            .O(N__26279),
            .I(N__26276));
    Odrv4 I__4529 (
            .O(N__26276),
            .I(\c0.n18444 ));
    InMux I__4528 (
            .O(N__26273),
            .I(N__26270));
    LocalMux I__4527 (
            .O(N__26270),
            .I(N__26267));
    Odrv12 I__4526 (
            .O(N__26267),
            .I(\c0.n9 ));
    InMux I__4525 (
            .O(N__26264),
            .I(N__26261));
    LocalMux I__4524 (
            .O(N__26261),
            .I(N__26257));
    InMux I__4523 (
            .O(N__26260),
            .I(N__26254));
    Span4Mux_h I__4522 (
            .O(N__26257),
            .I(N__26251));
    LocalMux I__4521 (
            .O(N__26254),
            .I(N__26246));
    Span4Mux_v I__4520 (
            .O(N__26251),
            .I(N__26246));
    Odrv4 I__4519 (
            .O(N__26246),
            .I(data_out_frame2_18_4));
    CascadeMux I__4518 (
            .O(N__26243),
            .I(N__26240));
    InMux I__4517 (
            .O(N__26240),
            .I(N__26237));
    LocalMux I__4516 (
            .O(N__26237),
            .I(N__26234));
    Span4Mux_v I__4515 (
            .O(N__26234),
            .I(N__26231));
    Span4Mux_v I__4514 (
            .O(N__26231),
            .I(N__26228));
    Odrv4 I__4513 (
            .O(N__26228),
            .I(\c0.data_out_frame2_19_4 ));
    InMux I__4512 (
            .O(N__26225),
            .I(N__26222));
    LocalMux I__4511 (
            .O(N__26222),
            .I(N__26218));
    InMux I__4510 (
            .O(N__26221),
            .I(N__26215));
    Span4Mux_s3_v I__4509 (
            .O(N__26218),
            .I(N__26212));
    LocalMux I__4508 (
            .O(N__26215),
            .I(data_out_frame2_16_4));
    Odrv4 I__4507 (
            .O(N__26212),
            .I(data_out_frame2_16_4));
    CascadeMux I__4506 (
            .O(N__26207),
            .I(\c0.n18528_cascade_ ));
    InMux I__4505 (
            .O(N__26204),
            .I(N__26201));
    LocalMux I__4504 (
            .O(N__26201),
            .I(N__26197));
    InMux I__4503 (
            .O(N__26200),
            .I(N__26194));
    Span12Mux_s6_v I__4502 (
            .O(N__26197),
            .I(N__26191));
    LocalMux I__4501 (
            .O(N__26194),
            .I(data_out_frame2_17_4));
    Odrv12 I__4500 (
            .O(N__26191),
            .I(data_out_frame2_17_4));
    InMux I__4499 (
            .O(N__26186),
            .I(N__26182));
    InMux I__4498 (
            .O(N__26185),
            .I(N__26177));
    LocalMux I__4497 (
            .O(N__26182),
            .I(N__26174));
    InMux I__4496 (
            .O(N__26181),
            .I(N__26171));
    CascadeMux I__4495 (
            .O(N__26180),
            .I(N__26164));
    LocalMux I__4494 (
            .O(N__26177),
            .I(N__26161));
    Span4Mux_h I__4493 (
            .O(N__26174),
            .I(N__26156));
    LocalMux I__4492 (
            .O(N__26171),
            .I(N__26156));
    InMux I__4491 (
            .O(N__26170),
            .I(N__26153));
    InMux I__4490 (
            .O(N__26169),
            .I(N__26144));
    InMux I__4489 (
            .O(N__26168),
            .I(N__26144));
    InMux I__4488 (
            .O(N__26167),
            .I(N__26144));
    InMux I__4487 (
            .O(N__26164),
            .I(N__26144));
    Odrv4 I__4486 (
            .O(N__26161),
            .I(r_Bit_Index_1_adj_2636));
    Odrv4 I__4485 (
            .O(N__26156),
            .I(r_Bit_Index_1_adj_2636));
    LocalMux I__4484 (
            .O(N__26153),
            .I(r_Bit_Index_1_adj_2636));
    LocalMux I__4483 (
            .O(N__26144),
            .I(r_Bit_Index_1_adj_2636));
    InMux I__4482 (
            .O(N__26135),
            .I(N__26132));
    LocalMux I__4481 (
            .O(N__26132),
            .I(N__26126));
    InMux I__4480 (
            .O(N__26131),
            .I(N__26121));
    InMux I__4479 (
            .O(N__26130),
            .I(N__26121));
    CascadeMux I__4478 (
            .O(N__26129),
            .I(N__26115));
    Span4Mux_h I__4477 (
            .O(N__26126),
            .I(N__26110));
    LocalMux I__4476 (
            .O(N__26121),
            .I(N__26110));
    InMux I__4475 (
            .O(N__26120),
            .I(N__26103));
    InMux I__4474 (
            .O(N__26119),
            .I(N__26103));
    InMux I__4473 (
            .O(N__26118),
            .I(N__26103));
    InMux I__4472 (
            .O(N__26115),
            .I(N__26100));
    Odrv4 I__4471 (
            .O(N__26110),
            .I(r_Bit_Index_0_adj_2637));
    LocalMux I__4470 (
            .O(N__26103),
            .I(r_Bit_Index_0_adj_2637));
    LocalMux I__4469 (
            .O(N__26100),
            .I(r_Bit_Index_0_adj_2637));
    CascadeMux I__4468 (
            .O(N__26093),
            .I(N__26090));
    InMux I__4467 (
            .O(N__26090),
            .I(N__26087));
    LocalMux I__4466 (
            .O(N__26087),
            .I(n4980));
    InMux I__4465 (
            .O(N__26084),
            .I(bfn_6_30_0_));
    InMux I__4464 (
            .O(N__26081),
            .I(N__26078));
    LocalMux I__4463 (
            .O(N__26078),
            .I(n225));
    InMux I__4462 (
            .O(N__26075),
            .I(\c0.rx.n16365 ));
    InMux I__4461 (
            .O(N__26072),
            .I(\c0.rx.n16366 ));
    InMux I__4460 (
            .O(N__26069),
            .I(\c0.rx.n16367 ));
    InMux I__4459 (
            .O(N__26066),
            .I(\c0.rx.n16368 ));
    InMux I__4458 (
            .O(N__26063),
            .I(\c0.rx.n16369 ));
    InMux I__4457 (
            .O(N__26060),
            .I(\c0.rx.n16370 ));
    InMux I__4456 (
            .O(N__26057),
            .I(\c0.rx.n16371 ));
    CascadeMux I__4455 (
            .O(N__26054),
            .I(\c0.n18375_cascade_ ));
    InMux I__4454 (
            .O(N__26051),
            .I(N__26048));
    LocalMux I__4453 (
            .O(N__26048),
            .I(N__26045));
    Span4Mux_v I__4452 (
            .O(N__26045),
            .I(N__26042));
    Odrv4 I__4451 (
            .O(N__26042),
            .I(\c0.tx2.r_Tx_Data_3 ));
    InMux I__4450 (
            .O(N__26039),
            .I(N__26036));
    LocalMux I__4449 (
            .O(N__26036),
            .I(N__26032));
    InMux I__4448 (
            .O(N__26035),
            .I(N__26029));
    Span4Mux_h I__4447 (
            .O(N__26032),
            .I(N__26026));
    LocalMux I__4446 (
            .O(N__26029),
            .I(data_out_frame2_18_3));
    Odrv4 I__4445 (
            .O(N__26026),
            .I(data_out_frame2_18_3));
    CascadeMux I__4444 (
            .O(N__26021),
            .I(N__26018));
    InMux I__4443 (
            .O(N__26018),
            .I(N__26015));
    LocalMux I__4442 (
            .O(N__26015),
            .I(N__26012));
    Span4Mux_h I__4441 (
            .O(N__26012),
            .I(N__26009));
    Span4Mux_v I__4440 (
            .O(N__26009),
            .I(N__26006));
    Odrv4 I__4439 (
            .O(N__26006),
            .I(\c0.data_out_frame2_19_3 ));
    InMux I__4438 (
            .O(N__26003),
            .I(N__26000));
    LocalMux I__4437 (
            .O(N__26000),
            .I(N__25996));
    InMux I__4436 (
            .O(N__25999),
            .I(N__25993));
    Span4Mux_h I__4435 (
            .O(N__25996),
            .I(N__25990));
    LocalMux I__4434 (
            .O(N__25993),
            .I(data_out_frame2_16_3));
    Odrv4 I__4433 (
            .O(N__25990),
            .I(data_out_frame2_16_3));
    CascadeMux I__4432 (
            .O(N__25985),
            .I(\c0.n18510_cascade_ ));
    InMux I__4431 (
            .O(N__25982),
            .I(N__25979));
    LocalMux I__4430 (
            .O(N__25979),
            .I(N__25975));
    InMux I__4429 (
            .O(N__25978),
            .I(N__25972));
    Span4Mux_h I__4428 (
            .O(N__25975),
            .I(N__25969));
    LocalMux I__4427 (
            .O(N__25972),
            .I(data_out_frame2_17_3));
    Odrv4 I__4426 (
            .O(N__25969),
            .I(data_out_frame2_17_3));
    InMux I__4425 (
            .O(N__25964),
            .I(N__25961));
    LocalMux I__4424 (
            .O(N__25961),
            .I(N__25958));
    Span4Mux_v I__4423 (
            .O(N__25958),
            .I(N__25955));
    Odrv4 I__4422 (
            .O(N__25955),
            .I(\c0.data_out_frame2_20_3 ));
    CascadeMux I__4421 (
            .O(N__25952),
            .I(\c0.n18513_cascade_ ));
    InMux I__4420 (
            .O(N__25949),
            .I(N__25946));
    LocalMux I__4419 (
            .O(N__25946),
            .I(\c0.n22_adj_2527 ));
    InMux I__4418 (
            .O(N__25943),
            .I(N__25939));
    CascadeMux I__4417 (
            .O(N__25942),
            .I(N__25936));
    LocalMux I__4416 (
            .O(N__25939),
            .I(N__25932));
    InMux I__4415 (
            .O(N__25936),
            .I(N__25927));
    InMux I__4414 (
            .O(N__25935),
            .I(N__25927));
    Span4Mux_h I__4413 (
            .O(N__25932),
            .I(N__25923));
    LocalMux I__4412 (
            .O(N__25927),
            .I(N__25920));
    InMux I__4411 (
            .O(N__25926),
            .I(N__25917));
    Odrv4 I__4410 (
            .O(N__25923),
            .I(n9652));
    Odrv4 I__4409 (
            .O(N__25920),
            .I(n9652));
    LocalMux I__4408 (
            .O(N__25917),
            .I(n9652));
    InMux I__4407 (
            .O(N__25910),
            .I(N__25907));
    LocalMux I__4406 (
            .O(N__25907),
            .I(N__25902));
    InMux I__4405 (
            .O(N__25906),
            .I(N__25897));
    InMux I__4404 (
            .O(N__25905),
            .I(N__25897));
    Span4Mux_h I__4403 (
            .O(N__25902),
            .I(N__25892));
    LocalMux I__4402 (
            .O(N__25897),
            .I(N__25892));
    Odrv4 I__4401 (
            .O(N__25892),
            .I(n9922));
    InMux I__4400 (
            .O(N__25889),
            .I(N__25885));
    InMux I__4399 (
            .O(N__25888),
            .I(N__25881));
    LocalMux I__4398 (
            .O(N__25885),
            .I(N__25878));
    InMux I__4397 (
            .O(N__25884),
            .I(N__25875));
    LocalMux I__4396 (
            .O(N__25881),
            .I(N__25872));
    Sp12to4 I__4395 (
            .O(N__25878),
            .I(N__25866));
    LocalMux I__4394 (
            .O(N__25875),
            .I(N__25866));
    Span4Mux_s3_v I__4393 (
            .O(N__25872),
            .I(N__25863));
    InMux I__4392 (
            .O(N__25871),
            .I(N__25860));
    Span12Mux_s3_v I__4391 (
            .O(N__25866),
            .I(N__25857));
    Span4Mux_h I__4390 (
            .O(N__25863),
            .I(N__25854));
    LocalMux I__4389 (
            .O(N__25860),
            .I(r_Bit_Index_2_adj_2635));
    Odrv12 I__4388 (
            .O(N__25857),
            .I(r_Bit_Index_2_adj_2635));
    Odrv4 I__4387 (
            .O(N__25854),
            .I(r_Bit_Index_2_adj_2635));
    CascadeMux I__4386 (
            .O(N__25847),
            .I(N__25844));
    InMux I__4385 (
            .O(N__25844),
            .I(N__25841));
    LocalMux I__4384 (
            .O(N__25841),
            .I(N__25838));
    Odrv4 I__4383 (
            .O(N__25838),
            .I(\c0.n17559 ));
    InMux I__4382 (
            .O(N__25835),
            .I(N__25832));
    LocalMux I__4381 (
            .O(N__25832),
            .I(N__25828));
    InMux I__4380 (
            .O(N__25831),
            .I(N__25825));
    Span4Mux_v I__4379 (
            .O(N__25828),
            .I(N__25822));
    LocalMux I__4378 (
            .O(N__25825),
            .I(N__25819));
    Span4Mux_h I__4377 (
            .O(N__25822),
            .I(N__25816));
    Odrv4 I__4376 (
            .O(N__25819),
            .I(n9135));
    Odrv4 I__4375 (
            .O(N__25816),
            .I(n9135));
    InMux I__4374 (
            .O(N__25811),
            .I(N__25807));
    InMux I__4373 (
            .O(N__25810),
            .I(N__25804));
    LocalMux I__4372 (
            .O(N__25807),
            .I(N__25801));
    LocalMux I__4371 (
            .O(N__25804),
            .I(\c0.data_out_frame2_0_3 ));
    Odrv4 I__4370 (
            .O(N__25801),
            .I(\c0.data_out_frame2_0_3 ));
    InMux I__4369 (
            .O(N__25796),
            .I(N__25793));
    LocalMux I__4368 (
            .O(N__25793),
            .I(\c0.n18082 ));
    InMux I__4367 (
            .O(N__25790),
            .I(N__25786));
    InMux I__4366 (
            .O(N__25789),
            .I(N__25783));
    LocalMux I__4365 (
            .O(N__25786),
            .I(\c0.n14631 ));
    LocalMux I__4364 (
            .O(N__25783),
            .I(\c0.n14631 ));
    InMux I__4363 (
            .O(N__25778),
            .I(N__25774));
    InMux I__4362 (
            .O(N__25777),
            .I(N__25771));
    LocalMux I__4361 (
            .O(N__25774),
            .I(data_out_frame2_12_3));
    LocalMux I__4360 (
            .O(N__25771),
            .I(data_out_frame2_12_3));
    InMux I__4359 (
            .O(N__25766),
            .I(N__25760));
    InMux I__4358 (
            .O(N__25765),
            .I(N__25760));
    LocalMux I__4357 (
            .O(N__25760),
            .I(data_in_20_2));
    InMux I__4356 (
            .O(N__25757),
            .I(N__25754));
    LocalMux I__4355 (
            .O(N__25754),
            .I(\c0.n17815 ));
    CascadeMux I__4354 (
            .O(N__25751),
            .I(N__25748));
    InMux I__4353 (
            .O(N__25748),
            .I(N__25745));
    LocalMux I__4352 (
            .O(N__25745),
            .I(\c0.n17818 ));
    InMux I__4351 (
            .O(N__25742),
            .I(N__25739));
    LocalMux I__4350 (
            .O(N__25739),
            .I(N__25736));
    Span4Mux_h I__4349 (
            .O(N__25736),
            .I(N__25733));
    Odrv4 I__4348 (
            .O(N__25733),
            .I(\c0.n6_adj_2432 ));
    CascadeMux I__4347 (
            .O(N__25730),
            .I(\c0.n18372_cascade_ ));
    InMux I__4346 (
            .O(N__25727),
            .I(N__25724));
    LocalMux I__4345 (
            .O(N__25724),
            .I(N__25720));
    CascadeMux I__4344 (
            .O(N__25723),
            .I(N__25717));
    Span4Mux_h I__4343 (
            .O(N__25720),
            .I(N__25714));
    InMux I__4342 (
            .O(N__25717),
            .I(N__25711));
    Span4Mux_v I__4341 (
            .O(N__25714),
            .I(N__25705));
    LocalMux I__4340 (
            .O(N__25711),
            .I(N__25705));
    InMux I__4339 (
            .O(N__25710),
            .I(N__25702));
    Span4Mux_v I__4338 (
            .O(N__25705),
            .I(N__25699));
    LocalMux I__4337 (
            .O(N__25702),
            .I(data_in_7_3));
    Odrv4 I__4336 (
            .O(N__25699),
            .I(data_in_7_3));
    InMux I__4335 (
            .O(N__25694),
            .I(N__25691));
    LocalMux I__4334 (
            .O(N__25691),
            .I(n18054));
    InMux I__4333 (
            .O(N__25688),
            .I(N__25684));
    InMux I__4332 (
            .O(N__25687),
            .I(N__25681));
    LocalMux I__4331 (
            .O(N__25684),
            .I(N__25678));
    LocalMux I__4330 (
            .O(N__25681),
            .I(N__25673));
    Span4Mux_v I__4329 (
            .O(N__25678),
            .I(N__25673));
    Odrv4 I__4328 (
            .O(N__25673),
            .I(data_out_frame2_10_4));
    InMux I__4327 (
            .O(N__25670),
            .I(N__25666));
    InMux I__4326 (
            .O(N__25669),
            .I(N__25663));
    LocalMux I__4325 (
            .O(N__25666),
            .I(N__25658));
    LocalMux I__4324 (
            .O(N__25663),
            .I(N__25658));
    Odrv12 I__4323 (
            .O(N__25658),
            .I(data_out_frame2_11_4));
    InMux I__4322 (
            .O(N__25655),
            .I(N__25652));
    LocalMux I__4321 (
            .O(N__25652),
            .I(N__25648));
    InMux I__4320 (
            .O(N__25651),
            .I(N__25645));
    Span12Mux_v I__4319 (
            .O(N__25648),
            .I(N__25642));
    LocalMux I__4318 (
            .O(N__25645),
            .I(data_out_frame2_14_5));
    Odrv12 I__4317 (
            .O(N__25642),
            .I(data_out_frame2_14_5));
    InMux I__4316 (
            .O(N__25637),
            .I(N__25632));
    InMux I__4315 (
            .O(N__25636),
            .I(N__25628));
    InMux I__4314 (
            .O(N__25635),
            .I(N__25625));
    LocalMux I__4313 (
            .O(N__25632),
            .I(N__25622));
    CascadeMux I__4312 (
            .O(N__25631),
            .I(N__25619));
    LocalMux I__4311 (
            .O(N__25628),
            .I(N__25614));
    LocalMux I__4310 (
            .O(N__25625),
            .I(N__25614));
    Span4Mux_v I__4309 (
            .O(N__25622),
            .I(N__25611));
    InMux I__4308 (
            .O(N__25619),
            .I(N__25608));
    Span4Mux_v I__4307 (
            .O(N__25614),
            .I(N__25605));
    Span4Mux_v I__4306 (
            .O(N__25611),
            .I(N__25600));
    LocalMux I__4305 (
            .O(N__25608),
            .I(N__25600));
    Span4Mux_h I__4304 (
            .O(N__25605),
            .I(N__25597));
    Span4Mux_h I__4303 (
            .O(N__25600),
            .I(N__25594));
    Odrv4 I__4302 (
            .O(N__25597),
            .I(\c0.data_in_frame_10_0 ));
    Odrv4 I__4301 (
            .O(N__25594),
            .I(\c0.data_in_frame_10_0 ));
    CascadeMux I__4300 (
            .O(N__25589),
            .I(N__25584));
    InMux I__4299 (
            .O(N__25588),
            .I(N__25579));
    InMux I__4298 (
            .O(N__25587),
            .I(N__25576));
    InMux I__4297 (
            .O(N__25584),
            .I(N__25573));
    InMux I__4296 (
            .O(N__25583),
            .I(N__25570));
    InMux I__4295 (
            .O(N__25582),
            .I(N__25567));
    LocalMux I__4294 (
            .O(N__25579),
            .I(N__25564));
    LocalMux I__4293 (
            .O(N__25576),
            .I(N__25561));
    LocalMux I__4292 (
            .O(N__25573),
            .I(N__25556));
    LocalMux I__4291 (
            .O(N__25570),
            .I(N__25556));
    LocalMux I__4290 (
            .O(N__25567),
            .I(N__25550));
    Span4Mux_h I__4289 (
            .O(N__25564),
            .I(N__25550));
    Span4Mux_v I__4288 (
            .O(N__25561),
            .I(N__25545));
    Span4Mux_v I__4287 (
            .O(N__25556),
            .I(N__25545));
    InMux I__4286 (
            .O(N__25555),
            .I(N__25542));
    Span4Mux_v I__4285 (
            .O(N__25550),
            .I(N__25539));
    Span4Mux_h I__4284 (
            .O(N__25545),
            .I(N__25536));
    LocalMux I__4283 (
            .O(N__25542),
            .I(data_in_frame_8_3));
    Odrv4 I__4282 (
            .O(N__25539),
            .I(data_in_frame_8_3));
    Odrv4 I__4281 (
            .O(N__25536),
            .I(data_in_frame_8_3));
    InMux I__4280 (
            .O(N__25529),
            .I(N__25526));
    LocalMux I__4279 (
            .O(N__25526),
            .I(N__25522));
    InMux I__4278 (
            .O(N__25525),
            .I(N__25519));
    Span4Mux_v I__4277 (
            .O(N__25522),
            .I(N__25516));
    LocalMux I__4276 (
            .O(N__25519),
            .I(N__25513));
    Span4Mux_h I__4275 (
            .O(N__25516),
            .I(N__25510));
    Span4Mux_h I__4274 (
            .O(N__25513),
            .I(N__25507));
    Odrv4 I__4273 (
            .O(N__25510),
            .I(n9380));
    Odrv4 I__4272 (
            .O(N__25507),
            .I(n9380));
    InMux I__4271 (
            .O(N__25502),
            .I(N__25498));
    InMux I__4270 (
            .O(N__25501),
            .I(N__25495));
    LocalMux I__4269 (
            .O(N__25498),
            .I(N__25492));
    LocalMux I__4268 (
            .O(N__25495),
            .I(N__25489));
    Span4Mux_s3_h I__4267 (
            .O(N__25492),
            .I(N__25486));
    Span4Mux_v I__4266 (
            .O(N__25489),
            .I(N__25483));
    Span4Mux_v I__4265 (
            .O(N__25486),
            .I(N__25480));
    Odrv4 I__4264 (
            .O(N__25483),
            .I(n9054));
    Odrv4 I__4263 (
            .O(N__25480),
            .I(n9054));
    CascadeMux I__4262 (
            .O(N__25475),
            .I(n6_adj_2604_cascade_));
    InMux I__4261 (
            .O(N__25472),
            .I(N__25468));
    InMux I__4260 (
            .O(N__25471),
            .I(N__25465));
    LocalMux I__4259 (
            .O(N__25468),
            .I(N__25462));
    LocalMux I__4258 (
            .O(N__25465),
            .I(N__25458));
    Span4Mux_h I__4257 (
            .O(N__25462),
            .I(N__25455));
    InMux I__4256 (
            .O(N__25461),
            .I(N__25452));
    Odrv12 I__4255 (
            .O(N__25458),
            .I(data_in_frame_7_0));
    Odrv4 I__4254 (
            .O(N__25455),
            .I(data_in_frame_7_0));
    LocalMux I__4253 (
            .O(N__25452),
            .I(data_in_frame_7_0));
    InMux I__4252 (
            .O(N__25445),
            .I(N__25440));
    InMux I__4251 (
            .O(N__25444),
            .I(N__25437));
    InMux I__4250 (
            .O(N__25443),
            .I(N__25434));
    LocalMux I__4249 (
            .O(N__25440),
            .I(N__25429));
    LocalMux I__4248 (
            .O(N__25437),
            .I(N__25424));
    LocalMux I__4247 (
            .O(N__25434),
            .I(N__25424));
    InMux I__4246 (
            .O(N__25433),
            .I(N__25421));
    InMux I__4245 (
            .O(N__25432),
            .I(N__25418));
    Span4Mux_v I__4244 (
            .O(N__25429),
            .I(N__25413));
    Span4Mux_v I__4243 (
            .O(N__25424),
            .I(N__25413));
    LocalMux I__4242 (
            .O(N__25421),
            .I(N__25410));
    LocalMux I__4241 (
            .O(N__25418),
            .I(\c0.data_in_frame_1_7 ));
    Odrv4 I__4240 (
            .O(N__25413),
            .I(\c0.data_in_frame_1_7 ));
    Odrv12 I__4239 (
            .O(N__25410),
            .I(\c0.data_in_frame_1_7 ));
    CascadeMux I__4238 (
            .O(N__25403),
            .I(N__25400));
    InMux I__4237 (
            .O(N__25400),
            .I(N__25396));
    CascadeMux I__4236 (
            .O(N__25399),
            .I(N__25393));
    LocalMux I__4235 (
            .O(N__25396),
            .I(N__25390));
    InMux I__4234 (
            .O(N__25393),
            .I(N__25386));
    Span4Mux_v I__4233 (
            .O(N__25390),
            .I(N__25382));
    InMux I__4232 (
            .O(N__25389),
            .I(N__25379));
    LocalMux I__4231 (
            .O(N__25386),
            .I(N__25376));
    InMux I__4230 (
            .O(N__25385),
            .I(N__25373));
    Span4Mux_h I__4229 (
            .O(N__25382),
            .I(N__25366));
    LocalMux I__4228 (
            .O(N__25379),
            .I(N__25366));
    Span4Mux_v I__4227 (
            .O(N__25376),
            .I(N__25366));
    LocalMux I__4226 (
            .O(N__25373),
            .I(\c0.data_in_frame_3_5 ));
    Odrv4 I__4225 (
            .O(N__25366),
            .I(\c0.data_in_frame_3_5 ));
    InMux I__4224 (
            .O(N__25361),
            .I(N__25358));
    LocalMux I__4223 (
            .O(N__25358),
            .I(N__25355));
    Span4Mux_v I__4222 (
            .O(N__25355),
            .I(N__25352));
    Span4Mux_h I__4221 (
            .O(N__25352),
            .I(N__25349));
    Odrv4 I__4220 (
            .O(N__25349),
            .I(\c0.n17614 ));
    InMux I__4219 (
            .O(N__25346),
            .I(N__25342));
    InMux I__4218 (
            .O(N__25345),
            .I(N__25339));
    LocalMux I__4217 (
            .O(N__25342),
            .I(N__25336));
    LocalMux I__4216 (
            .O(N__25339),
            .I(N__25333));
    Span4Mux_v I__4215 (
            .O(N__25336),
            .I(N__25326));
    Span4Mux_h I__4214 (
            .O(N__25333),
            .I(N__25326));
    InMux I__4213 (
            .O(N__25332),
            .I(N__25321));
    InMux I__4212 (
            .O(N__25331),
            .I(N__25321));
    Odrv4 I__4211 (
            .O(N__25326),
            .I(\c0.n8666 ));
    LocalMux I__4210 (
            .O(N__25321),
            .I(\c0.n8666 ));
    InMux I__4209 (
            .O(N__25316),
            .I(N__25313));
    LocalMux I__4208 (
            .O(N__25313),
            .I(N__25310));
    Span4Mux_s1_h I__4207 (
            .O(N__25310),
            .I(N__25306));
    InMux I__4206 (
            .O(N__25309),
            .I(N__25303));
    Span4Mux_h I__4205 (
            .O(N__25306),
            .I(N__25300));
    LocalMux I__4204 (
            .O(N__25303),
            .I(data_out_frame2_14_1));
    Odrv4 I__4203 (
            .O(N__25300),
            .I(data_out_frame2_14_1));
    InMux I__4202 (
            .O(N__25295),
            .I(N__25292));
    LocalMux I__4201 (
            .O(N__25292),
            .I(n18104));
    InMux I__4200 (
            .O(N__25289),
            .I(N__25286));
    LocalMux I__4199 (
            .O(N__25286),
            .I(n18097));
    InMux I__4198 (
            .O(N__25283),
            .I(N__25280));
    LocalMux I__4197 (
            .O(N__25280),
            .I(n18103));
    InMux I__4196 (
            .O(N__25277),
            .I(N__25274));
    LocalMux I__4195 (
            .O(N__25274),
            .I(N__25267));
    InMux I__4194 (
            .O(N__25273),
            .I(N__25264));
    CascadeMux I__4193 (
            .O(N__25272),
            .I(N__25260));
    CascadeMux I__4192 (
            .O(N__25271),
            .I(N__25257));
    InMux I__4191 (
            .O(N__25270),
            .I(N__25254));
    Span4Mux_h I__4190 (
            .O(N__25267),
            .I(N__25251));
    LocalMux I__4189 (
            .O(N__25264),
            .I(N__25248));
    InMux I__4188 (
            .O(N__25263),
            .I(N__25241));
    InMux I__4187 (
            .O(N__25260),
            .I(N__25241));
    InMux I__4186 (
            .O(N__25257),
            .I(N__25241));
    LocalMux I__4185 (
            .O(N__25254),
            .I(data_in_frame_5_4));
    Odrv4 I__4184 (
            .O(N__25251),
            .I(data_in_frame_5_4));
    Odrv12 I__4183 (
            .O(N__25248),
            .I(data_in_frame_5_4));
    LocalMux I__4182 (
            .O(N__25241),
            .I(data_in_frame_5_4));
    InMux I__4181 (
            .O(N__25232),
            .I(N__25229));
    LocalMux I__4180 (
            .O(N__25229),
            .I(N__25226));
    Span4Mux_h I__4179 (
            .O(N__25226),
            .I(N__25223));
    Odrv4 I__4178 (
            .O(N__25223),
            .I(\c0.n2603 ));
    InMux I__4177 (
            .O(N__25220),
            .I(N__25217));
    LocalMux I__4176 (
            .O(N__25217),
            .I(N__25214));
    Span4Mux_h I__4175 (
            .O(N__25214),
            .I(N__25211));
    Odrv4 I__4174 (
            .O(N__25211),
            .I(n2568));
    InMux I__4173 (
            .O(N__25208),
            .I(N__25204));
    InMux I__4172 (
            .O(N__25207),
            .I(N__25201));
    LocalMux I__4171 (
            .O(N__25204),
            .I(N__25198));
    LocalMux I__4170 (
            .O(N__25201),
            .I(\c0.n17538 ));
    Odrv12 I__4169 (
            .O(N__25198),
            .I(\c0.n17538 ));
    InMux I__4168 (
            .O(N__25193),
            .I(N__25190));
    LocalMux I__4167 (
            .O(N__25190),
            .I(N__25186));
    InMux I__4166 (
            .O(N__25189),
            .I(N__25183));
    Odrv4 I__4165 (
            .O(N__25186),
            .I(\c0.n9355 ));
    LocalMux I__4164 (
            .O(N__25183),
            .I(\c0.n9355 ));
    CascadeMux I__4163 (
            .O(N__25178),
            .I(n2568_cascade_));
    InMux I__4162 (
            .O(N__25175),
            .I(N__25171));
    InMux I__4161 (
            .O(N__25174),
            .I(N__25168));
    LocalMux I__4160 (
            .O(N__25171),
            .I(N__25165));
    LocalMux I__4159 (
            .O(N__25168),
            .I(N__25162));
    Span4Mux_h I__4158 (
            .O(N__25165),
            .I(N__25159));
    Span4Mux_v I__4157 (
            .O(N__25162),
            .I(N__25156));
    Span4Mux_v I__4156 (
            .O(N__25159),
            .I(N__25153));
    Span4Mux_h I__4155 (
            .O(N__25156),
            .I(N__25150));
    Odrv4 I__4154 (
            .O(N__25153),
            .I(\c0.n17541 ));
    Odrv4 I__4153 (
            .O(N__25150),
            .I(\c0.n17541 ));
    CascadeMux I__4152 (
            .O(N__25145),
            .I(\c0.n21_cascade_ ));
    InMux I__4151 (
            .O(N__25142),
            .I(N__25139));
    LocalMux I__4150 (
            .O(N__25139),
            .I(\c0.n25 ));
    CascadeMux I__4149 (
            .O(N__25136),
            .I(\c0.n27_cascade_ ));
    InMux I__4148 (
            .O(N__25133),
            .I(N__25129));
    InMux I__4147 (
            .O(N__25132),
            .I(N__25126));
    LocalMux I__4146 (
            .O(N__25129),
            .I(N__25123));
    LocalMux I__4145 (
            .O(N__25126),
            .I(N__25120));
    Span4Mux_h I__4144 (
            .O(N__25123),
            .I(N__25117));
    Odrv4 I__4143 (
            .O(N__25120),
            .I(\c0.n5_adj_2438 ));
    Odrv4 I__4142 (
            .O(N__25117),
            .I(\c0.n5_adj_2438 ));
    InMux I__4141 (
            .O(N__25112),
            .I(N__25109));
    LocalMux I__4140 (
            .O(N__25109),
            .I(N__25103));
    InMux I__4139 (
            .O(N__25108),
            .I(N__25100));
    CascadeMux I__4138 (
            .O(N__25107),
            .I(N__25097));
    InMux I__4137 (
            .O(N__25106),
            .I(N__25094));
    Span4Mux_v I__4136 (
            .O(N__25103),
            .I(N__25089));
    LocalMux I__4135 (
            .O(N__25100),
            .I(N__25089));
    InMux I__4134 (
            .O(N__25097),
            .I(N__25086));
    LocalMux I__4133 (
            .O(N__25094),
            .I(N__25083));
    Span4Mux_v I__4132 (
            .O(N__25089),
            .I(N__25080));
    LocalMux I__4131 (
            .O(N__25086),
            .I(\c0.data_in_frame_6_7 ));
    Odrv4 I__4130 (
            .O(N__25083),
            .I(\c0.data_in_frame_6_7 ));
    Odrv4 I__4129 (
            .O(N__25080),
            .I(\c0.data_in_frame_6_7 ));
    InMux I__4128 (
            .O(N__25073),
            .I(N__25070));
    LocalMux I__4127 (
            .O(N__25070),
            .I(N__25067));
    Odrv12 I__4126 (
            .O(N__25067),
            .I(\c0.n4_adj_2548 ));
    InMux I__4125 (
            .O(N__25064),
            .I(N__25059));
    InMux I__4124 (
            .O(N__25063),
            .I(N__25056));
    InMux I__4123 (
            .O(N__25062),
            .I(N__25053));
    LocalMux I__4122 (
            .O(N__25059),
            .I(N__25049));
    LocalMux I__4121 (
            .O(N__25056),
            .I(N__25046));
    LocalMux I__4120 (
            .O(N__25053),
            .I(N__25043));
    InMux I__4119 (
            .O(N__25052),
            .I(N__25040));
    Span4Mux_v I__4118 (
            .O(N__25049),
            .I(N__25037));
    Span4Mux_h I__4117 (
            .O(N__25046),
            .I(N__25032));
    Span4Mux_s3_h I__4116 (
            .O(N__25043),
            .I(N__25032));
    LocalMux I__4115 (
            .O(N__25040),
            .I(data_in_frame_8_4));
    Odrv4 I__4114 (
            .O(N__25037),
            .I(data_in_frame_8_4));
    Odrv4 I__4113 (
            .O(N__25032),
            .I(data_in_frame_8_4));
    InMux I__4112 (
            .O(N__25025),
            .I(N__25022));
    LocalMux I__4111 (
            .O(N__25022),
            .I(N__25018));
    InMux I__4110 (
            .O(N__25021),
            .I(N__25015));
    Span4Mux_v I__4109 (
            .O(N__25018),
            .I(N__25012));
    LocalMux I__4108 (
            .O(N__25015),
            .I(N__25009));
    Span4Mux_h I__4107 (
            .O(N__25012),
            .I(N__25006));
    Span4Mux_h I__4106 (
            .O(N__25009),
            .I(N__25003));
    Span4Mux_h I__4105 (
            .O(N__25006),
            .I(N__25000));
    Odrv4 I__4104 (
            .O(N__25003),
            .I(n19_adj_2651));
    Odrv4 I__4103 (
            .O(N__25000),
            .I(n19_adj_2651));
    InMux I__4102 (
            .O(N__24995),
            .I(N__24991));
    InMux I__4101 (
            .O(N__24994),
            .I(N__24988));
    LocalMux I__4100 (
            .O(N__24991),
            .I(N__24985));
    LocalMux I__4099 (
            .O(N__24988),
            .I(N__24982));
    Span4Mux_v I__4098 (
            .O(N__24985),
            .I(N__24979));
    Span4Mux_h I__4097 (
            .O(N__24982),
            .I(N__24976));
    Odrv4 I__4096 (
            .O(N__24979),
            .I(\c0.n8658 ));
    Odrv4 I__4095 (
            .O(N__24976),
            .I(\c0.n8658 ));
    InMux I__4094 (
            .O(N__24971),
            .I(N__24967));
    InMux I__4093 (
            .O(N__24970),
            .I(N__24964));
    LocalMux I__4092 (
            .O(N__24967),
            .I(N__24960));
    LocalMux I__4091 (
            .O(N__24964),
            .I(N__24957));
    InMux I__4090 (
            .O(N__24963),
            .I(N__24952));
    Span4Mux_h I__4089 (
            .O(N__24960),
            .I(N__24947));
    Span4Mux_h I__4088 (
            .O(N__24957),
            .I(N__24947));
    InMux I__4087 (
            .O(N__24956),
            .I(N__24942));
    InMux I__4086 (
            .O(N__24955),
            .I(N__24942));
    LocalMux I__4085 (
            .O(N__24952),
            .I(data_in_frame_5_1));
    Odrv4 I__4084 (
            .O(N__24947),
            .I(data_in_frame_5_1));
    LocalMux I__4083 (
            .O(N__24942),
            .I(data_in_frame_5_1));
    InMux I__4082 (
            .O(N__24935),
            .I(N__24932));
    LocalMux I__4081 (
            .O(N__24932),
            .I(N__24928));
    InMux I__4080 (
            .O(N__24931),
            .I(N__24925));
    Span4Mux_h I__4079 (
            .O(N__24928),
            .I(N__24922));
    LocalMux I__4078 (
            .O(N__24925),
            .I(N__24919));
    Span4Mux_h I__4077 (
            .O(N__24922),
            .I(N__24916));
    Odrv4 I__4076 (
            .O(N__24919),
            .I(\c0.n17516 ));
    Odrv4 I__4075 (
            .O(N__24916),
            .I(\c0.n17516 ));
    CascadeMux I__4074 (
            .O(N__24911),
            .I(\c0.n2601_cascade_ ));
    InMux I__4073 (
            .O(N__24908),
            .I(N__24905));
    LocalMux I__4072 (
            .O(N__24905),
            .I(N__24902));
    Span4Mux_v I__4071 (
            .O(N__24902),
            .I(N__24897));
    InMux I__4070 (
            .O(N__24901),
            .I(N__24894));
    InMux I__4069 (
            .O(N__24900),
            .I(N__24891));
    Odrv4 I__4068 (
            .O(N__24897),
            .I(n2597));
    LocalMux I__4067 (
            .O(N__24894),
            .I(n2597));
    LocalMux I__4066 (
            .O(N__24891),
            .I(n2597));
    InMux I__4065 (
            .O(N__24884),
            .I(N__24880));
    InMux I__4064 (
            .O(N__24883),
            .I(N__24876));
    LocalMux I__4063 (
            .O(N__24880),
            .I(N__24873));
    InMux I__4062 (
            .O(N__24879),
            .I(N__24870));
    LocalMux I__4061 (
            .O(N__24876),
            .I(N__24867));
    Span4Mux_s3_h I__4060 (
            .O(N__24873),
            .I(N__24864));
    LocalMux I__4059 (
            .O(N__24870),
            .I(N__24861));
    Span4Mux_h I__4058 (
            .O(N__24867),
            .I(N__24856));
    Span4Mux_v I__4057 (
            .O(N__24864),
            .I(N__24856));
    Span4Mux_h I__4056 (
            .O(N__24861),
            .I(N__24853));
    Odrv4 I__4055 (
            .O(N__24856),
            .I(\c0.n9039 ));
    Odrv4 I__4054 (
            .O(N__24853),
            .I(\c0.n9039 ));
    InMux I__4053 (
            .O(N__24848),
            .I(N__24845));
    LocalMux I__4052 (
            .O(N__24845),
            .I(N__24842));
    Span4Mux_v I__4051 (
            .O(N__24842),
            .I(N__24839));
    Span4Mux_h I__4050 (
            .O(N__24839),
            .I(N__24835));
    InMux I__4049 (
            .O(N__24838),
            .I(N__24832));
    Span4Mux_s2_h I__4048 (
            .O(N__24835),
            .I(N__24829));
    LocalMux I__4047 (
            .O(N__24832),
            .I(N__24826));
    Odrv4 I__4046 (
            .O(N__24829),
            .I(\c0.n17522 ));
    Odrv12 I__4045 (
            .O(N__24826),
            .I(\c0.n17522 ));
    InMux I__4044 (
            .O(N__24821),
            .I(N__24818));
    LocalMux I__4043 (
            .O(N__24818),
            .I(\c0.n2606 ));
    CascadeMux I__4042 (
            .O(N__24815),
            .I(\c0.n17428_cascade_ ));
    InMux I__4041 (
            .O(N__24812),
            .I(N__24809));
    LocalMux I__4040 (
            .O(N__24809),
            .I(\c0.n11_adj_2494 ));
    InMux I__4039 (
            .O(N__24806),
            .I(N__24803));
    LocalMux I__4038 (
            .O(N__24803),
            .I(N__24800));
    Span4Mux_v I__4037 (
            .O(N__24800),
            .I(N__24797));
    Span4Mux_s2_h I__4036 (
            .O(N__24797),
            .I(N__24794));
    Odrv4 I__4035 (
            .O(N__24794),
            .I(\c0.n14 ));
    InMux I__4034 (
            .O(N__24791),
            .I(N__24785));
    InMux I__4033 (
            .O(N__24790),
            .I(N__24785));
    LocalMux I__4032 (
            .O(N__24785),
            .I(\c0.n17575 ));
    InMux I__4031 (
            .O(N__24782),
            .I(N__24778));
    InMux I__4030 (
            .O(N__24781),
            .I(N__24775));
    LocalMux I__4029 (
            .O(N__24778),
            .I(N__24772));
    LocalMux I__4028 (
            .O(N__24775),
            .I(N__24769));
    Odrv4 I__4027 (
            .O(N__24772),
            .I(\c0.n9103 ));
    Odrv4 I__4026 (
            .O(N__24769),
            .I(\c0.n9103 ));
    CascadeMux I__4025 (
            .O(N__24764),
            .I(N__24760));
    InMux I__4024 (
            .O(N__24763),
            .I(N__24755));
    InMux I__4023 (
            .O(N__24760),
            .I(N__24750));
    InMux I__4022 (
            .O(N__24759),
            .I(N__24747));
    InMux I__4021 (
            .O(N__24758),
            .I(N__24744));
    LocalMux I__4020 (
            .O(N__24755),
            .I(N__24741));
    InMux I__4019 (
            .O(N__24754),
            .I(N__24736));
    InMux I__4018 (
            .O(N__24753),
            .I(N__24736));
    LocalMux I__4017 (
            .O(N__24750),
            .I(N__24733));
    LocalMux I__4016 (
            .O(N__24747),
            .I(N__24730));
    LocalMux I__4015 (
            .O(N__24744),
            .I(N__24725));
    Span4Mux_v I__4014 (
            .O(N__24741),
            .I(N__24725));
    LocalMux I__4013 (
            .O(N__24736),
            .I(N__24722));
    Span4Mux_v I__4012 (
            .O(N__24733),
            .I(N__24715));
    Span4Mux_v I__4011 (
            .O(N__24730),
            .I(N__24715));
    Sp12to4 I__4010 (
            .O(N__24725),
            .I(N__24710));
    Span12Mux_s11_v I__4009 (
            .O(N__24722),
            .I(N__24710));
    InMux I__4008 (
            .O(N__24721),
            .I(N__24705));
    InMux I__4007 (
            .O(N__24720),
            .I(N__24705));
    Odrv4 I__4006 (
            .O(N__24715),
            .I(data_in_frame_5_2));
    Odrv12 I__4005 (
            .O(N__24710),
            .I(data_in_frame_5_2));
    LocalMux I__4004 (
            .O(N__24705),
            .I(data_in_frame_5_2));
    CascadeMux I__4003 (
            .O(N__24698),
            .I(N__24695));
    InMux I__4002 (
            .O(N__24695),
            .I(N__24688));
    InMux I__4001 (
            .O(N__24694),
            .I(N__24683));
    InMux I__4000 (
            .O(N__24693),
            .I(N__24683));
    CascadeMux I__3999 (
            .O(N__24692),
            .I(N__24679));
    CascadeMux I__3998 (
            .O(N__24691),
            .I(N__24674));
    LocalMux I__3997 (
            .O(N__24688),
            .I(N__24670));
    LocalMux I__3996 (
            .O(N__24683),
            .I(N__24667));
    InMux I__3995 (
            .O(N__24682),
            .I(N__24660));
    InMux I__3994 (
            .O(N__24679),
            .I(N__24660));
    InMux I__3993 (
            .O(N__24678),
            .I(N__24660));
    CascadeMux I__3992 (
            .O(N__24677),
            .I(N__24657));
    InMux I__3991 (
            .O(N__24674),
            .I(N__24654));
    InMux I__3990 (
            .O(N__24673),
            .I(N__24651));
    Span4Mux_v I__3989 (
            .O(N__24670),
            .I(N__24648));
    Span4Mux_h I__3988 (
            .O(N__24667),
            .I(N__24643));
    LocalMux I__3987 (
            .O(N__24660),
            .I(N__24643));
    InMux I__3986 (
            .O(N__24657),
            .I(N__24640));
    LocalMux I__3985 (
            .O(N__24654),
            .I(N__24637));
    LocalMux I__3984 (
            .O(N__24651),
            .I(N__24634));
    Sp12to4 I__3983 (
            .O(N__24648),
            .I(N__24631));
    Span4Mux_v I__3982 (
            .O(N__24643),
            .I(N__24628));
    LocalMux I__3981 (
            .O(N__24640),
            .I(N__24621));
    Span4Mux_h I__3980 (
            .O(N__24637),
            .I(N__24621));
    Span4Mux_s2_h I__3979 (
            .O(N__24634),
            .I(N__24621));
    Odrv12 I__3978 (
            .O(N__24631),
            .I(data_in_frame_5_6));
    Odrv4 I__3977 (
            .O(N__24628),
            .I(data_in_frame_5_6));
    Odrv4 I__3976 (
            .O(N__24621),
            .I(data_in_frame_5_6));
    CascadeMux I__3975 (
            .O(N__24614),
            .I(N__24611));
    InMux I__3974 (
            .O(N__24611),
            .I(N__24608));
    LocalMux I__3973 (
            .O(N__24608),
            .I(\c0.n17430 ));
    CascadeMux I__3972 (
            .O(N__24605),
            .I(N__24602));
    InMux I__3971 (
            .O(N__24602),
            .I(N__24599));
    LocalMux I__3970 (
            .O(N__24599),
            .I(N__24595));
    InMux I__3969 (
            .O(N__24598),
            .I(N__24591));
    Span12Mux_s4_h I__3968 (
            .O(N__24595),
            .I(N__24588));
    InMux I__3967 (
            .O(N__24594),
            .I(N__24585));
    LocalMux I__3966 (
            .O(N__24591),
            .I(data_in_7_0));
    Odrv12 I__3965 (
            .O(N__24588),
            .I(data_in_7_0));
    LocalMux I__3964 (
            .O(N__24585),
            .I(data_in_7_0));
    CascadeMux I__3963 (
            .O(N__24578),
            .I(\c0.n4_adj_2512_cascade_ ));
    InMux I__3962 (
            .O(N__24575),
            .I(N__24572));
    LocalMux I__3961 (
            .O(N__24572),
            .I(N__24569));
    Span4Mux_s3_h I__3960 (
            .O(N__24569),
            .I(N__24566));
    Span4Mux_v I__3959 (
            .O(N__24566),
            .I(N__24563));
    Odrv4 I__3958 (
            .O(N__24563),
            .I(n2591));
    InMux I__3957 (
            .O(N__24560),
            .I(N__24557));
    LocalMux I__3956 (
            .O(N__24557),
            .I(N__24552));
    InMux I__3955 (
            .O(N__24556),
            .I(N__24549));
    InMux I__3954 (
            .O(N__24555),
            .I(N__24546));
    Span4Mux_h I__3953 (
            .O(N__24552),
            .I(N__24543));
    LocalMux I__3952 (
            .O(N__24549),
            .I(N__24540));
    LocalMux I__3951 (
            .O(N__24546),
            .I(N__24537));
    Span4Mux_v I__3950 (
            .O(N__24543),
            .I(N__24532));
    Span4Mux_s3_h I__3949 (
            .O(N__24540),
            .I(N__24532));
    Span4Mux_h I__3948 (
            .O(N__24537),
            .I(N__24529));
    Odrv4 I__3947 (
            .O(N__24532),
            .I(\c0.n8751 ));
    Odrv4 I__3946 (
            .O(N__24529),
            .I(\c0.n8751 ));
    InMux I__3945 (
            .O(N__24524),
            .I(N__24520));
    InMux I__3944 (
            .O(N__24523),
            .I(N__24517));
    LocalMux I__3943 (
            .O(N__24520),
            .I(N__24514));
    LocalMux I__3942 (
            .O(N__24517),
            .I(N__24509));
    Span4Mux_h I__3941 (
            .O(N__24514),
            .I(N__24509));
    Odrv4 I__3940 (
            .O(N__24509),
            .I(\c0.n17532 ));
    CascadeMux I__3939 (
            .O(N__24506),
            .I(n2591_cascade_));
    InMux I__3938 (
            .O(N__24503),
            .I(N__24500));
    LocalMux I__3937 (
            .O(N__24500),
            .I(N__24496));
    InMux I__3936 (
            .O(N__24499),
            .I(N__24493));
    Span4Mux_h I__3935 (
            .O(N__24496),
            .I(N__24490));
    LocalMux I__3934 (
            .O(N__24493),
            .I(N__24487));
    Odrv4 I__3933 (
            .O(N__24490),
            .I(\c0.n9324 ));
    Odrv12 I__3932 (
            .O(N__24487),
            .I(\c0.n9324 ));
    InMux I__3931 (
            .O(N__24482),
            .I(N__24479));
    LocalMux I__3930 (
            .O(N__24479),
            .I(\c0.n17533 ));
    InMux I__3929 (
            .O(N__24476),
            .I(N__24473));
    LocalMux I__3928 (
            .O(N__24473),
            .I(\c0.n2605 ));
    InMux I__3927 (
            .O(N__24470),
            .I(N__24467));
    LocalMux I__3926 (
            .O(N__24467),
            .I(N__24464));
    Span4Mux_v I__3925 (
            .O(N__24464),
            .I(N__24461));
    Odrv4 I__3924 (
            .O(N__24461),
            .I(n2570));
    CascadeMux I__3923 (
            .O(N__24458),
            .I(n2570_cascade_));
    InMux I__3922 (
            .O(N__24455),
            .I(N__24452));
    LocalMux I__3921 (
            .O(N__24452),
            .I(N__24449));
    Odrv4 I__3920 (
            .O(N__24449),
            .I(\c0.n8556 ));
    CascadeMux I__3919 (
            .O(N__24446),
            .I(\c0.n17_adj_2514_cascade_ ));
    InMux I__3918 (
            .O(N__24443),
            .I(N__24440));
    LocalMux I__3917 (
            .O(N__24440),
            .I(N__24435));
    InMux I__3916 (
            .O(N__24439),
            .I(N__24430));
    InMux I__3915 (
            .O(N__24438),
            .I(N__24430));
    Span4Mux_h I__3914 (
            .O(N__24435),
            .I(N__24427));
    LocalMux I__3913 (
            .O(N__24430),
            .I(N__24424));
    Odrv4 I__3912 (
            .O(N__24427),
            .I(\c0.data_in_frame_6_2 ));
    Odrv12 I__3911 (
            .O(N__24424),
            .I(\c0.data_in_frame_6_2 ));
    CascadeMux I__3910 (
            .O(N__24419),
            .I(FRAME_MATCHER_next_state_31_N_2026_1_cascade_));
    InMux I__3909 (
            .O(N__24416),
            .I(N__24412));
    InMux I__3908 (
            .O(N__24415),
            .I(N__24409));
    LocalMux I__3907 (
            .O(N__24412),
            .I(N__24406));
    LocalMux I__3906 (
            .O(N__24409),
            .I(N__24403));
    Span4Mux_h I__3905 (
            .O(N__24406),
            .I(N__24400));
    Odrv12 I__3904 (
            .O(N__24403),
            .I(n2567));
    Odrv4 I__3903 (
            .O(N__24400),
            .I(n2567));
    CascadeMux I__3902 (
            .O(N__24395),
            .I(\c0.n8556_cascade_ ));
    CascadeMux I__3901 (
            .O(N__24392),
            .I(\c0.n7_cascade_ ));
    InMux I__3900 (
            .O(N__24389),
            .I(N__24386));
    LocalMux I__3899 (
            .O(N__24386),
            .I(\c0.n6_adj_2478 ));
    InMux I__3898 (
            .O(N__24383),
            .I(N__24380));
    LocalMux I__3897 (
            .O(N__24380),
            .I(N__24374));
    InMux I__3896 (
            .O(N__24379),
            .I(N__24371));
    InMux I__3895 (
            .O(N__24378),
            .I(N__24367));
    InMux I__3894 (
            .O(N__24377),
            .I(N__24364));
    Span4Mux_v I__3893 (
            .O(N__24374),
            .I(N__24361));
    LocalMux I__3892 (
            .O(N__24371),
            .I(N__24358));
    InMux I__3891 (
            .O(N__24370),
            .I(N__24355));
    LocalMux I__3890 (
            .O(N__24367),
            .I(data_in_2_2));
    LocalMux I__3889 (
            .O(N__24364),
            .I(data_in_2_2));
    Odrv4 I__3888 (
            .O(N__24361),
            .I(data_in_2_2));
    Odrv4 I__3887 (
            .O(N__24358),
            .I(data_in_2_2));
    LocalMux I__3886 (
            .O(N__24355),
            .I(data_in_2_2));
    InMux I__3885 (
            .O(N__24344),
            .I(N__24340));
    InMux I__3884 (
            .O(N__24343),
            .I(N__24337));
    LocalMux I__3883 (
            .O(N__24340),
            .I(\c0.n8460 ));
    LocalMux I__3882 (
            .O(N__24337),
            .I(\c0.n8460 ));
    InMux I__3881 (
            .O(N__24332),
            .I(N__24329));
    LocalMux I__3880 (
            .O(N__24329),
            .I(N__24326));
    Odrv12 I__3879 (
            .O(N__24326),
            .I(\c0.n17745 ));
    CascadeMux I__3878 (
            .O(N__24323),
            .I(\c0.n16_adj_2485_cascade_ ));
    InMux I__3877 (
            .O(N__24320),
            .I(N__24310));
    InMux I__3876 (
            .O(N__24319),
            .I(N__24310));
    InMux I__3875 (
            .O(N__24318),
            .I(N__24307));
    InMux I__3874 (
            .O(N__24317),
            .I(N__24304));
    InMux I__3873 (
            .O(N__24316),
            .I(N__24299));
    InMux I__3872 (
            .O(N__24315),
            .I(N__24299));
    LocalMux I__3871 (
            .O(N__24310),
            .I(N__24294));
    LocalMux I__3870 (
            .O(N__24307),
            .I(N__24294));
    LocalMux I__3869 (
            .O(N__24304),
            .I(N__24291));
    LocalMux I__3868 (
            .O(N__24299),
            .I(N__24284));
    Span4Mux_v I__3867 (
            .O(N__24294),
            .I(N__24284));
    Span4Mux_h I__3866 (
            .O(N__24291),
            .I(N__24284));
    Odrv4 I__3865 (
            .O(N__24284),
            .I(data_in_frame_10_6));
    CascadeMux I__3864 (
            .O(N__24281),
            .I(n63_adj_2642_cascade_));
    CascadeMux I__3863 (
            .O(N__24278),
            .I(N__24247));
    InMux I__3862 (
            .O(N__24277),
            .I(N__24230));
    InMux I__3861 (
            .O(N__24276),
            .I(N__24230));
    InMux I__3860 (
            .O(N__24275),
            .I(N__24230));
    InMux I__3859 (
            .O(N__24274),
            .I(N__24227));
    InMux I__3858 (
            .O(N__24273),
            .I(N__24222));
    InMux I__3857 (
            .O(N__24272),
            .I(N__24222));
    InMux I__3856 (
            .O(N__24271),
            .I(N__24219));
    InMux I__3855 (
            .O(N__24270),
            .I(N__24205));
    InMux I__3854 (
            .O(N__24269),
            .I(N__24205));
    InMux I__3853 (
            .O(N__24268),
            .I(N__24205));
    InMux I__3852 (
            .O(N__24267),
            .I(N__24202));
    InMux I__3851 (
            .O(N__24266),
            .I(N__24193));
    InMux I__3850 (
            .O(N__24265),
            .I(N__24193));
    InMux I__3849 (
            .O(N__24264),
            .I(N__24193));
    InMux I__3848 (
            .O(N__24263),
            .I(N__24193));
    InMux I__3847 (
            .O(N__24262),
            .I(N__24184));
    InMux I__3846 (
            .O(N__24261),
            .I(N__24184));
    InMux I__3845 (
            .O(N__24260),
            .I(N__24184));
    InMux I__3844 (
            .O(N__24259),
            .I(N__24184));
    InMux I__3843 (
            .O(N__24258),
            .I(N__24181));
    InMux I__3842 (
            .O(N__24257),
            .I(N__24176));
    InMux I__3841 (
            .O(N__24256),
            .I(N__24176));
    InMux I__3840 (
            .O(N__24255),
            .I(N__24171));
    InMux I__3839 (
            .O(N__24254),
            .I(N__24171));
    InMux I__3838 (
            .O(N__24253),
            .I(N__24162));
    InMux I__3837 (
            .O(N__24252),
            .I(N__24162));
    InMux I__3836 (
            .O(N__24251),
            .I(N__24162));
    InMux I__3835 (
            .O(N__24250),
            .I(N__24162));
    InMux I__3834 (
            .O(N__24247),
            .I(N__24159));
    InMux I__3833 (
            .O(N__24246),
            .I(N__24152));
    InMux I__3832 (
            .O(N__24245),
            .I(N__24152));
    InMux I__3831 (
            .O(N__24244),
            .I(N__24152));
    InMux I__3830 (
            .O(N__24243),
            .I(N__24143));
    InMux I__3829 (
            .O(N__24242),
            .I(N__24143));
    InMux I__3828 (
            .O(N__24241),
            .I(N__24143));
    InMux I__3827 (
            .O(N__24240),
            .I(N__24143));
    InMux I__3826 (
            .O(N__24239),
            .I(N__24136));
    InMux I__3825 (
            .O(N__24238),
            .I(N__24136));
    InMux I__3824 (
            .O(N__24237),
            .I(N__24136));
    LocalMux I__3823 (
            .O(N__24230),
            .I(N__24131));
    LocalMux I__3822 (
            .O(N__24227),
            .I(N__24131));
    LocalMux I__3821 (
            .O(N__24222),
            .I(N__24126));
    LocalMux I__3820 (
            .O(N__24219),
            .I(N__24126));
    InMux I__3819 (
            .O(N__24218),
            .I(N__24122));
    InMux I__3818 (
            .O(N__24217),
            .I(N__24119));
    InMux I__3817 (
            .O(N__24216),
            .I(N__24115));
    InMux I__3816 (
            .O(N__24215),
            .I(N__24106));
    InMux I__3815 (
            .O(N__24214),
            .I(N__24106));
    InMux I__3814 (
            .O(N__24213),
            .I(N__24106));
    InMux I__3813 (
            .O(N__24212),
            .I(N__24106));
    LocalMux I__3812 (
            .O(N__24205),
            .I(N__24103));
    LocalMux I__3811 (
            .O(N__24202),
            .I(N__24096));
    LocalMux I__3810 (
            .O(N__24193),
            .I(N__24096));
    LocalMux I__3809 (
            .O(N__24184),
            .I(N__24096));
    LocalMux I__3808 (
            .O(N__24181),
            .I(N__24091));
    LocalMux I__3807 (
            .O(N__24176),
            .I(N__24091));
    LocalMux I__3806 (
            .O(N__24171),
            .I(N__24086));
    LocalMux I__3805 (
            .O(N__24162),
            .I(N__24086));
    LocalMux I__3804 (
            .O(N__24159),
            .I(N__24073));
    LocalMux I__3803 (
            .O(N__24152),
            .I(N__24073));
    LocalMux I__3802 (
            .O(N__24143),
            .I(N__24073));
    LocalMux I__3801 (
            .O(N__24136),
            .I(N__24073));
    Span4Mux_v I__3800 (
            .O(N__24131),
            .I(N__24073));
    Span4Mux_v I__3799 (
            .O(N__24126),
            .I(N__24073));
    InMux I__3798 (
            .O(N__24125),
            .I(N__24066));
    LocalMux I__3797 (
            .O(N__24122),
            .I(N__24061));
    LocalMux I__3796 (
            .O(N__24119),
            .I(N__24061));
    InMux I__3795 (
            .O(N__24118),
            .I(N__24058));
    LocalMux I__3794 (
            .O(N__24115),
            .I(N__24049));
    LocalMux I__3793 (
            .O(N__24106),
            .I(N__24049));
    Span4Mux_v I__3792 (
            .O(N__24103),
            .I(N__24049));
    Span4Mux_v I__3791 (
            .O(N__24096),
            .I(N__24049));
    Span4Mux_v I__3790 (
            .O(N__24091),
            .I(N__24044));
    Span4Mux_v I__3789 (
            .O(N__24086),
            .I(N__24044));
    Span4Mux_h I__3788 (
            .O(N__24073),
            .I(N__24041));
    InMux I__3787 (
            .O(N__24072),
            .I(N__24032));
    InMux I__3786 (
            .O(N__24071),
            .I(N__24032));
    InMux I__3785 (
            .O(N__24070),
            .I(N__24032));
    InMux I__3784 (
            .O(N__24069),
            .I(N__24032));
    LocalMux I__3783 (
            .O(N__24066),
            .I(N__24025));
    Span4Mux_h I__3782 (
            .O(N__24061),
            .I(N__24025));
    LocalMux I__3781 (
            .O(N__24058),
            .I(N__24025));
    Odrv4 I__3780 (
            .O(N__24049),
            .I(n16468));
    Odrv4 I__3779 (
            .O(N__24044),
            .I(n16468));
    Odrv4 I__3778 (
            .O(N__24041),
            .I(n16468));
    LocalMux I__3777 (
            .O(N__24032),
            .I(n16468));
    Odrv4 I__3776 (
            .O(N__24025),
            .I(n16468));
    InMux I__3775 (
            .O(N__24014),
            .I(N__24011));
    LocalMux I__3774 (
            .O(N__24011),
            .I(N__24008));
    Span4Mux_h I__3773 (
            .O(N__24008),
            .I(N__24004));
    InMux I__3772 (
            .O(N__24007),
            .I(N__23999));
    Span4Mux_v I__3771 (
            .O(N__24004),
            .I(N__23996));
    InMux I__3770 (
            .O(N__24003),
            .I(N__23991));
    InMux I__3769 (
            .O(N__24002),
            .I(N__23991));
    LocalMux I__3768 (
            .O(N__23999),
            .I(\c0.data_in_1_0 ));
    Odrv4 I__3767 (
            .O(N__23996),
            .I(\c0.data_in_1_0 ));
    LocalMux I__3766 (
            .O(N__23991),
            .I(\c0.data_in_1_0 ));
    InMux I__3765 (
            .O(N__23984),
            .I(N__23981));
    LocalMux I__3764 (
            .O(N__23981),
            .I(N__23978));
    Span4Mux_h I__3763 (
            .O(N__23978),
            .I(N__23974));
    CascadeMux I__3762 (
            .O(N__23977),
            .I(N__23970));
    Span4Mux_h I__3761 (
            .O(N__23974),
            .I(N__23966));
    InMux I__3760 (
            .O(N__23973),
            .I(N__23959));
    InMux I__3759 (
            .O(N__23970),
            .I(N__23959));
    InMux I__3758 (
            .O(N__23969),
            .I(N__23959));
    Odrv4 I__3757 (
            .O(N__23966),
            .I(\c0.data_in_0_0 ));
    LocalMux I__3756 (
            .O(N__23959),
            .I(\c0.data_in_0_0 ));
    InMux I__3755 (
            .O(N__23954),
            .I(N__23951));
    LocalMux I__3754 (
            .O(N__23951),
            .I(N__23948));
    Span4Mux_v I__3753 (
            .O(N__23948),
            .I(N__23941));
    InMux I__3752 (
            .O(N__23947),
            .I(N__23938));
    InMux I__3751 (
            .O(N__23946),
            .I(N__23931));
    InMux I__3750 (
            .O(N__23945),
            .I(N__23931));
    InMux I__3749 (
            .O(N__23944),
            .I(N__23931));
    Odrv4 I__3748 (
            .O(N__23941),
            .I(data_in_3_7));
    LocalMux I__3747 (
            .O(N__23938),
            .I(data_in_3_7));
    LocalMux I__3746 (
            .O(N__23931),
            .I(data_in_3_7));
    InMux I__3745 (
            .O(N__23924),
            .I(N__23921));
    LocalMux I__3744 (
            .O(N__23921),
            .I(\c0.n6_adj_2473 ));
    CascadeMux I__3743 (
            .O(N__23918),
            .I(N__23915));
    InMux I__3742 (
            .O(N__23915),
            .I(N__23912));
    LocalMux I__3741 (
            .O(N__23912),
            .I(N__23909));
    Span4Mux_v I__3740 (
            .O(N__23909),
            .I(N__23906));
    Span4Mux_h I__3739 (
            .O(N__23906),
            .I(N__23902));
    InMux I__3738 (
            .O(N__23905),
            .I(N__23899));
    Span4Mux_h I__3737 (
            .O(N__23902),
            .I(N__23894));
    LocalMux I__3736 (
            .O(N__23899),
            .I(N__23894));
    Span4Mux_v I__3735 (
            .O(N__23894),
            .I(N__23890));
    InMux I__3734 (
            .O(N__23893),
            .I(N__23887));
    Odrv4 I__3733 (
            .O(N__23890),
            .I(data_in_8_0));
    LocalMux I__3732 (
            .O(N__23887),
            .I(data_in_8_0));
    InMux I__3731 (
            .O(N__23882),
            .I(N__23878));
    InMux I__3730 (
            .O(N__23881),
            .I(N__23874));
    LocalMux I__3729 (
            .O(N__23878),
            .I(N__23870));
    InMux I__3728 (
            .O(N__23877),
            .I(N__23867));
    LocalMux I__3727 (
            .O(N__23874),
            .I(N__23863));
    InMux I__3726 (
            .O(N__23873),
            .I(N__23860));
    Span4Mux_h I__3725 (
            .O(N__23870),
            .I(N__23856));
    LocalMux I__3724 (
            .O(N__23867),
            .I(N__23853));
    InMux I__3723 (
            .O(N__23866),
            .I(N__23850));
    Span4Mux_v I__3722 (
            .O(N__23863),
            .I(N__23845));
    LocalMux I__3721 (
            .O(N__23860),
            .I(N__23845));
    InMux I__3720 (
            .O(N__23859),
            .I(N__23842));
    Odrv4 I__3719 (
            .O(N__23856),
            .I(\c0.n81 ));
    Odrv12 I__3718 (
            .O(N__23853),
            .I(\c0.n81 ));
    LocalMux I__3717 (
            .O(N__23850),
            .I(\c0.n81 ));
    Odrv4 I__3716 (
            .O(N__23845),
            .I(\c0.n81 ));
    LocalMux I__3715 (
            .O(N__23842),
            .I(\c0.n81 ));
    InMux I__3714 (
            .O(N__23831),
            .I(N__23827));
    InMux I__3713 (
            .O(N__23830),
            .I(N__23824));
    LocalMux I__3712 (
            .O(N__23827),
            .I(N__23820));
    LocalMux I__3711 (
            .O(N__23824),
            .I(N__23817));
    InMux I__3710 (
            .O(N__23823),
            .I(N__23814));
    Span12Mux_h I__3709 (
            .O(N__23820),
            .I(N__23811));
    Odrv12 I__3708 (
            .O(N__23817),
            .I(data_in_6_0));
    LocalMux I__3707 (
            .O(N__23814),
            .I(data_in_6_0));
    Odrv12 I__3706 (
            .O(N__23811),
            .I(data_in_6_0));
    InMux I__3705 (
            .O(N__23804),
            .I(N__23801));
    LocalMux I__3704 (
            .O(N__23801),
            .I(N__23798));
    Span4Mux_v I__3703 (
            .O(N__23798),
            .I(N__23795));
    Span4Mux_h I__3702 (
            .O(N__23795),
            .I(N__23790));
    InMux I__3701 (
            .O(N__23794),
            .I(N__23787));
    InMux I__3700 (
            .O(N__23793),
            .I(N__23784));
    Odrv4 I__3699 (
            .O(N__23790),
            .I(\c0.data_in_frame_6_0 ));
    LocalMux I__3698 (
            .O(N__23787),
            .I(\c0.data_in_frame_6_0 ));
    LocalMux I__3697 (
            .O(N__23784),
            .I(\c0.data_in_frame_6_0 ));
    InMux I__3696 (
            .O(N__23777),
            .I(N__23774));
    LocalMux I__3695 (
            .O(N__23774),
            .I(N__23770));
    InMux I__3694 (
            .O(N__23773),
            .I(N__23767));
    Span4Mux_h I__3693 (
            .O(N__23770),
            .I(N__23764));
    LocalMux I__3692 (
            .O(N__23767),
            .I(N__23761));
    Odrv4 I__3691 (
            .O(N__23764),
            .I(n2599));
    Odrv12 I__3690 (
            .O(N__23761),
            .I(n2599));
    CascadeMux I__3689 (
            .O(N__23756),
            .I(n2599_cascade_));
    InMux I__3688 (
            .O(N__23753),
            .I(N__23750));
    LocalMux I__3687 (
            .O(N__23750),
            .I(N__23747));
    Span4Mux_h I__3686 (
            .O(N__23747),
            .I(N__23744));
    Odrv4 I__3685 (
            .O(N__23744),
            .I(\c0.n20_adj_2452 ));
    InMux I__3684 (
            .O(N__23741),
            .I(N__23738));
    LocalMux I__3683 (
            .O(N__23738),
            .I(N__23733));
    InMux I__3682 (
            .O(N__23737),
            .I(N__23730));
    InMux I__3681 (
            .O(N__23736),
            .I(N__23727));
    Odrv12 I__3680 (
            .O(N__23733),
            .I(data_in_0_2));
    LocalMux I__3679 (
            .O(N__23730),
            .I(data_in_0_2));
    LocalMux I__3678 (
            .O(N__23727),
            .I(data_in_0_2));
    CascadeMux I__3677 (
            .O(N__23720),
            .I(\c0.n12_adj_2472_cascade_ ));
    InMux I__3676 (
            .O(N__23717),
            .I(N__23714));
    LocalMux I__3675 (
            .O(N__23714),
            .I(N__23711));
    Span4Mux_v I__3674 (
            .O(N__23711),
            .I(N__23708));
    Odrv4 I__3673 (
            .O(N__23708),
            .I(\c0.n17765 ));
    InMux I__3672 (
            .O(N__23705),
            .I(n16349));
    CascadeMux I__3671 (
            .O(N__23702),
            .I(N__23699));
    InMux I__3670 (
            .O(N__23699),
            .I(N__23695));
    CascadeMux I__3669 (
            .O(N__23698),
            .I(N__23692));
    LocalMux I__3668 (
            .O(N__23695),
            .I(N__23689));
    InMux I__3667 (
            .O(N__23692),
            .I(N__23686));
    Span4Mux_s2_h I__3666 (
            .O(N__23689),
            .I(N__23683));
    LocalMux I__3665 (
            .O(N__23686),
            .I(N__23680));
    Span4Mux_v I__3664 (
            .O(N__23683),
            .I(N__23675));
    Span4Mux_v I__3663 (
            .O(N__23680),
            .I(N__23672));
    InMux I__3662 (
            .O(N__23679),
            .I(N__23669));
    InMux I__3661 (
            .O(N__23678),
            .I(N__23666));
    Span4Mux_v I__3660 (
            .O(N__23675),
            .I(N__23663));
    Odrv4 I__3659 (
            .O(N__23672),
            .I(data_in_5_3));
    LocalMux I__3658 (
            .O(N__23669),
            .I(data_in_5_3));
    LocalMux I__3657 (
            .O(N__23666),
            .I(data_in_5_3));
    Odrv4 I__3656 (
            .O(N__23663),
            .I(data_in_5_3));
    CascadeMux I__3655 (
            .O(N__23654),
            .I(\c0.n17715_cascade_ ));
    CascadeMux I__3654 (
            .O(N__23651),
            .I(N__23648));
    InMux I__3653 (
            .O(N__23648),
            .I(N__23645));
    LocalMux I__3652 (
            .O(N__23645),
            .I(N__23642));
    Span4Mux_h I__3651 (
            .O(N__23642),
            .I(N__23638));
    InMux I__3650 (
            .O(N__23641),
            .I(N__23635));
    Span4Mux_v I__3649 (
            .O(N__23638),
            .I(N__23632));
    LocalMux I__3648 (
            .O(N__23635),
            .I(data_out_frame2_15_5));
    Odrv4 I__3647 (
            .O(N__23632),
            .I(data_out_frame2_15_5));
    InMux I__3646 (
            .O(N__23627),
            .I(N__23624));
    LocalMux I__3645 (
            .O(N__23624),
            .I(N__23621));
    Span4Mux_h I__3644 (
            .O(N__23621),
            .I(N__23618));
    Span4Mux_v I__3643 (
            .O(N__23618),
            .I(N__23615));
    Odrv4 I__3642 (
            .O(N__23615),
            .I(\c0.n18540 ));
    InMux I__3641 (
            .O(N__23612),
            .I(n16340));
    InMux I__3640 (
            .O(N__23609),
            .I(n16341));
    InMux I__3639 (
            .O(N__23606),
            .I(bfn_5_32_0_));
    InMux I__3638 (
            .O(N__23603),
            .I(n16343));
    InMux I__3637 (
            .O(N__23600),
            .I(n16344));
    InMux I__3636 (
            .O(N__23597),
            .I(n16345));
    InMux I__3635 (
            .O(N__23594),
            .I(n16346));
    InMux I__3634 (
            .O(N__23591),
            .I(n16347));
    InMux I__3633 (
            .O(N__23588),
            .I(n16348));
    InMux I__3632 (
            .O(N__23585),
            .I(n16330));
    InMux I__3631 (
            .O(N__23582),
            .I(n16331));
    InMux I__3630 (
            .O(N__23579),
            .I(n16332));
    InMux I__3629 (
            .O(N__23576),
            .I(n16333));
    InMux I__3628 (
            .O(N__23573),
            .I(bfn_5_31_0_));
    InMux I__3627 (
            .O(N__23570),
            .I(n16335));
    InMux I__3626 (
            .O(N__23567),
            .I(n16336));
    InMux I__3625 (
            .O(N__23564),
            .I(n16337));
    InMux I__3624 (
            .O(N__23561),
            .I(n16338));
    InMux I__3623 (
            .O(N__23558),
            .I(n16339));
    InMux I__3622 (
            .O(N__23555),
            .I(n16321));
    InMux I__3621 (
            .O(N__23552),
            .I(n16322));
    InMux I__3620 (
            .O(N__23549),
            .I(n16323));
    InMux I__3619 (
            .O(N__23546),
            .I(n16324));
    InMux I__3618 (
            .O(N__23543),
            .I(n16325));
    InMux I__3617 (
            .O(N__23540),
            .I(bfn_5_30_0_));
    InMux I__3616 (
            .O(N__23537),
            .I(n16327));
    InMux I__3615 (
            .O(N__23534),
            .I(n16328));
    InMux I__3614 (
            .O(N__23531),
            .I(n16329));
    InMux I__3613 (
            .O(N__23528),
            .I(N__23524));
    InMux I__3612 (
            .O(N__23527),
            .I(N__23521));
    LocalMux I__3611 (
            .O(N__23524),
            .I(N__23516));
    LocalMux I__3610 (
            .O(N__23521),
            .I(N__23516));
    Span4Mux_v I__3609 (
            .O(N__23516),
            .I(N__23513));
    Odrv4 I__3608 (
            .O(N__23513),
            .I(\c0.n17482 ));
    CascadeMux I__3607 (
            .O(N__23510),
            .I(N__23506));
    InMux I__3606 (
            .O(N__23509),
            .I(N__23503));
    InMux I__3605 (
            .O(N__23506),
            .I(N__23500));
    LocalMux I__3604 (
            .O(N__23503),
            .I(N__23497));
    LocalMux I__3603 (
            .O(N__23500),
            .I(data_out_frame2_9_3));
    Odrv4 I__3602 (
            .O(N__23497),
            .I(data_out_frame2_9_3));
    CascadeMux I__3601 (
            .O(N__23492),
            .I(N__23488));
    CascadeMux I__3600 (
            .O(N__23491),
            .I(N__23485));
    InMux I__3599 (
            .O(N__23488),
            .I(N__23480));
    InMux I__3598 (
            .O(N__23485),
            .I(N__23480));
    LocalMux I__3597 (
            .O(N__23480),
            .I(data_out_frame2_8_3));
    InMux I__3596 (
            .O(N__23477),
            .I(N__23474));
    LocalMux I__3595 (
            .O(N__23474),
            .I(N__23471));
    Odrv12 I__3594 (
            .O(N__23471),
            .I(\c0.n18522 ));
    InMux I__3593 (
            .O(N__23468),
            .I(N__23465));
    LocalMux I__3592 (
            .O(N__23465),
            .I(N__23461));
    InMux I__3591 (
            .O(N__23464),
            .I(N__23458));
    Span4Mux_h I__3590 (
            .O(N__23461),
            .I(N__23455));
    LocalMux I__3589 (
            .O(N__23458),
            .I(\c0.data_out_frame2_0_7 ));
    Odrv4 I__3588 (
            .O(N__23455),
            .I(\c0.data_out_frame2_0_7 ));
    CascadeMux I__3587 (
            .O(N__23450),
            .I(N__23447));
    InMux I__3586 (
            .O(N__23447),
            .I(N__23444));
    LocalMux I__3585 (
            .O(N__23444),
            .I(N__23441));
    Sp12to4 I__3584 (
            .O(N__23441),
            .I(N__23438));
    Odrv12 I__3583 (
            .O(N__23438),
            .I(\c0.n18076 ));
    CascadeMux I__3582 (
            .O(N__23435),
            .I(N__23432));
    InMux I__3581 (
            .O(N__23432),
            .I(N__23428));
    InMux I__3580 (
            .O(N__23431),
            .I(N__23425));
    LocalMux I__3579 (
            .O(N__23428),
            .I(data_out_frame2_9_7));
    LocalMux I__3578 (
            .O(N__23425),
            .I(data_out_frame2_9_7));
    CascadeMux I__3577 (
            .O(N__23420),
            .I(N__23416));
    InMux I__3576 (
            .O(N__23419),
            .I(N__23413));
    InMux I__3575 (
            .O(N__23416),
            .I(N__23410));
    LocalMux I__3574 (
            .O(N__23413),
            .I(data_out_frame2_8_7));
    LocalMux I__3573 (
            .O(N__23410),
            .I(data_out_frame2_8_7));
    InMux I__3572 (
            .O(N__23405),
            .I(N__23402));
    LocalMux I__3571 (
            .O(N__23402),
            .I(N__23399));
    Odrv4 I__3570 (
            .O(N__23399),
            .I(\c0.n18588 ));
    InMux I__3569 (
            .O(N__23396),
            .I(N__23393));
    LocalMux I__3568 (
            .O(N__23393),
            .I(N__23390));
    Odrv4 I__3567 (
            .O(N__23390),
            .I(\c0.n17785 ));
    InMux I__3566 (
            .O(N__23387),
            .I(bfn_5_29_0_));
    InMux I__3565 (
            .O(N__23384),
            .I(n16319));
    InMux I__3564 (
            .O(N__23381),
            .I(n16320));
    InMux I__3563 (
            .O(N__23378),
            .I(N__23374));
    InMux I__3562 (
            .O(N__23377),
            .I(N__23371));
    LocalMux I__3561 (
            .O(N__23374),
            .I(N__23368));
    LocalMux I__3560 (
            .O(N__23371),
            .I(data_out_frame2_9_6));
    Odrv12 I__3559 (
            .O(N__23368),
            .I(data_out_frame2_9_6));
    InMux I__3558 (
            .O(N__23363),
            .I(N__23359));
    InMux I__3557 (
            .O(N__23362),
            .I(N__23356));
    LocalMux I__3556 (
            .O(N__23359),
            .I(data_out_frame2_15_3));
    LocalMux I__3555 (
            .O(N__23356),
            .I(data_out_frame2_15_3));
    CascadeMux I__3554 (
            .O(N__23351),
            .I(N__23347));
    InMux I__3553 (
            .O(N__23350),
            .I(N__23344));
    InMux I__3552 (
            .O(N__23347),
            .I(N__23341));
    LocalMux I__3551 (
            .O(N__23344),
            .I(data_out_frame2_14_3));
    LocalMux I__3550 (
            .O(N__23341),
            .I(data_out_frame2_14_3));
    CascadeMux I__3549 (
            .O(N__23336),
            .I(\c0.n18516_cascade_ ));
    InMux I__3548 (
            .O(N__23333),
            .I(N__23330));
    LocalMux I__3547 (
            .O(N__23330),
            .I(N__23326));
    InMux I__3546 (
            .O(N__23329),
            .I(N__23323));
    Span4Mux_h I__3545 (
            .O(N__23326),
            .I(N__23320));
    LocalMux I__3544 (
            .O(N__23323),
            .I(data_out_frame2_13_3));
    Odrv4 I__3543 (
            .O(N__23320),
            .I(data_out_frame2_13_3));
    CascadeMux I__3542 (
            .O(N__23315),
            .I(N__23312));
    InMux I__3541 (
            .O(N__23312),
            .I(N__23308));
    InMux I__3540 (
            .O(N__23311),
            .I(N__23305));
    LocalMux I__3539 (
            .O(N__23308),
            .I(data_out_frame2_11_1));
    LocalMux I__3538 (
            .O(N__23305),
            .I(data_out_frame2_11_1));
    InMux I__3537 (
            .O(N__23300),
            .I(N__23296));
    InMux I__3536 (
            .O(N__23299),
            .I(N__23293));
    LocalMux I__3535 (
            .O(N__23296),
            .I(data_out_frame2_10_1));
    LocalMux I__3534 (
            .O(N__23293),
            .I(data_out_frame2_10_1));
    InMux I__3533 (
            .O(N__23288),
            .I(N__23285));
    LocalMux I__3532 (
            .O(N__23285),
            .I(N__23282));
    Span4Mux_h I__3531 (
            .O(N__23282),
            .I(N__23279));
    Odrv4 I__3530 (
            .O(N__23279),
            .I(\c0.n18480 ));
    InMux I__3529 (
            .O(N__23276),
            .I(N__23273));
    LocalMux I__3528 (
            .O(N__23273),
            .I(\c0.n136 ));
    InMux I__3527 (
            .O(N__23270),
            .I(N__23267));
    LocalMux I__3526 (
            .O(N__23267),
            .I(N__23264));
    Span4Mux_v I__3525 (
            .O(N__23264),
            .I(N__23260));
    InMux I__3524 (
            .O(N__23263),
            .I(N__23257));
    Odrv4 I__3523 (
            .O(N__23260),
            .I(\c0.n1_adj_2443 ));
    LocalMux I__3522 (
            .O(N__23257),
            .I(\c0.n1_adj_2443 ));
    CascadeMux I__3521 (
            .O(N__23252),
            .I(\c0.n14631_cascade_ ));
    CascadeMux I__3520 (
            .O(N__23249),
            .I(N__23246));
    InMux I__3519 (
            .O(N__23246),
            .I(N__23243));
    LocalMux I__3518 (
            .O(N__23243),
            .I(N__23239));
    InMux I__3517 (
            .O(N__23242),
            .I(N__23236));
    Span4Mux_h I__3516 (
            .O(N__23239),
            .I(N__23233));
    LocalMux I__3515 (
            .O(N__23236),
            .I(\c0.data_out_frame2_0_2 ));
    Odrv4 I__3514 (
            .O(N__23233),
            .I(\c0.data_out_frame2_0_2 ));
    InMux I__3513 (
            .O(N__23228),
            .I(\c0.tx.n16358 ));
    InMux I__3512 (
            .O(N__23225),
            .I(\c0.tx.n16359 ));
    InMux I__3511 (
            .O(N__23222),
            .I(\c0.tx.n16360 ));
    InMux I__3510 (
            .O(N__23219),
            .I(\c0.tx.n16361 ));
    InMux I__3509 (
            .O(N__23216),
            .I(\c0.tx.n16362 ));
    InMux I__3508 (
            .O(N__23213),
            .I(\c0.tx.n16363 ));
    InMux I__3507 (
            .O(N__23210),
            .I(bfn_5_26_0_));
    InMux I__3506 (
            .O(N__23207),
            .I(N__23203));
    InMux I__3505 (
            .O(N__23206),
            .I(N__23200));
    LocalMux I__3504 (
            .O(N__23203),
            .I(N__23195));
    LocalMux I__3503 (
            .O(N__23200),
            .I(N__23192));
    InMux I__3502 (
            .O(N__23199),
            .I(N__23187));
    InMux I__3501 (
            .O(N__23198),
            .I(N__23187));
    Span4Mux_v I__3500 (
            .O(N__23195),
            .I(N__23184));
    Span4Mux_v I__3499 (
            .O(N__23192),
            .I(N__23181));
    LocalMux I__3498 (
            .O(N__23187),
            .I(\c0.n31 ));
    Odrv4 I__3497 (
            .O(N__23184),
            .I(\c0.n31 ));
    Odrv4 I__3496 (
            .O(N__23181),
            .I(\c0.n31 ));
    CascadeMux I__3495 (
            .O(N__23174),
            .I(\c0.n17582_cascade_ ));
    InMux I__3494 (
            .O(N__23171),
            .I(N__23168));
    LocalMux I__3493 (
            .O(N__23168),
            .I(N__23165));
    Span4Mux_h I__3492 (
            .O(N__23165),
            .I(N__23162));
    Span4Mux_v I__3491 (
            .O(N__23162),
            .I(N__23159));
    Odrv4 I__3490 (
            .O(N__23159),
            .I(\c0.data_out_frame2_20_7 ));
    InMux I__3489 (
            .O(N__23156),
            .I(N__23153));
    LocalMux I__3488 (
            .O(N__23153),
            .I(N__23150));
    Span4Mux_h I__3487 (
            .O(N__23150),
            .I(N__23147));
    Odrv4 I__3486 (
            .O(N__23147),
            .I(n2560));
    InMux I__3485 (
            .O(N__23144),
            .I(N__23141));
    LocalMux I__3484 (
            .O(N__23141),
            .I(N__23138));
    Odrv4 I__3483 (
            .O(N__23138),
            .I(\c0.n17588 ));
    InMux I__3482 (
            .O(N__23135),
            .I(N__23132));
    LocalMux I__3481 (
            .O(N__23132),
            .I(\c0.n17582 ));
    CascadeMux I__3480 (
            .O(N__23129),
            .I(n2560_cascade_));
    InMux I__3479 (
            .O(N__23126),
            .I(N__23122));
    InMux I__3478 (
            .O(N__23125),
            .I(N__23119));
    LocalMux I__3477 (
            .O(N__23122),
            .I(N__23116));
    LocalMux I__3476 (
            .O(N__23119),
            .I(N__23113));
    Odrv12 I__3475 (
            .O(N__23116),
            .I(n17585));
    Odrv4 I__3474 (
            .O(N__23113),
            .I(n17585));
    InMux I__3473 (
            .O(N__23108),
            .I(N__23105));
    LocalMux I__3472 (
            .O(N__23105),
            .I(\c0.n17648 ));
    CascadeMux I__3471 (
            .O(N__23102),
            .I(\c0.n18_cascade_ ));
    InMux I__3470 (
            .O(N__23099),
            .I(N__23095));
    InMux I__3469 (
            .O(N__23098),
            .I(N__23092));
    LocalMux I__3468 (
            .O(N__23095),
            .I(\c0.n17418 ));
    LocalMux I__3467 (
            .O(N__23092),
            .I(\c0.n17418 ));
    InMux I__3466 (
            .O(N__23087),
            .I(N__23084));
    LocalMux I__3465 (
            .O(N__23084),
            .I(N__23080));
    InMux I__3464 (
            .O(N__23083),
            .I(N__23077));
    Odrv4 I__3463 (
            .O(N__23080),
            .I(n2572));
    LocalMux I__3462 (
            .O(N__23077),
            .I(n2572));
    InMux I__3461 (
            .O(N__23072),
            .I(bfn_5_25_0_));
    InMux I__3460 (
            .O(N__23069),
            .I(\c0.tx.n16357 ));
    InMux I__3459 (
            .O(N__23066),
            .I(N__23062));
    InMux I__3458 (
            .O(N__23065),
            .I(N__23059));
    LocalMux I__3457 (
            .O(N__23062),
            .I(N__23056));
    LocalMux I__3456 (
            .O(N__23059),
            .I(\c0.n8695 ));
    Odrv12 I__3455 (
            .O(N__23056),
            .I(\c0.n8695 ));
    InMux I__3454 (
            .O(N__23051),
            .I(N__23047));
    InMux I__3453 (
            .O(N__23050),
            .I(N__23044));
    LocalMux I__3452 (
            .O(N__23047),
            .I(N__23040));
    LocalMux I__3451 (
            .O(N__23044),
            .I(N__23037));
    InMux I__3450 (
            .O(N__23043),
            .I(N__23034));
    Span4Mux_v I__3449 (
            .O(N__23040),
            .I(N__23029));
    Span4Mux_v I__3448 (
            .O(N__23037),
            .I(N__23029));
    LocalMux I__3447 (
            .O(N__23034),
            .I(\c0.data_in_frame_6_6 ));
    Odrv4 I__3446 (
            .O(N__23029),
            .I(\c0.data_in_frame_6_6 ));
    InMux I__3445 (
            .O(N__23024),
            .I(N__23019));
    InMux I__3444 (
            .O(N__23023),
            .I(N__23016));
    InMux I__3443 (
            .O(N__23022),
            .I(N__23013));
    LocalMux I__3442 (
            .O(N__23019),
            .I(N__23010));
    LocalMux I__3441 (
            .O(N__23016),
            .I(N__23007));
    LocalMux I__3440 (
            .O(N__23013),
            .I(N__23004));
    Span4Mux_v I__3439 (
            .O(N__23010),
            .I(N__23001));
    Span4Mux_v I__3438 (
            .O(N__23007),
            .I(N__22998));
    Odrv12 I__3437 (
            .O(N__23004),
            .I(\c0.n9208 ));
    Odrv4 I__3436 (
            .O(N__23001),
            .I(\c0.n9208 ));
    Odrv4 I__3435 (
            .O(N__22998),
            .I(\c0.n9208 ));
    CascadeMux I__3434 (
            .O(N__22991),
            .I(\c0.n22_cascade_ ));
    InMux I__3433 (
            .O(N__22988),
            .I(N__22985));
    LocalMux I__3432 (
            .O(N__22985),
            .I(n16_adj_2656));
    InMux I__3431 (
            .O(N__22982),
            .I(N__22979));
    LocalMux I__3430 (
            .O(N__22979),
            .I(\c0.n17519 ));
    CascadeMux I__3429 (
            .O(N__22976),
            .I(\c0.n24_cascade_ ));
    InMux I__3428 (
            .O(N__22973),
            .I(N__22970));
    LocalMux I__3427 (
            .O(N__22970),
            .I(N__22967));
    Span4Mux_h I__3426 (
            .O(N__22967),
            .I(N__22964));
    Odrv4 I__3425 (
            .O(N__22964),
            .I(\c0.n11_adj_2453 ));
    InMux I__3424 (
            .O(N__22961),
            .I(N__22957));
    InMux I__3423 (
            .O(N__22960),
            .I(N__22954));
    LocalMux I__3422 (
            .O(N__22957),
            .I(N__22949));
    LocalMux I__3421 (
            .O(N__22954),
            .I(N__22946));
    InMux I__3420 (
            .O(N__22953),
            .I(N__22943));
    InMux I__3419 (
            .O(N__22952),
            .I(N__22940));
    Span4Mux_h I__3418 (
            .O(N__22949),
            .I(N__22935));
    Span4Mux_s2_h I__3417 (
            .O(N__22946),
            .I(N__22935));
    LocalMux I__3416 (
            .O(N__22943),
            .I(data_in_frame_8_2));
    LocalMux I__3415 (
            .O(N__22940),
            .I(data_in_frame_8_2));
    Odrv4 I__3414 (
            .O(N__22935),
            .I(data_in_frame_8_2));
    InMux I__3413 (
            .O(N__22928),
            .I(N__22922));
    InMux I__3412 (
            .O(N__22927),
            .I(N__22917));
    InMux I__3411 (
            .O(N__22926),
            .I(N__22917));
    InMux I__3410 (
            .O(N__22925),
            .I(N__22914));
    LocalMux I__3409 (
            .O(N__22922),
            .I(N__22909));
    LocalMux I__3408 (
            .O(N__22917),
            .I(N__22909));
    LocalMux I__3407 (
            .O(N__22914),
            .I(data_in_frame_8_1));
    Odrv4 I__3406 (
            .O(N__22909),
            .I(data_in_frame_8_1));
    InMux I__3405 (
            .O(N__22904),
            .I(N__22897));
    InMux I__3404 (
            .O(N__22903),
            .I(N__22897));
    InMux I__3403 (
            .O(N__22902),
            .I(N__22894));
    LocalMux I__3402 (
            .O(N__22897),
            .I(N__22890));
    LocalMux I__3401 (
            .O(N__22894),
            .I(N__22887));
    InMux I__3400 (
            .O(N__22893),
            .I(N__22884));
    Span4Mux_v I__3399 (
            .O(N__22890),
            .I(N__22881));
    Span4Mux_h I__3398 (
            .O(N__22887),
            .I(N__22876));
    LocalMux I__3397 (
            .O(N__22884),
            .I(N__22876));
    Odrv4 I__3396 (
            .O(N__22881),
            .I(\c0.data_in_frame_6_3 ));
    Odrv4 I__3395 (
            .O(N__22876),
            .I(\c0.data_in_frame_6_3 ));
    InMux I__3394 (
            .O(N__22871),
            .I(N__22865));
    InMux I__3393 (
            .O(N__22870),
            .I(N__22865));
    LocalMux I__3392 (
            .O(N__22865),
            .I(\c0.n17605 ));
    InMux I__3391 (
            .O(N__22862),
            .I(N__22859));
    LocalMux I__3390 (
            .O(N__22859),
            .I(\c0.n20 ));
    InMux I__3389 (
            .O(N__22856),
            .I(N__22853));
    LocalMux I__3388 (
            .O(N__22853),
            .I(N__22850));
    Span4Mux_v I__3387 (
            .O(N__22850),
            .I(N__22847));
    Span4Mux_h I__3386 (
            .O(N__22847),
            .I(N__22843));
    InMux I__3385 (
            .O(N__22846),
            .I(N__22840));
    Span4Mux_s1_h I__3384 (
            .O(N__22843),
            .I(N__22836));
    LocalMux I__3383 (
            .O(N__22840),
            .I(N__22833));
    InMux I__3382 (
            .O(N__22839),
            .I(N__22828));
    Span4Mux_v I__3381 (
            .O(N__22836),
            .I(N__22823));
    Span4Mux_h I__3380 (
            .O(N__22833),
            .I(N__22823));
    InMux I__3379 (
            .O(N__22832),
            .I(N__22820));
    InMux I__3378 (
            .O(N__22831),
            .I(N__22817));
    LocalMux I__3377 (
            .O(N__22828),
            .I(N__22814));
    Odrv4 I__3376 (
            .O(N__22823),
            .I(\c0.data_in_frame_7_6 ));
    LocalMux I__3375 (
            .O(N__22820),
            .I(\c0.data_in_frame_7_6 ));
    LocalMux I__3374 (
            .O(N__22817),
            .I(\c0.data_in_frame_7_6 ));
    Odrv12 I__3373 (
            .O(N__22814),
            .I(\c0.data_in_frame_7_6 ));
    InMux I__3372 (
            .O(N__22805),
            .I(N__22802));
    LocalMux I__3371 (
            .O(N__22802),
            .I(N__22798));
    CascadeMux I__3370 (
            .O(N__22801),
            .I(N__22795));
    Span4Mux_v I__3369 (
            .O(N__22798),
            .I(N__22792));
    InMux I__3368 (
            .O(N__22795),
            .I(N__22789));
    Odrv4 I__3367 (
            .O(N__22792),
            .I(\c0.n9144 ));
    LocalMux I__3366 (
            .O(N__22789),
            .I(\c0.n9144 ));
    InMux I__3365 (
            .O(N__22784),
            .I(N__22780));
    InMux I__3364 (
            .O(N__22783),
            .I(N__22777));
    LocalMux I__3363 (
            .O(N__22780),
            .I(N__22774));
    LocalMux I__3362 (
            .O(N__22777),
            .I(\c0.n8064 ));
    Odrv12 I__3361 (
            .O(N__22774),
            .I(\c0.n8064 ));
    InMux I__3360 (
            .O(N__22769),
            .I(N__22762));
    InMux I__3359 (
            .O(N__22768),
            .I(N__22762));
    InMux I__3358 (
            .O(N__22767),
            .I(N__22759));
    LocalMux I__3357 (
            .O(N__22762),
            .I(N__22756));
    LocalMux I__3356 (
            .O(N__22759),
            .I(N__22752));
    Span4Mux_v I__3355 (
            .O(N__22756),
            .I(N__22749));
    InMux I__3354 (
            .O(N__22755),
            .I(N__22746));
    Span4Mux_v I__3353 (
            .O(N__22752),
            .I(N__22739));
    Span4Mux_h I__3352 (
            .O(N__22749),
            .I(N__22739));
    LocalMux I__3351 (
            .O(N__22746),
            .I(N__22739));
    Odrv4 I__3350 (
            .O(N__22739),
            .I(\c0.n8687 ));
    InMux I__3349 (
            .O(N__22736),
            .I(N__22733));
    LocalMux I__3348 (
            .O(N__22733),
            .I(N__22730));
    Span4Mux_h I__3347 (
            .O(N__22730),
            .I(N__22726));
    InMux I__3346 (
            .O(N__22729),
            .I(N__22723));
    Odrv4 I__3345 (
            .O(N__22726),
            .I(n2585));
    LocalMux I__3344 (
            .O(N__22723),
            .I(n2585));
    InMux I__3343 (
            .O(N__22718),
            .I(N__22715));
    LocalMux I__3342 (
            .O(N__22715),
            .I(\c0.n17 ));
    InMux I__3341 (
            .O(N__22712),
            .I(N__22709));
    LocalMux I__3340 (
            .O(N__22709),
            .I(n2590));
    InMux I__3339 (
            .O(N__22706),
            .I(N__22702));
    CascadeMux I__3338 (
            .O(N__22705),
            .I(N__22699));
    LocalMux I__3337 (
            .O(N__22702),
            .I(N__22696));
    InMux I__3336 (
            .O(N__22699),
            .I(N__22692));
    Span4Mux_h I__3335 (
            .O(N__22696),
            .I(N__22689));
    CascadeMux I__3334 (
            .O(N__22695),
            .I(N__22686));
    LocalMux I__3333 (
            .O(N__22692),
            .I(N__22683));
    Span4Mux_h I__3332 (
            .O(N__22689),
            .I(N__22680));
    InMux I__3331 (
            .O(N__22686),
            .I(N__22677));
    Odrv4 I__3330 (
            .O(N__22683),
            .I(\c0.data_in_frame_7_1 ));
    Odrv4 I__3329 (
            .O(N__22680),
            .I(\c0.data_in_frame_7_1 ));
    LocalMux I__3328 (
            .O(N__22677),
            .I(\c0.data_in_frame_7_1 ));
    InMux I__3327 (
            .O(N__22670),
            .I(N__22665));
    InMux I__3326 (
            .O(N__22669),
            .I(N__22662));
    CascadeMux I__3325 (
            .O(N__22668),
            .I(N__22659));
    LocalMux I__3324 (
            .O(N__22665),
            .I(N__22654));
    LocalMux I__3323 (
            .O(N__22662),
            .I(N__22654));
    InMux I__3322 (
            .O(N__22659),
            .I(N__22650));
    Span4Mux_s3_h I__3321 (
            .O(N__22654),
            .I(N__22647));
    InMux I__3320 (
            .O(N__22653),
            .I(N__22644));
    LocalMux I__3319 (
            .O(N__22650),
            .I(\c0.data_in_frame_1_0 ));
    Odrv4 I__3318 (
            .O(N__22647),
            .I(\c0.data_in_frame_1_0 ));
    LocalMux I__3317 (
            .O(N__22644),
            .I(\c0.data_in_frame_1_0 ));
    InMux I__3316 (
            .O(N__22637),
            .I(N__22632));
    InMux I__3315 (
            .O(N__22636),
            .I(N__22629));
    InMux I__3314 (
            .O(N__22635),
            .I(N__22624));
    LocalMux I__3313 (
            .O(N__22632),
            .I(N__22621));
    LocalMux I__3312 (
            .O(N__22629),
            .I(N__22618));
    InMux I__3311 (
            .O(N__22628),
            .I(N__22615));
    InMux I__3310 (
            .O(N__22627),
            .I(N__22612));
    LocalMux I__3309 (
            .O(N__22624),
            .I(N__22609));
    Span4Mux_s2_h I__3308 (
            .O(N__22621),
            .I(N__22604));
    Span4Mux_h I__3307 (
            .O(N__22618),
            .I(N__22604));
    LocalMux I__3306 (
            .O(N__22615),
            .I(\c0.data_in_frame_4_6 ));
    LocalMux I__3305 (
            .O(N__22612),
            .I(\c0.data_in_frame_4_6 ));
    Odrv4 I__3304 (
            .O(N__22609),
            .I(\c0.data_in_frame_4_6 ));
    Odrv4 I__3303 (
            .O(N__22604),
            .I(\c0.data_in_frame_4_6 ));
    InMux I__3302 (
            .O(N__22595),
            .I(N__22592));
    LocalMux I__3301 (
            .O(N__22592),
            .I(N__22587));
    InMux I__3300 (
            .O(N__22591),
            .I(N__22584));
    CascadeMux I__3299 (
            .O(N__22590),
            .I(N__22581));
    Span4Mux_h I__3298 (
            .O(N__22587),
            .I(N__22577));
    LocalMux I__3297 (
            .O(N__22584),
            .I(N__22574));
    InMux I__3296 (
            .O(N__22581),
            .I(N__22571));
    InMux I__3295 (
            .O(N__22580),
            .I(N__22568));
    Span4Mux_v I__3294 (
            .O(N__22577),
            .I(N__22563));
    Span4Mux_v I__3293 (
            .O(N__22574),
            .I(N__22563));
    LocalMux I__3292 (
            .O(N__22571),
            .I(N__22560));
    LocalMux I__3291 (
            .O(N__22568),
            .I(\c0.data_in_frame_3_0 ));
    Odrv4 I__3290 (
            .O(N__22563),
            .I(\c0.data_in_frame_3_0 ));
    Odrv12 I__3289 (
            .O(N__22560),
            .I(\c0.data_in_frame_3_0 ));
    InMux I__3288 (
            .O(N__22553),
            .I(N__22549));
    InMux I__3287 (
            .O(N__22552),
            .I(N__22545));
    LocalMux I__3286 (
            .O(N__22549),
            .I(N__22539));
    InMux I__3285 (
            .O(N__22548),
            .I(N__22536));
    LocalMux I__3284 (
            .O(N__22545),
            .I(N__22533));
    InMux I__3283 (
            .O(N__22544),
            .I(N__22530));
    InMux I__3282 (
            .O(N__22543),
            .I(N__22525));
    InMux I__3281 (
            .O(N__22542),
            .I(N__22525));
    Span4Mux_v I__3280 (
            .O(N__22539),
            .I(N__22518));
    LocalMux I__3279 (
            .O(N__22536),
            .I(N__22518));
    Span4Mux_v I__3278 (
            .O(N__22533),
            .I(N__22518));
    LocalMux I__3277 (
            .O(N__22530),
            .I(\c0.data_in_frame_4_7 ));
    LocalMux I__3276 (
            .O(N__22525),
            .I(\c0.data_in_frame_4_7 ));
    Odrv4 I__3275 (
            .O(N__22518),
            .I(\c0.data_in_frame_4_7 ));
    InMux I__3274 (
            .O(N__22511),
            .I(N__22508));
    LocalMux I__3273 (
            .O(N__22508),
            .I(N__22505));
    Span4Mux_h I__3272 (
            .O(N__22505),
            .I(N__22502));
    Odrv4 I__3271 (
            .O(N__22502),
            .I(\c0.n17403 ));
    CascadeMux I__3270 (
            .O(N__22499),
            .I(\c0.n17403_cascade_ ));
    InMux I__3269 (
            .O(N__22496),
            .I(N__22493));
    LocalMux I__3268 (
            .O(N__22493),
            .I(N__22489));
    InMux I__3267 (
            .O(N__22492),
            .I(N__22486));
    Span4Mux_v I__3266 (
            .O(N__22489),
            .I(N__22481));
    LocalMux I__3265 (
            .O(N__22486),
            .I(N__22477));
    InMux I__3264 (
            .O(N__22485),
            .I(N__22474));
    InMux I__3263 (
            .O(N__22484),
            .I(N__22471));
    Span4Mux_h I__3262 (
            .O(N__22481),
            .I(N__22468));
    InMux I__3261 (
            .O(N__22480),
            .I(N__22465));
    Span4Mux_h I__3260 (
            .O(N__22477),
            .I(N__22460));
    LocalMux I__3259 (
            .O(N__22474),
            .I(N__22460));
    LocalMux I__3258 (
            .O(N__22471),
            .I(\c0.data_in_frame_2_6 ));
    Odrv4 I__3257 (
            .O(N__22468),
            .I(\c0.data_in_frame_2_6 ));
    LocalMux I__3256 (
            .O(N__22465),
            .I(\c0.data_in_frame_2_6 ));
    Odrv4 I__3255 (
            .O(N__22460),
            .I(\c0.data_in_frame_2_6 ));
    InMux I__3254 (
            .O(N__22451),
            .I(N__22447));
    InMux I__3253 (
            .O(N__22450),
            .I(N__22444));
    LocalMux I__3252 (
            .O(N__22447),
            .I(N__22441));
    LocalMux I__3251 (
            .O(N__22444),
            .I(N__22438));
    Span4Mux_v I__3250 (
            .O(N__22441),
            .I(N__22433));
    Span4Mux_h I__3249 (
            .O(N__22438),
            .I(N__22433));
    Odrv4 I__3248 (
            .O(N__22433),
            .I(n9283));
    CascadeMux I__3247 (
            .O(N__22430),
            .I(n9283_cascade_));
    InMux I__3246 (
            .O(N__22427),
            .I(N__22424));
    LocalMux I__3245 (
            .O(N__22424),
            .I(N__22421));
    Sp12to4 I__3244 (
            .O(N__22421),
            .I(N__22417));
    InMux I__3243 (
            .O(N__22420),
            .I(N__22414));
    Span12Mux_s7_v I__3242 (
            .O(N__22417),
            .I(N__22411));
    LocalMux I__3241 (
            .O(N__22414),
            .I(data_out_frame2_16_7));
    Odrv12 I__3240 (
            .O(N__22411),
            .I(data_out_frame2_16_7));
    InMux I__3239 (
            .O(N__22406),
            .I(N__22402));
    CascadeMux I__3238 (
            .O(N__22405),
            .I(N__22399));
    LocalMux I__3237 (
            .O(N__22402),
            .I(N__22396));
    InMux I__3236 (
            .O(N__22399),
            .I(N__22393));
    Span4Mux_v I__3235 (
            .O(N__22396),
            .I(N__22390));
    LocalMux I__3234 (
            .O(N__22393),
            .I(N__22387));
    Span4Mux_h I__3233 (
            .O(N__22390),
            .I(N__22382));
    Span4Mux_h I__3232 (
            .O(N__22387),
            .I(N__22382));
    Odrv4 I__3231 (
            .O(N__22382),
            .I(\c0.n9219 ));
    InMux I__3230 (
            .O(N__22379),
            .I(N__22376));
    LocalMux I__3229 (
            .O(N__22376),
            .I(N__22372));
    InMux I__3228 (
            .O(N__22375),
            .I(N__22369));
    Span4Mux_h I__3227 (
            .O(N__22372),
            .I(N__22366));
    LocalMux I__3226 (
            .O(N__22369),
            .I(n2593));
    Odrv4 I__3225 (
            .O(N__22366),
            .I(n2593));
    CascadeMux I__3224 (
            .O(N__22361),
            .I(n2593_cascade_));
    InMux I__3223 (
            .O(N__22358),
            .I(N__22355));
    LocalMux I__3222 (
            .O(N__22355),
            .I(\c0.n22_adj_2461 ));
    InMux I__3221 (
            .O(N__22352),
            .I(N__22349));
    LocalMux I__3220 (
            .O(N__22349),
            .I(N__22346));
    Span4Mux_h I__3219 (
            .O(N__22346),
            .I(N__22342));
    InMux I__3218 (
            .O(N__22345),
            .I(N__22339));
    Odrv4 I__3217 (
            .O(N__22342),
            .I(n2586));
    LocalMux I__3216 (
            .O(N__22339),
            .I(n2586));
    InMux I__3215 (
            .O(N__22334),
            .I(N__22330));
    InMux I__3214 (
            .O(N__22333),
            .I(N__22327));
    LocalMux I__3213 (
            .O(N__22330),
            .I(N__22324));
    LocalMux I__3212 (
            .O(N__22327),
            .I(N__22321));
    Span4Mux_v I__3211 (
            .O(N__22324),
            .I(N__22316));
    Span4Mux_v I__3210 (
            .O(N__22321),
            .I(N__22316));
    Odrv4 I__3209 (
            .O(N__22316),
            .I(\c0.n9279 ));
    CascadeMux I__3208 (
            .O(N__22313),
            .I(n2590_cascade_));
    InMux I__3207 (
            .O(N__22310),
            .I(N__22307));
    LocalMux I__3206 (
            .O(N__22307),
            .I(\c0.n10_adj_2450 ));
    CascadeMux I__3205 (
            .O(N__22304),
            .I(N__22301));
    InMux I__3204 (
            .O(N__22301),
            .I(N__22298));
    LocalMux I__3203 (
            .O(N__22298),
            .I(N__22293));
    InMux I__3202 (
            .O(N__22297),
            .I(N__22288));
    InMux I__3201 (
            .O(N__22296),
            .I(N__22288));
    Span4Mux_v I__3200 (
            .O(N__22293),
            .I(N__22285));
    LocalMux I__3199 (
            .O(N__22288),
            .I(data_in_6_3));
    Odrv4 I__3198 (
            .O(N__22285),
            .I(data_in_6_3));
    InMux I__3197 (
            .O(N__22280),
            .I(N__22277));
    LocalMux I__3196 (
            .O(N__22277),
            .I(N__22274));
    Span4Mux_h I__3195 (
            .O(N__22274),
            .I(N__22270));
    InMux I__3194 (
            .O(N__22273),
            .I(N__22267));
    Odrv4 I__3193 (
            .O(N__22270),
            .I(n2596));
    LocalMux I__3192 (
            .O(N__22267),
            .I(n2596));
    InMux I__3191 (
            .O(N__22262),
            .I(N__22258));
    InMux I__3190 (
            .O(N__22261),
            .I(N__22255));
    LocalMux I__3189 (
            .O(N__22258),
            .I(N__22250));
    LocalMux I__3188 (
            .O(N__22255),
            .I(N__22250));
    Span4Mux_v I__3187 (
            .O(N__22250),
            .I(N__22247));
    Odrv4 I__3186 (
            .O(N__22247),
            .I(\c0.n17529 ));
    CascadeMux I__3185 (
            .O(N__22244),
            .I(n2596_cascade_));
    InMux I__3184 (
            .O(N__22241),
            .I(N__22238));
    LocalMux I__3183 (
            .O(N__22238),
            .I(N__22235));
    Span4Mux_h I__3182 (
            .O(N__22235),
            .I(N__22232));
    Odrv4 I__3181 (
            .O(N__22232),
            .I(\c0.n10_adj_2498 ));
    InMux I__3180 (
            .O(N__22229),
            .I(N__22226));
    LocalMux I__3179 (
            .O(N__22226),
            .I(N__22221));
    InMux I__3178 (
            .O(N__22225),
            .I(N__22218));
    InMux I__3177 (
            .O(N__22224),
            .I(N__22215));
    Span4Mux_s3_h I__3176 (
            .O(N__22221),
            .I(N__22212));
    LocalMux I__3175 (
            .O(N__22218),
            .I(N__22209));
    LocalMux I__3174 (
            .O(N__22215),
            .I(\c0.data_in_frame_7_3 ));
    Odrv4 I__3173 (
            .O(N__22212),
            .I(\c0.data_in_frame_7_3 ));
    Odrv12 I__3172 (
            .O(N__22209),
            .I(\c0.data_in_frame_7_3 ));
    InMux I__3171 (
            .O(N__22202),
            .I(N__22196));
    InMux I__3170 (
            .O(N__22201),
            .I(N__22196));
    LocalMux I__3169 (
            .O(N__22196),
            .I(n2588));
    CascadeMux I__3168 (
            .O(N__22193),
            .I(\c0.n8695_cascade_ ));
    InMux I__3167 (
            .O(N__22190),
            .I(N__22187));
    LocalMux I__3166 (
            .O(N__22187),
            .I(N__22184));
    Span4Mux_v I__3165 (
            .O(N__22184),
            .I(N__22180));
    InMux I__3164 (
            .O(N__22183),
            .I(N__22177));
    Odrv4 I__3163 (
            .O(N__22180),
            .I(\c0.n8867 ));
    LocalMux I__3162 (
            .O(N__22177),
            .I(\c0.n8867 ));
    InMux I__3161 (
            .O(N__22172),
            .I(N__22169));
    LocalMux I__3160 (
            .O(N__22169),
            .I(N__22165));
    InMux I__3159 (
            .O(N__22168),
            .I(N__22162));
    Span4Mux_v I__3158 (
            .O(N__22165),
            .I(N__22156));
    LocalMux I__3157 (
            .O(N__22162),
            .I(N__22156));
    InMux I__3156 (
            .O(N__22161),
            .I(N__22152));
    Span4Mux_v I__3155 (
            .O(N__22156),
            .I(N__22149));
    InMux I__3154 (
            .O(N__22155),
            .I(N__22146));
    LocalMux I__3153 (
            .O(N__22152),
            .I(\c0.data_in_frame_0_6 ));
    Odrv4 I__3152 (
            .O(N__22149),
            .I(\c0.data_in_frame_0_6 ));
    LocalMux I__3151 (
            .O(N__22146),
            .I(\c0.data_in_frame_0_6 ));
    InMux I__3150 (
            .O(N__22139),
            .I(N__22135));
    InMux I__3149 (
            .O(N__22138),
            .I(N__22130));
    LocalMux I__3148 (
            .O(N__22135),
            .I(N__22127));
    InMux I__3147 (
            .O(N__22134),
            .I(N__22124));
    CascadeMux I__3146 (
            .O(N__22133),
            .I(N__22121));
    LocalMux I__3145 (
            .O(N__22130),
            .I(N__22114));
    Span4Mux_v I__3144 (
            .O(N__22127),
            .I(N__22114));
    LocalMux I__3143 (
            .O(N__22124),
            .I(N__22114));
    InMux I__3142 (
            .O(N__22121),
            .I(N__22111));
    Span4Mux_h I__3141 (
            .O(N__22114),
            .I(N__22108));
    LocalMux I__3140 (
            .O(N__22111),
            .I(\c0.data_in_frame_3_4 ));
    Odrv4 I__3139 (
            .O(N__22108),
            .I(\c0.data_in_frame_3_4 ));
    InMux I__3138 (
            .O(N__22103),
            .I(N__22099));
    CascadeMux I__3137 (
            .O(N__22102),
            .I(N__22095));
    LocalMux I__3136 (
            .O(N__22099),
            .I(N__22092));
    InMux I__3135 (
            .O(N__22098),
            .I(N__22087));
    InMux I__3134 (
            .O(N__22095),
            .I(N__22087));
    Span4Mux_h I__3133 (
            .O(N__22092),
            .I(N__22083));
    LocalMux I__3132 (
            .O(N__22087),
            .I(N__22080));
    InMux I__3131 (
            .O(N__22086),
            .I(N__22077));
    Sp12to4 I__3130 (
            .O(N__22083),
            .I(N__22074));
    Span4Mux_v I__3129 (
            .O(N__22080),
            .I(N__22071));
    LocalMux I__3128 (
            .O(N__22077),
            .I(data_in_5_0));
    Odrv12 I__3127 (
            .O(N__22074),
            .I(data_in_5_0));
    Odrv4 I__3126 (
            .O(N__22071),
            .I(data_in_5_0));
    CascadeMux I__3125 (
            .O(N__22064),
            .I(N__22060));
    CascadeMux I__3124 (
            .O(N__22063),
            .I(N__22056));
    InMux I__3123 (
            .O(N__22060),
            .I(N__22049));
    InMux I__3122 (
            .O(N__22059),
            .I(N__22049));
    InMux I__3121 (
            .O(N__22056),
            .I(N__22049));
    LocalMux I__3120 (
            .O(N__22049),
            .I(data_in_7_6));
    InMux I__3119 (
            .O(N__22046),
            .I(N__22043));
    LocalMux I__3118 (
            .O(N__22043),
            .I(N__22038));
    CascadeMux I__3117 (
            .O(N__22042),
            .I(N__22035));
    CascadeMux I__3116 (
            .O(N__22041),
            .I(N__22030));
    Span4Mux_h I__3115 (
            .O(N__22038),
            .I(N__22027));
    InMux I__3114 (
            .O(N__22035),
            .I(N__22022));
    InMux I__3113 (
            .O(N__22034),
            .I(N__22022));
    InMux I__3112 (
            .O(N__22033),
            .I(N__22017));
    InMux I__3111 (
            .O(N__22030),
            .I(N__22017));
    Odrv4 I__3110 (
            .O(N__22027),
            .I(\c0.data_in_frame_1_2 ));
    LocalMux I__3109 (
            .O(N__22022),
            .I(\c0.data_in_frame_1_2 ));
    LocalMux I__3108 (
            .O(N__22017),
            .I(\c0.data_in_frame_1_2 ));
    InMux I__3107 (
            .O(N__22010),
            .I(N__22006));
    InMux I__3106 (
            .O(N__22009),
            .I(N__22003));
    LocalMux I__3105 (
            .O(N__22006),
            .I(N__21999));
    LocalMux I__3104 (
            .O(N__22003),
            .I(N__21996));
    InMux I__3103 (
            .O(N__22002),
            .I(N__21993));
    Span4Mux_v I__3102 (
            .O(N__21999),
            .I(N__21990));
    Span4Mux_h I__3101 (
            .O(N__21996),
            .I(N__21985));
    LocalMux I__3100 (
            .O(N__21993),
            .I(N__21985));
    Span4Mux_h I__3099 (
            .O(N__21990),
            .I(N__21982));
    Odrv4 I__3098 (
            .O(N__21985),
            .I(\c0.data_in_frame_6_1 ));
    Odrv4 I__3097 (
            .O(N__21982),
            .I(\c0.data_in_frame_6_1 ));
    InMux I__3096 (
            .O(N__21977),
            .I(N__21973));
    InMux I__3095 (
            .O(N__21976),
            .I(N__21970));
    LocalMux I__3094 (
            .O(N__21973),
            .I(N__21967));
    LocalMux I__3093 (
            .O(N__21970),
            .I(N__21964));
    Span4Mux_h I__3092 (
            .O(N__21967),
            .I(N__21961));
    Span4Mux_v I__3091 (
            .O(N__21964),
            .I(N__21958));
    Odrv4 I__3090 (
            .O(N__21961),
            .I(\c0.n9328 ));
    Odrv4 I__3089 (
            .O(N__21958),
            .I(\c0.n9328 ));
    CascadeMux I__3088 (
            .O(N__21953),
            .I(N__21950));
    InMux I__3087 (
            .O(N__21950),
            .I(N__21947));
    LocalMux I__3086 (
            .O(N__21947),
            .I(N__21943));
    CascadeMux I__3085 (
            .O(N__21946),
            .I(N__21940));
    Span4Mux_v I__3084 (
            .O(N__21943),
            .I(N__21937));
    InMux I__3083 (
            .O(N__21940),
            .I(N__21934));
    Odrv4 I__3082 (
            .O(N__21937),
            .I(\c0.n8645 ));
    LocalMux I__3081 (
            .O(N__21934),
            .I(\c0.n8645 ));
    InMux I__3080 (
            .O(N__21929),
            .I(N__21925));
    InMux I__3079 (
            .O(N__21928),
            .I(N__21922));
    LocalMux I__3078 (
            .O(N__21925),
            .I(N__21919));
    LocalMux I__3077 (
            .O(N__21922),
            .I(N__21916));
    Span12Mux_s4_h I__3076 (
            .O(N__21919),
            .I(N__21913));
    Odrv4 I__3075 (
            .O(N__21916),
            .I(n9100));
    Odrv12 I__3074 (
            .O(N__21913),
            .I(n9100));
    InMux I__3073 (
            .O(N__21908),
            .I(N__21902));
    InMux I__3072 (
            .O(N__21907),
            .I(N__21899));
    InMux I__3071 (
            .O(N__21906),
            .I(N__21896));
    InMux I__3070 (
            .O(N__21905),
            .I(N__21892));
    LocalMux I__3069 (
            .O(N__21902),
            .I(N__21885));
    LocalMux I__3068 (
            .O(N__21899),
            .I(N__21885));
    LocalMux I__3067 (
            .O(N__21896),
            .I(N__21885));
    InMux I__3066 (
            .O(N__21895),
            .I(N__21882));
    LocalMux I__3065 (
            .O(N__21892),
            .I(N__21877));
    Span4Mux_h I__3064 (
            .O(N__21885),
            .I(N__21877));
    LocalMux I__3063 (
            .O(N__21882),
            .I(N__21874));
    Odrv4 I__3062 (
            .O(N__21877),
            .I(\c0.data_in_frame_4_5 ));
    Odrv4 I__3061 (
            .O(N__21874),
            .I(\c0.data_in_frame_4_5 ));
    InMux I__3060 (
            .O(N__21869),
            .I(N__21865));
    CascadeMux I__3059 (
            .O(N__21868),
            .I(N__21862));
    LocalMux I__3058 (
            .O(N__21865),
            .I(N__21859));
    InMux I__3057 (
            .O(N__21862),
            .I(N__21854));
    Span4Mux_h I__3056 (
            .O(N__21859),
            .I(N__21851));
    InMux I__3055 (
            .O(N__21858),
            .I(N__21846));
    InMux I__3054 (
            .O(N__21857),
            .I(N__21846));
    LocalMux I__3053 (
            .O(N__21854),
            .I(\c0.data_in_frame_0_5 ));
    Odrv4 I__3052 (
            .O(N__21851),
            .I(\c0.data_in_frame_0_5 ));
    LocalMux I__3051 (
            .O(N__21846),
            .I(\c0.data_in_frame_0_5 ));
    InMux I__3050 (
            .O(N__21839),
            .I(N__21834));
    CascadeMux I__3049 (
            .O(N__21838),
            .I(N__21830));
    InMux I__3048 (
            .O(N__21837),
            .I(N__21826));
    LocalMux I__3047 (
            .O(N__21834),
            .I(N__21823));
    InMux I__3046 (
            .O(N__21833),
            .I(N__21820));
    InMux I__3045 (
            .O(N__21830),
            .I(N__21817));
    InMux I__3044 (
            .O(N__21829),
            .I(N__21814));
    LocalMux I__3043 (
            .O(N__21826),
            .I(N__21811));
    Span4Mux_s2_h I__3042 (
            .O(N__21823),
            .I(N__21808));
    LocalMux I__3041 (
            .O(N__21820),
            .I(N__21805));
    LocalMux I__3040 (
            .O(N__21817),
            .I(N__21802));
    LocalMux I__3039 (
            .O(N__21814),
            .I(N__21795));
    Span4Mux_v I__3038 (
            .O(N__21811),
            .I(N__21795));
    Span4Mux_v I__3037 (
            .O(N__21808),
            .I(N__21795));
    Span4Mux_v I__3036 (
            .O(N__21805),
            .I(N__21790));
    Span4Mux_h I__3035 (
            .O(N__21802),
            .I(N__21790));
    Odrv4 I__3034 (
            .O(N__21795),
            .I(\c0.data_in_frame_4_4 ));
    Odrv4 I__3033 (
            .O(N__21790),
            .I(\c0.data_in_frame_4_4 ));
    InMux I__3032 (
            .O(N__21785),
            .I(N__21782));
    LocalMux I__3031 (
            .O(N__21782),
            .I(N__21779));
    Span4Mux_h I__3030 (
            .O(N__21779),
            .I(N__21776));
    Odrv4 I__3029 (
            .O(N__21776),
            .I(\c0.n9176 ));
    InMux I__3028 (
            .O(N__21773),
            .I(N__21769));
    InMux I__3027 (
            .O(N__21772),
            .I(N__21765));
    LocalMux I__3026 (
            .O(N__21769),
            .I(N__21761));
    InMux I__3025 (
            .O(N__21768),
            .I(N__21758));
    LocalMux I__3024 (
            .O(N__21765),
            .I(N__21755));
    CascadeMux I__3023 (
            .O(N__21764),
            .I(N__21751));
    Span4Mux_s3_h I__3022 (
            .O(N__21761),
            .I(N__21748));
    LocalMux I__3021 (
            .O(N__21758),
            .I(N__21745));
    Span4Mux_s2_h I__3020 (
            .O(N__21755),
            .I(N__21742));
    InMux I__3019 (
            .O(N__21754),
            .I(N__21737));
    InMux I__3018 (
            .O(N__21751),
            .I(N__21737));
    Odrv4 I__3017 (
            .O(N__21748),
            .I(\c0.data_in_frame_4_2 ));
    Odrv12 I__3016 (
            .O(N__21745),
            .I(\c0.data_in_frame_4_2 ));
    Odrv4 I__3015 (
            .O(N__21742),
            .I(\c0.data_in_frame_4_2 ));
    LocalMux I__3014 (
            .O(N__21737),
            .I(\c0.data_in_frame_4_2 ));
    InMux I__3013 (
            .O(N__21728),
            .I(N__21724));
    InMux I__3012 (
            .O(N__21727),
            .I(N__21719));
    LocalMux I__3011 (
            .O(N__21724),
            .I(N__21715));
    InMux I__3010 (
            .O(N__21723),
            .I(N__21712));
    InMux I__3009 (
            .O(N__21722),
            .I(N__21709));
    LocalMux I__3008 (
            .O(N__21719),
            .I(N__21706));
    InMux I__3007 (
            .O(N__21718),
            .I(N__21703));
    Span4Mux_s1_h I__3006 (
            .O(N__21715),
            .I(N__21700));
    LocalMux I__3005 (
            .O(N__21712),
            .I(\c0.data_in_frame_2_3 ));
    LocalMux I__3004 (
            .O(N__21709),
            .I(\c0.data_in_frame_2_3 ));
    Odrv12 I__3003 (
            .O(N__21706),
            .I(\c0.data_in_frame_2_3 ));
    LocalMux I__3002 (
            .O(N__21703),
            .I(\c0.data_in_frame_2_3 ));
    Odrv4 I__3001 (
            .O(N__21700),
            .I(\c0.data_in_frame_2_3 ));
    CascadeMux I__3000 (
            .O(N__21689),
            .I(\c0.n10_adj_2430_cascade_ ));
    InMux I__2999 (
            .O(N__21686),
            .I(N__21680));
    InMux I__2998 (
            .O(N__21685),
            .I(N__21677));
    InMux I__2997 (
            .O(N__21684),
            .I(N__21674));
    InMux I__2996 (
            .O(N__21683),
            .I(N__21671));
    LocalMux I__2995 (
            .O(N__21680),
            .I(N__21668));
    LocalMux I__2994 (
            .O(N__21677),
            .I(N__21665));
    LocalMux I__2993 (
            .O(N__21674),
            .I(N__21662));
    LocalMux I__2992 (
            .O(N__21671),
            .I(\c0.data_in_frame_4_1 ));
    Odrv4 I__2991 (
            .O(N__21668),
            .I(\c0.data_in_frame_4_1 ));
    Odrv4 I__2990 (
            .O(N__21665),
            .I(\c0.data_in_frame_4_1 ));
    Odrv12 I__2989 (
            .O(N__21662),
            .I(\c0.data_in_frame_4_1 ));
    InMux I__2988 (
            .O(N__21653),
            .I(N__21650));
    LocalMux I__2987 (
            .O(N__21650),
            .I(N__21647));
    Span4Mux_h I__2986 (
            .O(N__21647),
            .I(N__21642));
    InMux I__2985 (
            .O(N__21646),
            .I(N__21637));
    InMux I__2984 (
            .O(N__21645),
            .I(N__21637));
    Odrv4 I__2983 (
            .O(N__21642),
            .I(data_in_0_7));
    LocalMux I__2982 (
            .O(N__21637),
            .I(data_in_0_7));
    CascadeMux I__2981 (
            .O(N__21632),
            .I(\c0.n17697_cascade_ ));
    InMux I__2980 (
            .O(N__21629),
            .I(N__21625));
    InMux I__2979 (
            .O(N__21628),
            .I(N__21621));
    LocalMux I__2978 (
            .O(N__21625),
            .I(N__21618));
    InMux I__2977 (
            .O(N__21624),
            .I(N__21615));
    LocalMux I__2976 (
            .O(N__21621),
            .I(data_in_0_4));
    Odrv12 I__2975 (
            .O(N__21618),
            .I(data_in_0_4));
    LocalMux I__2974 (
            .O(N__21615),
            .I(data_in_0_4));
    InMux I__2973 (
            .O(N__21608),
            .I(N__21602));
    InMux I__2972 (
            .O(N__21607),
            .I(N__21599));
    InMux I__2971 (
            .O(N__21606),
            .I(N__21596));
    CascadeMux I__2970 (
            .O(N__21605),
            .I(N__21593));
    LocalMux I__2969 (
            .O(N__21602),
            .I(N__21589));
    LocalMux I__2968 (
            .O(N__21599),
            .I(N__21584));
    LocalMux I__2967 (
            .O(N__21596),
            .I(N__21584));
    InMux I__2966 (
            .O(N__21593),
            .I(N__21579));
    InMux I__2965 (
            .O(N__21592),
            .I(N__21576));
    Span4Mux_h I__2964 (
            .O(N__21589),
            .I(N__21573));
    Span4Mux_h I__2963 (
            .O(N__21584),
            .I(N__21570));
    InMux I__2962 (
            .O(N__21583),
            .I(N__21565));
    InMux I__2961 (
            .O(N__21582),
            .I(N__21565));
    LocalMux I__2960 (
            .O(N__21579),
            .I(data_in_frame_5_0));
    LocalMux I__2959 (
            .O(N__21576),
            .I(data_in_frame_5_0));
    Odrv4 I__2958 (
            .O(N__21573),
            .I(data_in_frame_5_0));
    Odrv4 I__2957 (
            .O(N__21570),
            .I(data_in_frame_5_0));
    LocalMux I__2956 (
            .O(N__21565),
            .I(data_in_frame_5_0));
    CascadeMux I__2955 (
            .O(N__21554),
            .I(N__21549));
    InMux I__2954 (
            .O(N__21553),
            .I(N__21546));
    InMux I__2953 (
            .O(N__21552),
            .I(N__21543));
    InMux I__2952 (
            .O(N__21549),
            .I(N__21540));
    LocalMux I__2951 (
            .O(N__21546),
            .I(\c0.n9306 ));
    LocalMux I__2950 (
            .O(N__21543),
            .I(\c0.n9306 ));
    LocalMux I__2949 (
            .O(N__21540),
            .I(\c0.n9306 ));
    InMux I__2948 (
            .O(N__21533),
            .I(N__21530));
    LocalMux I__2947 (
            .O(N__21530),
            .I(\c0.tx2.n4 ));
    CascadeMux I__2946 (
            .O(N__21527),
            .I(\c0.tx2.n9568_cascade_ ));
    InMux I__2945 (
            .O(N__21524),
            .I(N__21520));
    InMux I__2944 (
            .O(N__21523),
            .I(N__21517));
    LocalMux I__2943 (
            .O(N__21520),
            .I(\c0.tx2.tx2_active ));
    LocalMux I__2942 (
            .O(N__21517),
            .I(\c0.tx2.tx2_active ));
    InMux I__2941 (
            .O(N__21512),
            .I(N__21509));
    LocalMux I__2940 (
            .O(N__21509),
            .I(\c0.tx2.n23 ));
    InMux I__2939 (
            .O(N__21506),
            .I(N__21502));
    InMux I__2938 (
            .O(N__21505),
            .I(N__21497));
    LocalMux I__2937 (
            .O(N__21502),
            .I(N__21494));
    InMux I__2936 (
            .O(N__21501),
            .I(N__21491));
    InMux I__2935 (
            .O(N__21500),
            .I(N__21488));
    LocalMux I__2934 (
            .O(N__21497),
            .I(\c0.r_SM_Main_2_N_2326_0 ));
    Odrv4 I__2933 (
            .O(N__21494),
            .I(\c0.r_SM_Main_2_N_2326_0 ));
    LocalMux I__2932 (
            .O(N__21491),
            .I(\c0.r_SM_Main_2_N_2326_0 ));
    LocalMux I__2931 (
            .O(N__21488),
            .I(\c0.r_SM_Main_2_N_2326_0 ));
    InMux I__2930 (
            .O(N__21479),
            .I(N__21476));
    LocalMux I__2929 (
            .O(N__21476),
            .I(N__21473));
    Odrv4 I__2928 (
            .O(N__21473),
            .I(\c0.tx2.n17990 ));
    InMux I__2927 (
            .O(N__21470),
            .I(N__21462));
    InMux I__2926 (
            .O(N__21469),
            .I(N__21455));
    InMux I__2925 (
            .O(N__21468),
            .I(N__21455));
    InMux I__2924 (
            .O(N__21467),
            .I(N__21455));
    InMux I__2923 (
            .O(N__21466),
            .I(N__21452));
    InMux I__2922 (
            .O(N__21465),
            .I(N__21449));
    LocalMux I__2921 (
            .O(N__21462),
            .I(N__21444));
    LocalMux I__2920 (
            .O(N__21455),
            .I(N__21444));
    LocalMux I__2919 (
            .O(N__21452),
            .I(\c0.tx2.r_SM_Main_2_N_2323_1 ));
    LocalMux I__2918 (
            .O(N__21449),
            .I(\c0.tx2.r_SM_Main_2_N_2323_1 ));
    Odrv4 I__2917 (
            .O(N__21444),
            .I(\c0.tx2.r_SM_Main_2_N_2323_1 ));
    CascadeMux I__2916 (
            .O(N__21437),
            .I(\c0.tx2.n12_cascade_ ));
    CascadeMux I__2915 (
            .O(N__21434),
            .I(N__21427));
    CascadeMux I__2914 (
            .O(N__21433),
            .I(N__21422));
    CascadeMux I__2913 (
            .O(N__21432),
            .I(N__21418));
    CascadeMux I__2912 (
            .O(N__21431),
            .I(N__21406));
    InMux I__2911 (
            .O(N__21430),
            .I(N__21401));
    InMux I__2910 (
            .O(N__21427),
            .I(N__21401));
    InMux I__2909 (
            .O(N__21426),
            .I(N__21398));
    InMux I__2908 (
            .O(N__21425),
            .I(N__21391));
    InMux I__2907 (
            .O(N__21422),
            .I(N__21391));
    InMux I__2906 (
            .O(N__21421),
            .I(N__21391));
    InMux I__2905 (
            .O(N__21418),
            .I(N__21382));
    InMux I__2904 (
            .O(N__21417),
            .I(N__21382));
    InMux I__2903 (
            .O(N__21416),
            .I(N__21382));
    InMux I__2902 (
            .O(N__21415),
            .I(N__21382));
    InMux I__2901 (
            .O(N__21414),
            .I(N__21379));
    InMux I__2900 (
            .O(N__21413),
            .I(N__21368));
    InMux I__2899 (
            .O(N__21412),
            .I(N__21368));
    InMux I__2898 (
            .O(N__21411),
            .I(N__21368));
    InMux I__2897 (
            .O(N__21410),
            .I(N__21368));
    InMux I__2896 (
            .O(N__21409),
            .I(N__21368));
    InMux I__2895 (
            .O(N__21406),
            .I(N__21365));
    LocalMux I__2894 (
            .O(N__21401),
            .I(N__21360));
    LocalMux I__2893 (
            .O(N__21398),
            .I(N__21360));
    LocalMux I__2892 (
            .O(N__21391),
            .I(r_SM_Main_2_adj_2628));
    LocalMux I__2891 (
            .O(N__21382),
            .I(r_SM_Main_2_adj_2628));
    LocalMux I__2890 (
            .O(N__21379),
            .I(r_SM_Main_2_adj_2628));
    LocalMux I__2889 (
            .O(N__21368),
            .I(r_SM_Main_2_adj_2628));
    LocalMux I__2888 (
            .O(N__21365),
            .I(r_SM_Main_2_adj_2628));
    Odrv4 I__2887 (
            .O(N__21360),
            .I(r_SM_Main_2_adj_2628));
    InMux I__2886 (
            .O(N__21347),
            .I(N__21344));
    LocalMux I__2885 (
            .O(N__21344),
            .I(N__21337));
    InMux I__2884 (
            .O(N__21343),
            .I(N__21330));
    InMux I__2883 (
            .O(N__21342),
            .I(N__21330));
    InMux I__2882 (
            .O(N__21341),
            .I(N__21330));
    InMux I__2881 (
            .O(N__21340),
            .I(N__21327));
    Span4Mux_s3_h I__2880 (
            .O(N__21337),
            .I(N__21320));
    LocalMux I__2879 (
            .O(N__21330),
            .I(N__21315));
    LocalMux I__2878 (
            .O(N__21327),
            .I(N__21315));
    InMux I__2877 (
            .O(N__21326),
            .I(N__21312));
    InMux I__2876 (
            .O(N__21325),
            .I(N__21305));
    InMux I__2875 (
            .O(N__21324),
            .I(N__21305));
    InMux I__2874 (
            .O(N__21323),
            .I(N__21305));
    Odrv4 I__2873 (
            .O(N__21320),
            .I(\c0.tx2.r_SM_Main_0 ));
    Odrv12 I__2872 (
            .O(N__21315),
            .I(\c0.tx2.r_SM_Main_0 ));
    LocalMux I__2871 (
            .O(N__21312),
            .I(\c0.tx2.r_SM_Main_0 ));
    LocalMux I__2870 (
            .O(N__21305),
            .I(\c0.tx2.r_SM_Main_0 ));
    CascadeMux I__2869 (
            .O(N__21296),
            .I(N__21289));
    CascadeMux I__2868 (
            .O(N__21295),
            .I(N__21285));
    CascadeMux I__2867 (
            .O(N__21294),
            .I(N__21280));
    InMux I__2866 (
            .O(N__21293),
            .I(N__21276));
    InMux I__2865 (
            .O(N__21292),
            .I(N__21267));
    InMux I__2864 (
            .O(N__21289),
            .I(N__21267));
    InMux I__2863 (
            .O(N__21288),
            .I(N__21267));
    InMux I__2862 (
            .O(N__21285),
            .I(N__21267));
    InMux I__2861 (
            .O(N__21284),
            .I(N__21261));
    InMux I__2860 (
            .O(N__21283),
            .I(N__21261));
    InMux I__2859 (
            .O(N__21280),
            .I(N__21258));
    InMux I__2858 (
            .O(N__21279),
            .I(N__21255));
    LocalMux I__2857 (
            .O(N__21276),
            .I(N__21250));
    LocalMux I__2856 (
            .O(N__21267),
            .I(N__21250));
    InMux I__2855 (
            .O(N__21266),
            .I(N__21247));
    LocalMux I__2854 (
            .O(N__21261),
            .I(\c0.tx2.r_SM_Main_1 ));
    LocalMux I__2853 (
            .O(N__21258),
            .I(\c0.tx2.r_SM_Main_1 ));
    LocalMux I__2852 (
            .O(N__21255),
            .I(\c0.tx2.r_SM_Main_1 ));
    Odrv4 I__2851 (
            .O(N__21250),
            .I(\c0.tx2.r_SM_Main_1 ));
    LocalMux I__2850 (
            .O(N__21247),
            .I(\c0.tx2.r_SM_Main_1 ));
    CascadeMux I__2849 (
            .O(N__21236),
            .I(\c0.tx2.n6812_cascade_ ));
    InMux I__2848 (
            .O(N__21233),
            .I(N__21229));
    InMux I__2847 (
            .O(N__21232),
            .I(N__21226));
    LocalMux I__2846 (
            .O(N__21229),
            .I(data_out_frame2_18_7));
    LocalMux I__2845 (
            .O(N__21226),
            .I(data_out_frame2_18_7));
    CascadeMux I__2844 (
            .O(N__21221),
            .I(N__21218));
    InMux I__2843 (
            .O(N__21218),
            .I(N__21215));
    LocalMux I__2842 (
            .O(N__21215),
            .I(N__21212));
    Odrv12 I__2841 (
            .O(N__21212),
            .I(\c0.data_out_frame2_19_7 ));
    CascadeMux I__2840 (
            .O(N__21209),
            .I(\c0.n18576_cascade_ ));
    InMux I__2839 (
            .O(N__21206),
            .I(N__21202));
    InMux I__2838 (
            .O(N__21205),
            .I(N__21199));
    LocalMux I__2837 (
            .O(N__21202),
            .I(N__21196));
    LocalMux I__2836 (
            .O(N__21199),
            .I(data_out_frame2_17_7));
    Odrv4 I__2835 (
            .O(N__21196),
            .I(data_out_frame2_17_7));
    CascadeMux I__2834 (
            .O(N__21191),
            .I(\c0.n18579_cascade_ ));
    InMux I__2833 (
            .O(N__21188),
            .I(N__21185));
    LocalMux I__2832 (
            .O(N__21185),
            .I(\c0.n22_adj_2520 ));
    CascadeMux I__2831 (
            .O(N__21182),
            .I(N__21179));
    InMux I__2830 (
            .O(N__21179),
            .I(N__21176));
    LocalMux I__2829 (
            .O(N__21176),
            .I(\c0.n17788 ));
    InMux I__2828 (
            .O(N__21173),
            .I(N__21170));
    LocalMux I__2827 (
            .O(N__21170),
            .I(\c0.n18420 ));
    SRMux I__2826 (
            .O(N__21167),
            .I(N__21164));
    LocalMux I__2825 (
            .O(N__21164),
            .I(\c0.n4_adj_2480 ));
    IoInMux I__2824 (
            .O(N__21161),
            .I(N__21158));
    LocalMux I__2823 (
            .O(N__21158),
            .I(N__21155));
    Odrv12 I__2822 (
            .O(N__21155),
            .I(tx_enable));
    IoInMux I__2821 (
            .O(N__21152),
            .I(N__21149));
    LocalMux I__2820 (
            .O(N__21149),
            .I(N__21145));
    InMux I__2819 (
            .O(N__21148),
            .I(N__21142));
    Span4Mux_s0_h I__2818 (
            .O(N__21145),
            .I(N__21139));
    LocalMux I__2817 (
            .O(N__21142),
            .I(N__21136));
    Span4Mux_v I__2816 (
            .O(N__21139),
            .I(N__21130));
    Span4Mux_v I__2815 (
            .O(N__21136),
            .I(N__21130));
    InMux I__2814 (
            .O(N__21135),
            .I(N__21127));
    Odrv4 I__2813 (
            .O(N__21130),
            .I(tx2_o));
    LocalMux I__2812 (
            .O(N__21127),
            .I(tx2_o));
    IoInMux I__2811 (
            .O(N__21122),
            .I(N__21119));
    LocalMux I__2810 (
            .O(N__21119),
            .I(N__21116));
    IoSpan4Mux I__2809 (
            .O(N__21116),
            .I(N__21113));
    Span4Mux_s3_h I__2808 (
            .O(N__21113),
            .I(N__21110));
    Span4Mux_h I__2807 (
            .O(N__21110),
            .I(N__21107));
    Odrv4 I__2806 (
            .O(N__21107),
            .I(tx2_enable));
    CascadeMux I__2805 (
            .O(N__21104),
            .I(\c0.n17535_cascade_ ));
    CascadeMux I__2804 (
            .O(N__21101),
            .I(N__21098));
    InMux I__2803 (
            .O(N__21098),
            .I(N__21095));
    LocalMux I__2802 (
            .O(N__21095),
            .I(N__21092));
    Span4Mux_s3_h I__2801 (
            .O(N__21092),
            .I(N__21089));
    Odrv4 I__2800 (
            .O(N__21089),
            .I(\c0.data_out_frame2_19_6 ));
    InMux I__2799 (
            .O(N__21086),
            .I(N__21083));
    LocalMux I__2798 (
            .O(N__21083),
            .I(N__21080));
    Odrv4 I__2797 (
            .O(N__21080),
            .I(\c0.n9240 ));
    CascadeMux I__2796 (
            .O(N__21077),
            .I(\c0.n9240_cascade_ ));
    InMux I__2795 (
            .O(N__21074),
            .I(N__21068));
    InMux I__2794 (
            .O(N__21073),
            .I(N__21068));
    LocalMux I__2793 (
            .O(N__21068),
            .I(N__21065));
    Span4Mux_v I__2792 (
            .O(N__21065),
            .I(N__21061));
    InMux I__2791 (
            .O(N__21064),
            .I(N__21058));
    Odrv4 I__2790 (
            .O(N__21061),
            .I(\c0.n9131 ));
    LocalMux I__2789 (
            .O(N__21058),
            .I(\c0.n9131 ));
    CascadeMux I__2788 (
            .O(N__21053),
            .I(\c0.n17409_cascade_ ));
    InMux I__2787 (
            .O(N__21050),
            .I(N__21047));
    LocalMux I__2786 (
            .O(N__21047),
            .I(\c0.n10_adj_2470 ));
    InMux I__2785 (
            .O(N__21044),
            .I(N__21041));
    LocalMux I__2784 (
            .O(N__21041),
            .I(N__21038));
    Span4Mux_s3_v I__2783 (
            .O(N__21038),
            .I(N__21035));
    Odrv4 I__2782 (
            .O(N__21035),
            .I(\c0.data_out_frame2_20_1 ));
    CascadeMux I__2781 (
            .O(N__21032),
            .I(N__21029));
    InMux I__2780 (
            .O(N__21029),
            .I(N__21026));
    LocalMux I__2779 (
            .O(N__21026),
            .I(N__21023));
    Odrv12 I__2778 (
            .O(N__21023),
            .I(\c0.data_out_frame2_19_1 ));
    InMux I__2777 (
            .O(N__21020),
            .I(N__21017));
    LocalMux I__2776 (
            .O(N__21017),
            .I(N__21014));
    Span4Mux_h I__2775 (
            .O(N__21014),
            .I(N__21011));
    Odrv4 I__2774 (
            .O(N__21011),
            .I(\c0.n6_adj_2464 ));
    CascadeMux I__2773 (
            .O(N__21008),
            .I(\c0.n18423_cascade_ ));
    InMux I__2772 (
            .O(N__21005),
            .I(N__21002));
    LocalMux I__2771 (
            .O(N__21002),
            .I(N__20999));
    Odrv4 I__2770 (
            .O(N__20999),
            .I(\c0.tx2.r_Tx_Data_7 ));
    InMux I__2769 (
            .O(N__20996),
            .I(N__20992));
    InMux I__2768 (
            .O(N__20995),
            .I(N__20989));
    LocalMux I__2767 (
            .O(N__20992),
            .I(N__20986));
    LocalMux I__2766 (
            .O(N__20989),
            .I(data_out_frame2_15_4));
    Odrv12 I__2765 (
            .O(N__20986),
            .I(data_out_frame2_15_4));
    InMux I__2764 (
            .O(N__20981),
            .I(N__20977));
    InMux I__2763 (
            .O(N__20980),
            .I(N__20974));
    LocalMux I__2762 (
            .O(N__20977),
            .I(N__20971));
    LocalMux I__2761 (
            .O(N__20974),
            .I(data_out_frame2_12_4));
    Odrv4 I__2760 (
            .O(N__20971),
            .I(data_out_frame2_12_4));
    InMux I__2759 (
            .O(N__20966),
            .I(N__20963));
    LocalMux I__2758 (
            .O(N__20963),
            .I(N__20960));
    Span4Mux_v I__2757 (
            .O(N__20960),
            .I(N__20956));
    InMux I__2756 (
            .O(N__20959),
            .I(N__20953));
    Span4Mux_h I__2755 (
            .O(N__20956),
            .I(N__20950));
    LocalMux I__2754 (
            .O(N__20953),
            .I(data_out_frame2_13_6));
    Odrv4 I__2753 (
            .O(N__20950),
            .I(data_out_frame2_13_6));
    InMux I__2752 (
            .O(N__20945),
            .I(N__20942));
    LocalMux I__2751 (
            .O(N__20942),
            .I(N__20939));
    Span4Mux_v I__2750 (
            .O(N__20939),
            .I(N__20935));
    InMux I__2749 (
            .O(N__20938),
            .I(N__20932));
    Span4Mux_s1_h I__2748 (
            .O(N__20935),
            .I(N__20929));
    LocalMux I__2747 (
            .O(N__20932),
            .I(data_out_frame2_8_0));
    Odrv4 I__2746 (
            .O(N__20929),
            .I(data_out_frame2_8_0));
    InMux I__2745 (
            .O(N__20924),
            .I(N__20920));
    InMux I__2744 (
            .O(N__20923),
            .I(N__20917));
    LocalMux I__2743 (
            .O(N__20920),
            .I(data_out_frame2_10_7));
    LocalMux I__2742 (
            .O(N__20917),
            .I(data_out_frame2_10_7));
    InMux I__2741 (
            .O(N__20912),
            .I(N__20909));
    LocalMux I__2740 (
            .O(N__20909),
            .I(\c0.n17647 ));
    CascadeMux I__2739 (
            .O(N__20906),
            .I(N__20902));
    CascadeMux I__2738 (
            .O(N__20905),
            .I(N__20899));
    InMux I__2737 (
            .O(N__20902),
            .I(N__20894));
    InMux I__2736 (
            .O(N__20899),
            .I(N__20894));
    LocalMux I__2735 (
            .O(N__20894),
            .I(\c0.n8995 ));
    InMux I__2734 (
            .O(N__20891),
            .I(N__20888));
    LocalMux I__2733 (
            .O(N__20888),
            .I(N__20885));
    Span4Mux_h I__2732 (
            .O(N__20885),
            .I(N__20882));
    Odrv4 I__2731 (
            .O(N__20882),
            .I(\c0.n6_adj_2550 ));
    CascadeMux I__2730 (
            .O(N__20879),
            .I(N__20876));
    InMux I__2729 (
            .O(N__20876),
            .I(N__20873));
    LocalMux I__2728 (
            .O(N__20873),
            .I(N__20870));
    Span12Mux_s3_h I__2727 (
            .O(N__20870),
            .I(N__20867));
    Odrv12 I__2726 (
            .O(N__20867),
            .I(\c0.data_out_frame2_20_0 ));
    CascadeMux I__2725 (
            .O(N__20864),
            .I(\c0.n6_adj_2502_cascade_ ));
    InMux I__2724 (
            .O(N__20861),
            .I(N__20858));
    LocalMux I__2723 (
            .O(N__20858),
            .I(N__20855));
    Span4Mux_s3_h I__2722 (
            .O(N__20855),
            .I(N__20852));
    Odrv4 I__2721 (
            .O(N__20852),
            .I(\c0.data_out_frame2_20_2 ));
    CascadeMux I__2720 (
            .O(N__20849),
            .I(N__20846));
    InMux I__2719 (
            .O(N__20846),
            .I(N__20843));
    LocalMux I__2718 (
            .O(N__20843),
            .I(N__20840));
    Span4Mux_s1_h I__2717 (
            .O(N__20840),
            .I(N__20837));
    Odrv4 I__2716 (
            .O(N__20837),
            .I(\c0.data_out_frame2_19_5 ));
    InMux I__2715 (
            .O(N__20834),
            .I(N__20831));
    LocalMux I__2714 (
            .O(N__20831),
            .I(N__20827));
    InMux I__2713 (
            .O(N__20830),
            .I(N__20824));
    Span4Mux_v I__2712 (
            .O(N__20827),
            .I(N__20821));
    LocalMux I__2711 (
            .O(N__20824),
            .I(data_out_frame2_14_0));
    Odrv4 I__2710 (
            .O(N__20821),
            .I(data_out_frame2_14_0));
    InMux I__2709 (
            .O(N__20816),
            .I(N__20813));
    LocalMux I__2708 (
            .O(N__20813),
            .I(N__20809));
    InMux I__2707 (
            .O(N__20812),
            .I(N__20806));
    Span4Mux_h I__2706 (
            .O(N__20809),
            .I(N__20803));
    LocalMux I__2705 (
            .O(N__20806),
            .I(data_out_frame2_18_2));
    Odrv4 I__2704 (
            .O(N__20803),
            .I(data_out_frame2_18_2));
    InMux I__2703 (
            .O(N__20798),
            .I(N__20795));
    LocalMux I__2702 (
            .O(N__20795),
            .I(N__20792));
    Span4Mux_v I__2701 (
            .O(N__20792),
            .I(N__20788));
    InMux I__2700 (
            .O(N__20791),
            .I(N__20785));
    Span4Mux_v I__2699 (
            .O(N__20788),
            .I(N__20782));
    LocalMux I__2698 (
            .O(N__20785),
            .I(data_out_frame2_5_6));
    Odrv4 I__2697 (
            .O(N__20782),
            .I(data_out_frame2_5_6));
    InMux I__2696 (
            .O(N__20777),
            .I(N__20774));
    LocalMux I__2695 (
            .O(N__20774),
            .I(N__20770));
    InMux I__2694 (
            .O(N__20773),
            .I(N__20767));
    Span4Mux_s3_v I__2693 (
            .O(N__20770),
            .I(N__20764));
    LocalMux I__2692 (
            .O(N__20767),
            .I(data_out_frame2_6_3));
    Odrv4 I__2691 (
            .O(N__20764),
            .I(data_out_frame2_6_3));
    CascadeMux I__2690 (
            .O(N__20759),
            .I(N__20756));
    InMux I__2689 (
            .O(N__20756),
            .I(N__20753));
    LocalMux I__2688 (
            .O(N__20753),
            .I(N__20749));
    InMux I__2687 (
            .O(N__20752),
            .I(N__20746));
    Span4Mux_v I__2686 (
            .O(N__20749),
            .I(N__20743));
    LocalMux I__2685 (
            .O(N__20746),
            .I(data_out_frame2_12_6));
    Odrv4 I__2684 (
            .O(N__20743),
            .I(data_out_frame2_12_6));
    CascadeMux I__2683 (
            .O(N__20738),
            .I(\c0.n17647_cascade_ ));
    InMux I__2682 (
            .O(N__20735),
            .I(N__20732));
    LocalMux I__2681 (
            .O(N__20732),
            .I(\c0.n12_adj_2549 ));
    InMux I__2680 (
            .O(N__20729),
            .I(N__20725));
    InMux I__2679 (
            .O(N__20728),
            .I(N__20722));
    LocalMux I__2678 (
            .O(N__20725),
            .I(N__20719));
    LocalMux I__2677 (
            .O(N__20722),
            .I(N__20716));
    Sp12to4 I__2676 (
            .O(N__20719),
            .I(N__20713));
    Span4Mux_s3_h I__2675 (
            .O(N__20716),
            .I(N__20709));
    Span12Mux_v I__2674 (
            .O(N__20713),
            .I(N__20706));
    InMux I__2673 (
            .O(N__20712),
            .I(N__20703));
    Odrv4 I__2672 (
            .O(N__20709),
            .I(data_in_8_5));
    Odrv12 I__2671 (
            .O(N__20706),
            .I(data_in_8_5));
    LocalMux I__2670 (
            .O(N__20703),
            .I(data_in_8_5));
    CascadeMux I__2669 (
            .O(N__20696),
            .I(N__20693));
    InMux I__2668 (
            .O(N__20693),
            .I(N__20690));
    LocalMux I__2667 (
            .O(N__20690),
            .I(N__20686));
    CascadeMux I__2666 (
            .O(N__20689),
            .I(N__20683));
    Span4Mux_v I__2665 (
            .O(N__20686),
            .I(N__20680));
    InMux I__2664 (
            .O(N__20683),
            .I(N__20677));
    Span4Mux_v I__2663 (
            .O(N__20680),
            .I(N__20674));
    LocalMux I__2662 (
            .O(N__20677),
            .I(\c0.n17602 ));
    Odrv4 I__2661 (
            .O(N__20674),
            .I(\c0.n17602 ));
    InMux I__2660 (
            .O(N__20669),
            .I(N__20665));
    InMux I__2659 (
            .O(N__20668),
            .I(N__20662));
    LocalMux I__2658 (
            .O(N__20665),
            .I(N__20659));
    LocalMux I__2657 (
            .O(N__20662),
            .I(N__20656));
    Span4Mux_v I__2656 (
            .O(N__20659),
            .I(N__20653));
    Odrv4 I__2655 (
            .O(N__20656),
            .I(\c0.n30_adj_2489 ));
    Odrv4 I__2654 (
            .O(N__20653),
            .I(\c0.n30_adj_2489 ));
    InMux I__2653 (
            .O(N__20648),
            .I(N__20645));
    LocalMux I__2652 (
            .O(N__20645),
            .I(\c0.n9345 ));
    CascadeMux I__2651 (
            .O(N__20642),
            .I(\c0.n9345_cascade_ ));
    CascadeMux I__2650 (
            .O(N__20639),
            .I(\c0.n10_cascade_ ));
    InMux I__2649 (
            .O(N__20636),
            .I(N__20633));
    LocalMux I__2648 (
            .O(N__20633),
            .I(N__20630));
    Span4Mux_s3_v I__2647 (
            .O(N__20630),
            .I(N__20627));
    Span4Mux_v I__2646 (
            .O(N__20627),
            .I(N__20624));
    Odrv4 I__2645 (
            .O(N__20624),
            .I(\c0.data_out_frame2_20_6 ));
    InMux I__2644 (
            .O(N__20621),
            .I(N__20618));
    LocalMux I__2643 (
            .O(N__20618),
            .I(N__20615));
    Span4Mux_h I__2642 (
            .O(N__20615),
            .I(N__20612));
    Span4Mux_v I__2641 (
            .O(N__20612),
            .I(N__20608));
    InMux I__2640 (
            .O(N__20611),
            .I(N__20605));
    Odrv4 I__2639 (
            .O(N__20608),
            .I(\c0.n9163 ));
    LocalMux I__2638 (
            .O(N__20605),
            .I(\c0.n9163 ));
    InMux I__2637 (
            .O(N__20600),
            .I(N__20596));
    CascadeMux I__2636 (
            .O(N__20599),
            .I(N__20593));
    LocalMux I__2635 (
            .O(N__20596),
            .I(N__20590));
    InMux I__2634 (
            .O(N__20593),
            .I(N__20587));
    Span4Mux_s3_h I__2633 (
            .O(N__20590),
            .I(N__20584));
    LocalMux I__2632 (
            .O(N__20587),
            .I(\c0.n17470 ));
    Odrv4 I__2631 (
            .O(N__20584),
            .I(\c0.n17470 ));
    InMux I__2630 (
            .O(N__20579),
            .I(N__20576));
    LocalMux I__2629 (
            .O(N__20576),
            .I(n9148));
    CascadeMux I__2628 (
            .O(N__20573),
            .I(n9148_cascade_));
    CascadeMux I__2627 (
            .O(N__20570),
            .I(N__20567));
    InMux I__2626 (
            .O(N__20567),
            .I(N__20563));
    InMux I__2625 (
            .O(N__20566),
            .I(N__20560));
    LocalMux I__2624 (
            .O(N__20563),
            .I(N__20557));
    LocalMux I__2623 (
            .O(N__20560),
            .I(N__20553));
    Span4Mux_h I__2622 (
            .O(N__20557),
            .I(N__20550));
    InMux I__2621 (
            .O(N__20556),
            .I(N__20547));
    Span12Mux_h I__2620 (
            .O(N__20553),
            .I(N__20544));
    Odrv4 I__2619 (
            .O(N__20550),
            .I(\c0.n22_adj_2508 ));
    LocalMux I__2618 (
            .O(N__20547),
            .I(\c0.n22_adj_2508 ));
    Odrv12 I__2617 (
            .O(N__20544),
            .I(\c0.n22_adj_2508 ));
    InMux I__2616 (
            .O(N__20537),
            .I(N__20534));
    LocalMux I__2615 (
            .O(N__20534),
            .I(N__20531));
    Odrv12 I__2614 (
            .O(N__20531),
            .I(\c0.n12_adj_2542 ));
    InMux I__2613 (
            .O(N__20528),
            .I(N__20524));
    InMux I__2612 (
            .O(N__20527),
            .I(N__20520));
    LocalMux I__2611 (
            .O(N__20524),
            .I(N__20517));
    CascadeMux I__2610 (
            .O(N__20523),
            .I(N__20514));
    LocalMux I__2609 (
            .O(N__20520),
            .I(N__20510));
    Span4Mux_v I__2608 (
            .O(N__20517),
            .I(N__20507));
    InMux I__2607 (
            .O(N__20514),
            .I(N__20502));
    InMux I__2606 (
            .O(N__20513),
            .I(N__20502));
    Span4Mux_v I__2605 (
            .O(N__20510),
            .I(N__20499));
    Odrv4 I__2604 (
            .O(N__20507),
            .I(\c0.data_in_frame_2_2 ));
    LocalMux I__2603 (
            .O(N__20502),
            .I(\c0.data_in_frame_2_2 ));
    Odrv4 I__2602 (
            .O(N__20499),
            .I(\c0.data_in_frame_2_2 ));
    InMux I__2601 (
            .O(N__20492),
            .I(N__20486));
    InMux I__2600 (
            .O(N__20491),
            .I(N__20486));
    LocalMux I__2599 (
            .O(N__20486),
            .I(N__20483));
    Span4Mux_v I__2598 (
            .O(N__20483),
            .I(N__20478));
    InMux I__2597 (
            .O(N__20482),
            .I(N__20475));
    InMux I__2596 (
            .O(N__20481),
            .I(N__20472));
    Span4Mux_v I__2595 (
            .O(N__20478),
            .I(N__20467));
    LocalMux I__2594 (
            .O(N__20475),
            .I(N__20467));
    LocalMux I__2593 (
            .O(N__20472),
            .I(\c0.n9058 ));
    Odrv4 I__2592 (
            .O(N__20467),
            .I(\c0.n9058 ));
    InMux I__2591 (
            .O(N__20462),
            .I(N__20458));
    InMux I__2590 (
            .O(N__20461),
            .I(N__20455));
    LocalMux I__2589 (
            .O(N__20458),
            .I(N__20452));
    LocalMux I__2588 (
            .O(N__20455),
            .I(N__20449));
    Span4Mux_v I__2587 (
            .O(N__20452),
            .I(N__20446));
    Odrv12 I__2586 (
            .O(N__20449),
            .I(\c0.n17467 ));
    Odrv4 I__2585 (
            .O(N__20446),
            .I(\c0.n17467 ));
    InMux I__2584 (
            .O(N__20441),
            .I(N__20438));
    LocalMux I__2583 (
            .O(N__20438),
            .I(N__20434));
    InMux I__2582 (
            .O(N__20437),
            .I(N__20431));
    Span4Mux_h I__2581 (
            .O(N__20434),
            .I(N__20428));
    LocalMux I__2580 (
            .O(N__20431),
            .I(N__20419));
    Span4Mux_v I__2579 (
            .O(N__20428),
            .I(N__20419));
    InMux I__2578 (
            .O(N__20427),
            .I(N__20414));
    InMux I__2577 (
            .O(N__20426),
            .I(N__20414));
    InMux I__2576 (
            .O(N__20425),
            .I(N__20409));
    InMux I__2575 (
            .O(N__20424),
            .I(N__20409));
    Odrv4 I__2574 (
            .O(N__20419),
            .I(\c0.data_in_frame_4_3 ));
    LocalMux I__2573 (
            .O(N__20414),
            .I(\c0.data_in_frame_4_3 ));
    LocalMux I__2572 (
            .O(N__20409),
            .I(\c0.data_in_frame_4_3 ));
    InMux I__2571 (
            .O(N__20402),
            .I(N__20398));
    InMux I__2570 (
            .O(N__20401),
            .I(N__20395));
    LocalMux I__2569 (
            .O(N__20398),
            .I(N__20392));
    LocalMux I__2568 (
            .O(N__20395),
            .I(N__20389));
    Span4Mux_v I__2567 (
            .O(N__20392),
            .I(N__20386));
    Odrv4 I__2566 (
            .O(N__20389),
            .I(\c0.n17562 ));
    Odrv4 I__2565 (
            .O(N__20386),
            .I(\c0.n17562 ));
    CascadeMux I__2564 (
            .O(N__20381),
            .I(N__20377));
    InMux I__2563 (
            .O(N__20380),
            .I(N__20372));
    InMux I__2562 (
            .O(N__20377),
            .I(N__20369));
    InMux I__2561 (
            .O(N__20376),
            .I(N__20366));
    InMux I__2560 (
            .O(N__20375),
            .I(N__20363));
    LocalMux I__2559 (
            .O(N__20372),
            .I(N__20360));
    LocalMux I__2558 (
            .O(N__20369),
            .I(N__20355));
    LocalMux I__2557 (
            .O(N__20366),
            .I(N__20355));
    LocalMux I__2556 (
            .O(N__20363),
            .I(N__20350));
    Span4Mux_v I__2555 (
            .O(N__20360),
            .I(N__20350));
    Odrv12 I__2554 (
            .O(N__20355),
            .I(data_in_frame_8_7));
    Odrv4 I__2553 (
            .O(N__20350),
            .I(data_in_frame_8_7));
    InMux I__2552 (
            .O(N__20345),
            .I(N__20342));
    LocalMux I__2551 (
            .O(N__20342),
            .I(N__20338));
    InMux I__2550 (
            .O(N__20341),
            .I(N__20335));
    Span4Mux_h I__2549 (
            .O(N__20338),
            .I(N__20332));
    LocalMux I__2548 (
            .O(N__20335),
            .I(data_out_frame2_6_7));
    Odrv4 I__2547 (
            .O(N__20332),
            .I(data_out_frame2_6_7));
    InMux I__2546 (
            .O(N__20327),
            .I(N__20324));
    LocalMux I__2545 (
            .O(N__20324),
            .I(N__20321));
    Span4Mux_v I__2544 (
            .O(N__20321),
            .I(N__20318));
    Span4Mux_v I__2543 (
            .O(N__20318),
            .I(N__20315));
    Odrv4 I__2542 (
            .O(N__20315),
            .I(\c0.n5_adj_2501 ));
    InMux I__2541 (
            .O(N__20312),
            .I(N__20309));
    LocalMux I__2540 (
            .O(N__20309),
            .I(\c0.n17534 ));
    InMux I__2539 (
            .O(N__20306),
            .I(N__20302));
    InMux I__2538 (
            .O(N__20305),
            .I(N__20299));
    LocalMux I__2537 (
            .O(N__20302),
            .I(N__20296));
    LocalMux I__2536 (
            .O(N__20299),
            .I(N__20291));
    Span4Mux_s3_h I__2535 (
            .O(N__20296),
            .I(N__20291));
    Span4Mux_v I__2534 (
            .O(N__20291),
            .I(N__20286));
    InMux I__2533 (
            .O(N__20290),
            .I(N__20281));
    InMux I__2532 (
            .O(N__20289),
            .I(N__20281));
    Odrv4 I__2531 (
            .O(N__20286),
            .I(\c0.n8674 ));
    LocalMux I__2530 (
            .O(N__20281),
            .I(\c0.n8674 ));
    CascadeMux I__2529 (
            .O(N__20276),
            .I(N__20270));
    CascadeMux I__2528 (
            .O(N__20275),
            .I(N__20267));
    CascadeMux I__2527 (
            .O(N__20274),
            .I(N__20262));
    InMux I__2526 (
            .O(N__20273),
            .I(N__20254));
    InMux I__2525 (
            .O(N__20270),
            .I(N__20254));
    InMux I__2524 (
            .O(N__20267),
            .I(N__20254));
    InMux I__2523 (
            .O(N__20266),
            .I(N__20247));
    InMux I__2522 (
            .O(N__20265),
            .I(N__20247));
    InMux I__2521 (
            .O(N__20262),
            .I(N__20247));
    InMux I__2520 (
            .O(N__20261),
            .I(N__20244));
    LocalMux I__2519 (
            .O(N__20254),
            .I(n9419));
    LocalMux I__2518 (
            .O(N__20247),
            .I(n9419));
    LocalMux I__2517 (
            .O(N__20244),
            .I(n9419));
    CascadeMux I__2516 (
            .O(N__20237),
            .I(N__20234));
    InMux I__2515 (
            .O(N__20234),
            .I(N__20231));
    LocalMux I__2514 (
            .O(N__20231),
            .I(N__20228));
    Odrv4 I__2513 (
            .O(N__20228),
            .I(\c0.n8061 ));
    CascadeMux I__2512 (
            .O(N__20225),
            .I(N__20222));
    InMux I__2511 (
            .O(N__20222),
            .I(N__20219));
    LocalMux I__2510 (
            .O(N__20219),
            .I(N__20216));
    Span4Mux_h I__2509 (
            .O(N__20216),
            .I(N__20213));
    Span4Mux_s1_h I__2508 (
            .O(N__20213),
            .I(N__20210));
    Odrv4 I__2507 (
            .O(N__20210),
            .I(\c0.n8857 ));
    InMux I__2506 (
            .O(N__20207),
            .I(N__20204));
    LocalMux I__2505 (
            .O(N__20204),
            .I(\c0.n18_adj_2468 ));
    CascadeMux I__2504 (
            .O(N__20201),
            .I(\c0.n26_adj_2469_cascade_ ));
    InMux I__2503 (
            .O(N__20198),
            .I(N__20195));
    LocalMux I__2502 (
            .O(N__20195),
            .I(N__20192));
    Odrv12 I__2501 (
            .O(N__20192),
            .I(\c0.n30 ));
    CascadeMux I__2500 (
            .O(N__20189),
            .I(\c0.n12_adj_2449_cascade_ ));
    InMux I__2499 (
            .O(N__20186),
            .I(N__20183));
    LocalMux I__2498 (
            .O(N__20183),
            .I(N__20179));
    InMux I__2497 (
            .O(N__20182),
            .I(N__20175));
    Span4Mux_v I__2496 (
            .O(N__20179),
            .I(N__20172));
    InMux I__2495 (
            .O(N__20178),
            .I(N__20169));
    LocalMux I__2494 (
            .O(N__20175),
            .I(N__20166));
    Odrv4 I__2493 (
            .O(N__20172),
            .I(n2598));
    LocalMux I__2492 (
            .O(N__20169),
            .I(n2598));
    Odrv4 I__2491 (
            .O(N__20166),
            .I(n2598));
    InMux I__2490 (
            .O(N__20159),
            .I(N__20156));
    LocalMux I__2489 (
            .O(N__20156),
            .I(N__20153));
    Span4Mux_v I__2488 (
            .O(N__20153),
            .I(N__20150));
    Odrv4 I__2487 (
            .O(N__20150),
            .I(\c0.n23_adj_2462 ));
    CascadeMux I__2486 (
            .O(N__20147),
            .I(\c0.n24_adj_2454_cascade_ ));
    InMux I__2485 (
            .O(N__20144),
            .I(N__20140));
    InMux I__2484 (
            .O(N__20143),
            .I(N__20137));
    LocalMux I__2483 (
            .O(N__20140),
            .I(N__20132));
    LocalMux I__2482 (
            .O(N__20137),
            .I(N__20129));
    InMux I__2481 (
            .O(N__20136),
            .I(N__20126));
    CascadeMux I__2480 (
            .O(N__20135),
            .I(N__20123));
    Span4Mux_s3_h I__2479 (
            .O(N__20132),
            .I(N__20115));
    Span4Mux_s3_h I__2478 (
            .O(N__20129),
            .I(N__20115));
    LocalMux I__2477 (
            .O(N__20126),
            .I(N__20115));
    InMux I__2476 (
            .O(N__20123),
            .I(N__20112));
    InMux I__2475 (
            .O(N__20122),
            .I(N__20109));
    Span4Mux_v I__2474 (
            .O(N__20115),
            .I(N__20104));
    LocalMux I__2473 (
            .O(N__20112),
            .I(N__20104));
    LocalMux I__2472 (
            .O(N__20109),
            .I(data_in_frame_5_3));
    Odrv4 I__2471 (
            .O(N__20104),
            .I(data_in_frame_5_3));
    InMux I__2470 (
            .O(N__20099),
            .I(N__20095));
    InMux I__2469 (
            .O(N__20098),
            .I(N__20090));
    LocalMux I__2468 (
            .O(N__20095),
            .I(N__20087));
    InMux I__2467 (
            .O(N__20094),
            .I(N__20082));
    InMux I__2466 (
            .O(N__20093),
            .I(N__20082));
    LocalMux I__2465 (
            .O(N__20090),
            .I(\c0.data_in_frame_2_7 ));
    Odrv4 I__2464 (
            .O(N__20087),
            .I(\c0.data_in_frame_2_7 ));
    LocalMux I__2463 (
            .O(N__20082),
            .I(\c0.data_in_frame_2_7 ));
    InMux I__2462 (
            .O(N__20075),
            .I(N__20068));
    CascadeMux I__2461 (
            .O(N__20074),
            .I(N__20065));
    InMux I__2460 (
            .O(N__20073),
            .I(N__20062));
    InMux I__2459 (
            .O(N__20072),
            .I(N__20057));
    InMux I__2458 (
            .O(N__20071),
            .I(N__20057));
    LocalMux I__2457 (
            .O(N__20068),
            .I(N__20054));
    InMux I__2456 (
            .O(N__20065),
            .I(N__20051));
    LocalMux I__2455 (
            .O(N__20062),
            .I(N__20048));
    LocalMux I__2454 (
            .O(N__20057),
            .I(N__20045));
    Span4Mux_h I__2453 (
            .O(N__20054),
            .I(N__20036));
    LocalMux I__2452 (
            .O(N__20051),
            .I(N__20036));
    Span4Mux_v I__2451 (
            .O(N__20048),
            .I(N__20036));
    Span4Mux_v I__2450 (
            .O(N__20045),
            .I(N__20036));
    Odrv4 I__2449 (
            .O(N__20036),
            .I(\c0.data_in_frame_7_7 ));
    InMux I__2448 (
            .O(N__20033),
            .I(N__20030));
    LocalMux I__2447 (
            .O(N__20030),
            .I(N__20027));
    Span4Mux_s3_h I__2446 (
            .O(N__20027),
            .I(N__20024));
    Odrv4 I__2445 (
            .O(N__20024),
            .I(n2584));
    InMux I__2444 (
            .O(N__20021),
            .I(N__20018));
    LocalMux I__2443 (
            .O(N__20018),
            .I(N__20015));
    Span4Mux_h I__2442 (
            .O(N__20015),
            .I(N__20012));
    Span4Mux_v I__2441 (
            .O(N__20012),
            .I(N__20009));
    Odrv4 I__2440 (
            .O(N__20009),
            .I(\c0.n9151 ));
    CascadeMux I__2439 (
            .O(N__20006),
            .I(n2584_cascade_));
    InMux I__2438 (
            .O(N__20003),
            .I(N__20000));
    LocalMux I__2437 (
            .O(N__20000),
            .I(\c0.n21_adj_2465 ));
    InMux I__2436 (
            .O(N__19997),
            .I(N__19993));
    InMux I__2435 (
            .O(N__19996),
            .I(N__19990));
    LocalMux I__2434 (
            .O(N__19993),
            .I(N__19987));
    LocalMux I__2433 (
            .O(N__19990),
            .I(N__19984));
    Span4Mux_s3_h I__2432 (
            .O(N__19987),
            .I(N__19981));
    Span4Mux_s3_h I__2431 (
            .O(N__19984),
            .I(N__19978));
    Span4Mux_v I__2430 (
            .O(N__19981),
            .I(N__19975));
    Span4Mux_v I__2429 (
            .O(N__19978),
            .I(N__19972));
    Odrv4 I__2428 (
            .O(N__19975),
            .I(\c0.n8874 ));
    Odrv4 I__2427 (
            .O(N__19972),
            .I(\c0.n8874 ));
    InMux I__2426 (
            .O(N__19967),
            .I(N__19964));
    LocalMux I__2425 (
            .O(N__19964),
            .I(N__19960));
    InMux I__2424 (
            .O(N__19963),
            .I(N__19955));
    Span4Mux_v I__2423 (
            .O(N__19960),
            .I(N__19952));
    InMux I__2422 (
            .O(N__19959),
            .I(N__19947));
    InMux I__2421 (
            .O(N__19958),
            .I(N__19947));
    LocalMux I__2420 (
            .O(N__19955),
            .I(\c0.data_in_frame_1_4 ));
    Odrv4 I__2419 (
            .O(N__19952),
            .I(\c0.data_in_frame_1_4 ));
    LocalMux I__2418 (
            .O(N__19947),
            .I(\c0.data_in_frame_1_4 ));
    CascadeMux I__2417 (
            .O(N__19940),
            .I(\c0.n8874_cascade_ ));
    InMux I__2416 (
            .O(N__19937),
            .I(N__19933));
    InMux I__2415 (
            .O(N__19936),
            .I(N__19930));
    LocalMux I__2414 (
            .O(N__19933),
            .I(\c0.n9349 ));
    LocalMux I__2413 (
            .O(N__19930),
            .I(\c0.n9349 ));
    CascadeMux I__2412 (
            .O(N__19925),
            .I(\c0.n9368_cascade_ ));
    InMux I__2411 (
            .O(N__19922),
            .I(N__19919));
    LocalMux I__2410 (
            .O(N__19919),
            .I(N__19915));
    InMux I__2409 (
            .O(N__19918),
            .I(N__19912));
    Span4Mux_h I__2408 (
            .O(N__19915),
            .I(N__19909));
    LocalMux I__2407 (
            .O(N__19912),
            .I(\c0.n23_adj_2426 ));
    Odrv4 I__2406 (
            .O(N__19909),
            .I(\c0.n23_adj_2426 ));
    CascadeMux I__2405 (
            .O(N__19904),
            .I(N__19899));
    InMux I__2404 (
            .O(N__19903),
            .I(N__19893));
    InMux I__2403 (
            .O(N__19902),
            .I(N__19893));
    InMux I__2402 (
            .O(N__19899),
            .I(N__19888));
    InMux I__2401 (
            .O(N__19898),
            .I(N__19888));
    LocalMux I__2400 (
            .O(N__19893),
            .I(N__19885));
    LocalMux I__2399 (
            .O(N__19888),
            .I(\c0.data_in_frame_1_6 ));
    Odrv4 I__2398 (
            .O(N__19885),
            .I(\c0.data_in_frame_1_6 ));
    InMux I__2397 (
            .O(N__19880),
            .I(N__19877));
    LocalMux I__2396 (
            .O(N__19877),
            .I(N__19874));
    Odrv4 I__2395 (
            .O(N__19874),
            .I(\c0.n17632 ));
    InMux I__2394 (
            .O(N__19871),
            .I(N__19868));
    LocalMux I__2393 (
            .O(N__19868),
            .I(N__19865));
    Span4Mux_s3_h I__2392 (
            .O(N__19865),
            .I(N__19862));
    Odrv4 I__2391 (
            .O(N__19862),
            .I(\c0.n17485 ));
    InMux I__2390 (
            .O(N__19859),
            .I(N__19855));
    CascadeMux I__2389 (
            .O(N__19858),
            .I(N__19852));
    LocalMux I__2388 (
            .O(N__19855),
            .I(N__19848));
    InMux I__2387 (
            .O(N__19852),
            .I(N__19845));
    InMux I__2386 (
            .O(N__19851),
            .I(N__19842));
    Span4Mux_s3_h I__2385 (
            .O(N__19848),
            .I(N__19839));
    LocalMux I__2384 (
            .O(N__19845),
            .I(\c0.data_in_frame_3_1 ));
    LocalMux I__2383 (
            .O(N__19842),
            .I(\c0.data_in_frame_3_1 ));
    Odrv4 I__2382 (
            .O(N__19839),
            .I(\c0.data_in_frame_3_1 ));
    InMux I__2381 (
            .O(N__19832),
            .I(N__19829));
    LocalMux I__2380 (
            .O(N__19829),
            .I(N__19826));
    Odrv12 I__2379 (
            .O(N__19826),
            .I(\c0.n17406 ));
    InMux I__2378 (
            .O(N__19823),
            .I(N__19817));
    InMux I__2377 (
            .O(N__19822),
            .I(N__19817));
    LocalMux I__2376 (
            .O(N__19817),
            .I(\c0.n13530 ));
    InMux I__2375 (
            .O(N__19814),
            .I(N__19811));
    LocalMux I__2374 (
            .O(N__19811),
            .I(N__19808));
    Span4Mux_v I__2373 (
            .O(N__19808),
            .I(N__19804));
    InMux I__2372 (
            .O(N__19807),
            .I(N__19801));
    Odrv4 I__2371 (
            .O(N__19804),
            .I(\c0.n17656 ));
    LocalMux I__2370 (
            .O(N__19801),
            .I(\c0.n17656 ));
    InMux I__2369 (
            .O(N__19796),
            .I(N__19793));
    LocalMux I__2368 (
            .O(N__19793),
            .I(N__19790));
    Odrv4 I__2367 (
            .O(N__19790),
            .I(\c0.n20_adj_2427 ));
    CascadeMux I__2366 (
            .O(N__19787),
            .I(\c0.n10_adj_2428_cascade_ ));
    InMux I__2365 (
            .O(N__19784),
            .I(N__19781));
    LocalMux I__2364 (
            .O(N__19781),
            .I(N__19778));
    Odrv4 I__2363 (
            .O(N__19778),
            .I(\c0.n17442 ));
    InMux I__2362 (
            .O(N__19775),
            .I(N__19772));
    LocalMux I__2361 (
            .O(N__19772),
            .I(N__19769));
    Odrv4 I__2360 (
            .O(N__19769),
            .I(\c0.n17553 ));
    CascadeMux I__2359 (
            .O(N__19766),
            .I(\c0.n17442_cascade_ ));
    InMux I__2358 (
            .O(N__19763),
            .I(N__19760));
    LocalMux I__2357 (
            .O(N__19760),
            .I(N__19757));
    Odrv4 I__2356 (
            .O(N__19757),
            .I(\c0.n17550 ));
    InMux I__2355 (
            .O(N__19754),
            .I(N__19750));
    InMux I__2354 (
            .O(N__19753),
            .I(N__19745));
    LocalMux I__2353 (
            .O(N__19750),
            .I(N__19742));
    InMux I__2352 (
            .O(N__19749),
            .I(N__19737));
    InMux I__2351 (
            .O(N__19748),
            .I(N__19737));
    LocalMux I__2350 (
            .O(N__19745),
            .I(\c0.data_in_frame_4_0 ));
    Odrv4 I__2349 (
            .O(N__19742),
            .I(\c0.data_in_frame_4_0 ));
    LocalMux I__2348 (
            .O(N__19737),
            .I(\c0.data_in_frame_4_0 ));
    CascadeMux I__2347 (
            .O(N__19730),
            .I(N__19726));
    InMux I__2346 (
            .O(N__19729),
            .I(N__19721));
    InMux I__2345 (
            .O(N__19726),
            .I(N__19721));
    LocalMux I__2344 (
            .O(N__19721),
            .I(data_out_frame2_5_3));
    InMux I__2343 (
            .O(N__19718),
            .I(N__19714));
    InMux I__2342 (
            .O(N__19717),
            .I(N__19711));
    LocalMux I__2341 (
            .O(N__19714),
            .I(N__19708));
    LocalMux I__2340 (
            .O(N__19711),
            .I(data_out_frame2_7_3));
    Odrv12 I__2339 (
            .O(N__19708),
            .I(data_out_frame2_7_3));
    InMux I__2338 (
            .O(N__19703),
            .I(N__19700));
    LocalMux I__2337 (
            .O(N__19700),
            .I(\c0.n5_adj_2509 ));
    InMux I__2336 (
            .O(N__19697),
            .I(N__19694));
    LocalMux I__2335 (
            .O(N__19694),
            .I(N__19691));
    Span4Mux_s2_v I__2334 (
            .O(N__19691),
            .I(N__19688));
    Span4Mux_v I__2333 (
            .O(N__19688),
            .I(N__19684));
    InMux I__2332 (
            .O(N__19687),
            .I(N__19681));
    Span4Mux_v I__2331 (
            .O(N__19684),
            .I(N__19678));
    LocalMux I__2330 (
            .O(N__19681),
            .I(\c0.byte_transmit_counter2_5 ));
    Odrv4 I__2329 (
            .O(N__19678),
            .I(\c0.byte_transmit_counter2_5 ));
    InMux I__2328 (
            .O(N__19673),
            .I(N__19670));
    LocalMux I__2327 (
            .O(N__19670),
            .I(N__19667));
    Span4Mux_s2_v I__2326 (
            .O(N__19667),
            .I(N__19664));
    Span4Mux_v I__2325 (
            .O(N__19664),
            .I(N__19660));
    InMux I__2324 (
            .O(N__19663),
            .I(N__19657));
    Span4Mux_v I__2323 (
            .O(N__19660),
            .I(N__19654));
    LocalMux I__2322 (
            .O(N__19657),
            .I(\c0.byte_transmit_counter2_6 ));
    Odrv4 I__2321 (
            .O(N__19654),
            .I(\c0.byte_transmit_counter2_6 ));
    CascadeMux I__2320 (
            .O(N__19649),
            .I(\c0.n18_adj_2544_cascade_ ));
    InMux I__2319 (
            .O(N__19646),
            .I(N__19643));
    LocalMux I__2318 (
            .O(N__19643),
            .I(N__19640));
    Span4Mux_s2_v I__2317 (
            .O(N__19640),
            .I(N__19637));
    Span4Mux_v I__2316 (
            .O(N__19637),
            .I(N__19633));
    InMux I__2315 (
            .O(N__19636),
            .I(N__19630));
    Span4Mux_v I__2314 (
            .O(N__19633),
            .I(N__19627));
    LocalMux I__2313 (
            .O(N__19630),
            .I(\c0.byte_transmit_counter2_7 ));
    Odrv4 I__2312 (
            .O(N__19627),
            .I(\c0.byte_transmit_counter2_7 ));
    CascadeMux I__2311 (
            .O(N__19622),
            .I(\c0.n19_adj_2540_cascade_ ));
    InMux I__2310 (
            .O(N__19619),
            .I(N__19616));
    LocalMux I__2309 (
            .O(N__19616),
            .I(N__19613));
    Span12Mux_s2_h I__2308 (
            .O(N__19613),
            .I(N__19610));
    Odrv12 I__2307 (
            .O(N__19610),
            .I(\c0.tx2_transmit_N_2287 ));
    CascadeMux I__2306 (
            .O(N__19607),
            .I(\c0.tx2_transmit_N_2287_cascade_ ));
    InMux I__2305 (
            .O(N__19604),
            .I(N__19601));
    LocalMux I__2304 (
            .O(N__19601),
            .I(N__19598));
    Odrv4 I__2303 (
            .O(N__19598),
            .I(\c0.n19_adj_2540 ));
    CascadeMux I__2302 (
            .O(N__19595),
            .I(\c0.n67_cascade_ ));
    InMux I__2301 (
            .O(N__19592),
            .I(N__19589));
    LocalMux I__2300 (
            .O(N__19589),
            .I(N__19586));
    Span4Mux_s3_v I__2299 (
            .O(N__19586),
            .I(N__19583));
    Odrv4 I__2298 (
            .O(N__19583),
            .I(\c0.tx2.r_Tx_Data_0 ));
    InMux I__2297 (
            .O(N__19580),
            .I(N__19577));
    LocalMux I__2296 (
            .O(N__19577),
            .I(N__19574));
    Odrv4 I__2295 (
            .O(N__19574),
            .I(\c0.tx2.r_Tx_Data_1 ));
    CascadeMux I__2294 (
            .O(N__19571),
            .I(\c0.tx2.n18612_cascade_ ));
    InMux I__2293 (
            .O(N__19568),
            .I(N__19565));
    LocalMux I__2292 (
            .O(N__19565),
            .I(\c0.tx2.n18615 ));
    InMux I__2291 (
            .O(N__19562),
            .I(N__19559));
    LocalMux I__2290 (
            .O(N__19559),
            .I(\c0.tx2.r_Tx_Data_6 ));
    InMux I__2289 (
            .O(N__19556),
            .I(N__19552));
    InMux I__2288 (
            .O(N__19555),
            .I(N__19549));
    LocalMux I__2287 (
            .O(N__19552),
            .I(data_out_frame2_17_6));
    LocalMux I__2286 (
            .O(N__19549),
            .I(data_out_frame2_17_6));
    InMux I__2285 (
            .O(N__19544),
            .I(N__19541));
    LocalMux I__2284 (
            .O(N__19541),
            .I(N__19537));
    InMux I__2283 (
            .O(N__19540),
            .I(N__19534));
    Span12Mux_s8_v I__2282 (
            .O(N__19537),
            .I(N__19531));
    LocalMux I__2281 (
            .O(N__19534),
            .I(data_out_frame2_13_4));
    Odrv12 I__2280 (
            .O(N__19531),
            .I(data_out_frame2_13_4));
    InMux I__2279 (
            .O(N__19526),
            .I(N__19523));
    LocalMux I__2278 (
            .O(N__19523),
            .I(N__19520));
    Span4Mux_v I__2277 (
            .O(N__19520),
            .I(N__19517));
    Odrv4 I__2276 (
            .O(N__19517),
            .I(\c0.n12 ));
    CascadeMux I__2275 (
            .O(N__19514),
            .I(\c0.n11_cascade_ ));
    InMux I__2274 (
            .O(N__19511),
            .I(N__19508));
    LocalMux I__2273 (
            .O(N__19508),
            .I(N__19505));
    Span4Mux_h I__2272 (
            .O(N__19505),
            .I(N__19502));
    Span4Mux_v I__2271 (
            .O(N__19502),
            .I(N__19499));
    Odrv4 I__2270 (
            .O(N__19499),
            .I(\c0.tx2.r_Tx_Data_5 ));
    InMux I__2269 (
            .O(N__19496),
            .I(N__19493));
    LocalMux I__2268 (
            .O(N__19493),
            .I(\c0.tx2.n18450 ));
    InMux I__2267 (
            .O(N__19490),
            .I(N__19487));
    LocalMux I__2266 (
            .O(N__19487),
            .I(\c0.tx2.n18453 ));
    CascadeMux I__2265 (
            .O(N__19484),
            .I(N__19481));
    InMux I__2264 (
            .O(N__19481),
            .I(N__19478));
    LocalMux I__2263 (
            .O(N__19478),
            .I(N__19475));
    Span4Mux_v I__2262 (
            .O(N__19475),
            .I(N__19471));
    InMux I__2261 (
            .O(N__19474),
            .I(N__19468));
    Span4Mux_s3_v I__2260 (
            .O(N__19471),
            .I(N__19465));
    LocalMux I__2259 (
            .O(N__19468),
            .I(data_out_frame2_19_0));
    Odrv4 I__2258 (
            .O(N__19465),
            .I(data_out_frame2_19_0));
    InMux I__2257 (
            .O(N__19460),
            .I(N__19457));
    LocalMux I__2256 (
            .O(N__19457),
            .I(\c0.n18603 ));
    InMux I__2255 (
            .O(N__19454),
            .I(N__19451));
    LocalMux I__2254 (
            .O(N__19451),
            .I(N__19448));
    Odrv4 I__2253 (
            .O(N__19448),
            .I(\c0.n22_adj_2510 ));
    InMux I__2252 (
            .O(N__19445),
            .I(N__19441));
    InMux I__2251 (
            .O(N__19444),
            .I(N__19438));
    LocalMux I__2250 (
            .O(N__19441),
            .I(N__19435));
    LocalMux I__2249 (
            .O(N__19438),
            .I(data_out_frame2_14_7));
    Odrv12 I__2248 (
            .O(N__19435),
            .I(data_out_frame2_14_7));
    InMux I__2247 (
            .O(N__19430),
            .I(N__19426));
    InMux I__2246 (
            .O(N__19429),
            .I(N__19423));
    LocalMux I__2245 (
            .O(N__19426),
            .I(N__19420));
    LocalMux I__2244 (
            .O(N__19423),
            .I(data_out_frame2_15_7));
    Odrv12 I__2243 (
            .O(N__19420),
            .I(data_out_frame2_15_7));
    InMux I__2242 (
            .O(N__19415),
            .I(N__19409));
    InMux I__2241 (
            .O(N__19414),
            .I(N__19409));
    LocalMux I__2240 (
            .O(N__19409),
            .I(data_out_frame2_12_7));
    CascadeMux I__2239 (
            .O(N__19406),
            .I(\c0.n18582_cascade_ ));
    InMux I__2238 (
            .O(N__19403),
            .I(N__19399));
    InMux I__2237 (
            .O(N__19402),
            .I(N__19396));
    LocalMux I__2236 (
            .O(N__19399),
            .I(N__19393));
    LocalMux I__2235 (
            .O(N__19396),
            .I(data_out_frame2_13_7));
    Odrv4 I__2234 (
            .O(N__19393),
            .I(data_out_frame2_13_7));
    InMux I__2233 (
            .O(N__19388),
            .I(N__19384));
    InMux I__2232 (
            .O(N__19387),
            .I(N__19381));
    LocalMux I__2231 (
            .O(N__19384),
            .I(data_out_frame2_9_2));
    LocalMux I__2230 (
            .O(N__19381),
            .I(data_out_frame2_9_2));
    CascadeMux I__2229 (
            .O(N__19376),
            .I(N__19373));
    InMux I__2228 (
            .O(N__19373),
            .I(N__19369));
    InMux I__2227 (
            .O(N__19372),
            .I(N__19366));
    LocalMux I__2226 (
            .O(N__19369),
            .I(N__19363));
    LocalMux I__2225 (
            .O(N__19366),
            .I(data_out_frame2_8_2));
    Odrv4 I__2224 (
            .O(N__19363),
            .I(data_out_frame2_8_2));
    InMux I__2223 (
            .O(N__19358),
            .I(N__19355));
    LocalMux I__2222 (
            .O(N__19355),
            .I(\c0.n18504 ));
    InMux I__2221 (
            .O(N__19352),
            .I(N__19349));
    LocalMux I__2220 (
            .O(N__19349),
            .I(N__19346));
    Span4Mux_s2_h I__2219 (
            .O(N__19346),
            .I(N__19343));
    Odrv4 I__2218 (
            .O(N__19343),
            .I(\c0.n17824 ));
    InMux I__2217 (
            .O(N__19340),
            .I(N__19337));
    LocalMux I__2216 (
            .O(N__19337),
            .I(N__19334));
    Span4Mux_h I__2215 (
            .O(N__19334),
            .I(N__19331));
    Odrv4 I__2214 (
            .O(N__19331),
            .I(\c0.tx2.r_Tx_Data_2 ));
    CascadeMux I__2213 (
            .O(N__19328),
            .I(N__19325));
    InMux I__2212 (
            .O(N__19325),
            .I(N__19321));
    InMux I__2211 (
            .O(N__19324),
            .I(N__19318));
    LocalMux I__2210 (
            .O(N__19321),
            .I(N__19315));
    LocalMux I__2209 (
            .O(N__19318),
            .I(data_out_frame2_6_0));
    Odrv4 I__2208 (
            .O(N__19315),
            .I(data_out_frame2_6_0));
    InMux I__2207 (
            .O(N__19310),
            .I(N__19306));
    InMux I__2206 (
            .O(N__19309),
            .I(N__19303));
    LocalMux I__2205 (
            .O(N__19306),
            .I(N__19300));
    LocalMux I__2204 (
            .O(N__19303),
            .I(data_out_frame2_7_1));
    Odrv4 I__2203 (
            .O(N__19300),
            .I(data_out_frame2_7_1));
    InMux I__2202 (
            .O(N__19295),
            .I(N__19292));
    LocalMux I__2201 (
            .O(N__19292),
            .I(N__19288));
    InMux I__2200 (
            .O(N__19291),
            .I(N__19285));
    Span4Mux_s2_h I__2199 (
            .O(N__19288),
            .I(N__19282));
    LocalMux I__2198 (
            .O(N__19285),
            .I(data_out_frame2_16_6));
    Odrv4 I__2197 (
            .O(N__19282),
            .I(data_out_frame2_16_6));
    InMux I__2196 (
            .O(N__19277),
            .I(N__19271));
    InMux I__2195 (
            .O(N__19276),
            .I(N__19271));
    LocalMux I__2194 (
            .O(N__19271),
            .I(data_out_frame2_11_7));
    InMux I__2193 (
            .O(N__19268),
            .I(N__19264));
    InMux I__2192 (
            .O(N__19267),
            .I(N__19261));
    LocalMux I__2191 (
            .O(N__19264),
            .I(N__19258));
    LocalMux I__2190 (
            .O(N__19261),
            .I(data_out_frame2_9_1));
    Odrv4 I__2189 (
            .O(N__19258),
            .I(data_out_frame2_9_1));
    CascadeMux I__2188 (
            .O(N__19253),
            .I(N__19249));
    InMux I__2187 (
            .O(N__19252),
            .I(N__19244));
    InMux I__2186 (
            .O(N__19249),
            .I(N__19244));
    LocalMux I__2185 (
            .O(N__19244),
            .I(data_out_frame2_8_1));
    InMux I__2184 (
            .O(N__19241),
            .I(N__19238));
    LocalMux I__2183 (
            .O(N__19238),
            .I(N__19235));
    Span4Mux_s2_h I__2182 (
            .O(N__19235),
            .I(N__19232));
    Odrv4 I__2181 (
            .O(N__19232),
            .I(\c0.n17833 ));
    InMux I__2180 (
            .O(N__19229),
            .I(N__19225));
    InMux I__2179 (
            .O(N__19228),
            .I(N__19222));
    LocalMux I__2178 (
            .O(N__19225),
            .I(N__19219));
    LocalMux I__2177 (
            .O(N__19222),
            .I(N__19216));
    Span4Mux_s3_h I__2176 (
            .O(N__19219),
            .I(N__19213));
    Odrv4 I__2175 (
            .O(N__19216),
            .I(data_out_frame2_6_1));
    Odrv4 I__2174 (
            .O(N__19213),
            .I(data_out_frame2_6_1));
    InMux I__2173 (
            .O(N__19208),
            .I(N__19204));
    InMux I__2172 (
            .O(N__19207),
            .I(N__19201));
    LocalMux I__2171 (
            .O(N__19204),
            .I(N__19198));
    LocalMux I__2170 (
            .O(N__19201),
            .I(data_out_frame2_17_2));
    Odrv4 I__2169 (
            .O(N__19198),
            .I(data_out_frame2_17_2));
    InMux I__2168 (
            .O(N__19193),
            .I(N__19189));
    InMux I__2167 (
            .O(N__19192),
            .I(N__19186));
    LocalMux I__2166 (
            .O(N__19189),
            .I(data_out_frame2_5_7));
    LocalMux I__2165 (
            .O(N__19186),
            .I(data_out_frame2_5_7));
    CascadeMux I__2164 (
            .O(N__19181),
            .I(N__19178));
    InMux I__2163 (
            .O(N__19178),
            .I(N__19175));
    LocalMux I__2162 (
            .O(N__19175),
            .I(N__19171));
    InMux I__2161 (
            .O(N__19174),
            .I(N__19168));
    Span4Mux_v I__2160 (
            .O(N__19171),
            .I(N__19165));
    LocalMux I__2159 (
            .O(N__19168),
            .I(data_out_frame2_6_5));
    Odrv4 I__2158 (
            .O(N__19165),
            .I(data_out_frame2_6_5));
    CascadeMux I__2157 (
            .O(N__19160),
            .I(N__19157));
    InMux I__2156 (
            .O(N__19157),
            .I(N__19154));
    LocalMux I__2155 (
            .O(N__19154),
            .I(N__19150));
    InMux I__2154 (
            .O(N__19153),
            .I(N__19147));
    Span4Mux_s2_h I__2153 (
            .O(N__19150),
            .I(N__19144));
    LocalMux I__2152 (
            .O(N__19147),
            .I(data_out_frame2_12_1));
    Odrv4 I__2151 (
            .O(N__19144),
            .I(data_out_frame2_12_1));
    InMux I__2150 (
            .O(N__19139),
            .I(N__19136));
    LocalMux I__2149 (
            .O(N__19136),
            .I(N__19132));
    InMux I__2148 (
            .O(N__19135),
            .I(N__19129));
    Span4Mux_v I__2147 (
            .O(N__19132),
            .I(N__19126));
    LocalMux I__2146 (
            .O(N__19129),
            .I(data_out_frame2_7_0));
    Odrv4 I__2145 (
            .O(N__19126),
            .I(data_out_frame2_7_0));
    CascadeMux I__2144 (
            .O(N__19121),
            .I(n9606_cascade_));
    InMux I__2143 (
            .O(N__19118),
            .I(N__19114));
    InMux I__2142 (
            .O(N__19117),
            .I(N__19111));
    LocalMux I__2141 (
            .O(N__19114),
            .I(N__19108));
    LocalMux I__2140 (
            .O(N__19111),
            .I(N__19103));
    Span4Mux_v I__2139 (
            .O(N__19108),
            .I(N__19103));
    Odrv4 I__2138 (
            .O(N__19103),
            .I(data_out_frame2_10_5));
    CascadeMux I__2137 (
            .O(N__19100),
            .I(N__19097));
    InMux I__2136 (
            .O(N__19097),
            .I(N__19093));
    InMux I__2135 (
            .O(N__19096),
            .I(N__19090));
    LocalMux I__2134 (
            .O(N__19093),
            .I(N__19087));
    LocalMux I__2133 (
            .O(N__19090),
            .I(data_out_frame2_13_5));
    Odrv4 I__2132 (
            .O(N__19087),
            .I(data_out_frame2_13_5));
    InMux I__2131 (
            .O(N__19082),
            .I(N__19079));
    LocalMux I__2130 (
            .O(N__19079),
            .I(N__19075));
    InMux I__2129 (
            .O(N__19078),
            .I(N__19072));
    Span4Mux_s2_h I__2128 (
            .O(N__19075),
            .I(N__19069));
    LocalMux I__2127 (
            .O(N__19072),
            .I(data_out_frame2_9_0));
    Odrv4 I__2126 (
            .O(N__19069),
            .I(data_out_frame2_9_0));
    CascadeMux I__2125 (
            .O(N__19064),
            .I(\c0.n9151_cascade_ ));
    CascadeMux I__2124 (
            .O(N__19061),
            .I(\c0.n17588_cascade_ ));
    InMux I__2123 (
            .O(N__19058),
            .I(N__19054));
    InMux I__2122 (
            .O(N__19057),
            .I(N__19050));
    LocalMux I__2121 (
            .O(N__19054),
            .I(N__19047));
    InMux I__2120 (
            .O(N__19053),
            .I(N__19044));
    LocalMux I__2119 (
            .O(N__19050),
            .I(N__19041));
    Span4Mux_v I__2118 (
            .O(N__19047),
            .I(N__19038));
    LocalMux I__2117 (
            .O(N__19044),
            .I(data_in_frame_8_5));
    Odrv12 I__2116 (
            .O(N__19041),
            .I(data_in_frame_8_5));
    Odrv4 I__2115 (
            .O(N__19038),
            .I(data_in_frame_8_5));
    InMux I__2114 (
            .O(N__19031),
            .I(N__19028));
    LocalMux I__2113 (
            .O(N__19028),
            .I(\c0.n6_adj_2429 ));
    InMux I__2112 (
            .O(N__19025),
            .I(N__19022));
    LocalMux I__2111 (
            .O(N__19022),
            .I(N__19019));
    Span4Mux_s2_h I__2110 (
            .O(N__19019),
            .I(N__19016));
    Odrv4 I__2109 (
            .O(N__19016),
            .I(\c0.data_out_frame2_20_5 ));
    CascadeMux I__2108 (
            .O(N__19013),
            .I(N__19009));
    InMux I__2107 (
            .O(N__19012),
            .I(N__19006));
    InMux I__2106 (
            .O(N__19009),
            .I(N__19003));
    LocalMux I__2105 (
            .O(N__19006),
            .I(data_out_frame2_12_2));
    LocalMux I__2104 (
            .O(N__19003),
            .I(data_out_frame2_12_2));
    InMux I__2103 (
            .O(N__18998),
            .I(N__18995));
    LocalMux I__2102 (
            .O(N__18995),
            .I(N__18991));
    InMux I__2101 (
            .O(N__18994),
            .I(N__18988));
    Span4Mux_s2_h I__2100 (
            .O(N__18991),
            .I(N__18985));
    LocalMux I__2099 (
            .O(N__18988),
            .I(data_out_frame2_13_1));
    Odrv4 I__2098 (
            .O(N__18985),
            .I(data_out_frame2_13_1));
    InMux I__2097 (
            .O(N__18980),
            .I(N__18977));
    LocalMux I__2096 (
            .O(N__18977),
            .I(N__18974));
    Span4Mux_v I__2095 (
            .O(N__18974),
            .I(N__18971));
    Span4Mux_v I__2094 (
            .O(N__18971),
            .I(N__18968));
    Odrv4 I__2093 (
            .O(N__18968),
            .I(\c0.n17424 ));
    CascadeMux I__2092 (
            .O(N__18965),
            .I(N__18962));
    InMux I__2091 (
            .O(N__18962),
            .I(N__18959));
    LocalMux I__2090 (
            .O(N__18959),
            .I(N__18956));
    Odrv4 I__2089 (
            .O(N__18956),
            .I(\c0.n17569 ));
    InMux I__2088 (
            .O(N__18953),
            .I(N__18950));
    LocalMux I__2087 (
            .O(N__18950),
            .I(\c0.n10_adj_2505 ));
    InMux I__2086 (
            .O(N__18947),
            .I(N__18944));
    LocalMux I__2085 (
            .O(N__18944),
            .I(\c0.n9028 ));
    CascadeMux I__2084 (
            .O(N__18941),
            .I(\c0.n8061_cascade_ ));
    CascadeMux I__2083 (
            .O(N__18938),
            .I(N__18933));
    InMux I__2082 (
            .O(N__18937),
            .I(N__18930));
    InMux I__2081 (
            .O(N__18936),
            .I(N__18927));
    InMux I__2080 (
            .O(N__18933),
            .I(N__18924));
    LocalMux I__2079 (
            .O(N__18930),
            .I(N__18919));
    LocalMux I__2078 (
            .O(N__18927),
            .I(N__18919));
    LocalMux I__2077 (
            .O(N__18924),
            .I(N__18916));
    Span4Mux_s3_h I__2076 (
            .O(N__18919),
            .I(N__18911));
    Span4Mux_s3_h I__2075 (
            .O(N__18916),
            .I(N__18911));
    Odrv4 I__2074 (
            .O(N__18911),
            .I(\c0.data_in_frame_6_4 ));
    InMux I__2073 (
            .O(N__18908),
            .I(N__18904));
    CascadeMux I__2072 (
            .O(N__18907),
            .I(N__18900));
    LocalMux I__2071 (
            .O(N__18904),
            .I(N__18897));
    InMux I__2070 (
            .O(N__18903),
            .I(N__18894));
    InMux I__2069 (
            .O(N__18900),
            .I(N__18891));
    Odrv4 I__2068 (
            .O(N__18897),
            .I(n2595));
    LocalMux I__2067 (
            .O(N__18894),
            .I(n2595));
    LocalMux I__2066 (
            .O(N__18891),
            .I(n2595));
    InMux I__2065 (
            .O(N__18884),
            .I(N__18880));
    CascadeMux I__2064 (
            .O(N__18883),
            .I(N__18877));
    LocalMux I__2063 (
            .O(N__18880),
            .I(N__18873));
    InMux I__2062 (
            .O(N__18877),
            .I(N__18868));
    InMux I__2061 (
            .O(N__18876),
            .I(N__18868));
    Odrv12 I__2060 (
            .O(N__18873),
            .I(\c0.data_in_frame_0_0 ));
    LocalMux I__2059 (
            .O(N__18868),
            .I(\c0.data_in_frame_0_0 ));
    InMux I__2058 (
            .O(N__18863),
            .I(N__18859));
    InMux I__2057 (
            .O(N__18862),
            .I(N__18856));
    LocalMux I__2056 (
            .O(N__18859),
            .I(N__18850));
    LocalMux I__2055 (
            .O(N__18856),
            .I(N__18850));
    InMux I__2054 (
            .O(N__18855),
            .I(N__18847));
    Span4Mux_v I__2053 (
            .O(N__18850),
            .I(N__18842));
    LocalMux I__2052 (
            .O(N__18847),
            .I(N__18842));
    Odrv4 I__2051 (
            .O(N__18842),
            .I(\c0.n2839 ));
    CascadeMux I__2050 (
            .O(N__18839),
            .I(n1396_cascade_));
    CascadeMux I__2049 (
            .O(N__18836),
            .I(n2589_cascade_));
    InMux I__2048 (
            .O(N__18833),
            .I(N__18830));
    LocalMux I__2047 (
            .O(N__18830),
            .I(n2589));
    InMux I__2046 (
            .O(N__18827),
            .I(N__18824));
    LocalMux I__2045 (
            .O(N__18824),
            .I(N__18821));
    Span4Mux_v I__2044 (
            .O(N__18821),
            .I(N__18818));
    Odrv4 I__2043 (
            .O(N__18818),
            .I(\c0.n18558 ));
    CascadeMux I__2042 (
            .O(N__18815),
            .I(N__18812));
    InMux I__2041 (
            .O(N__18812),
            .I(N__18809));
    LocalMux I__2040 (
            .O(N__18809),
            .I(N__18806));
    Span4Mux_s3_v I__2039 (
            .O(N__18806),
            .I(N__18803));
    Span4Mux_v I__2038 (
            .O(N__18803),
            .I(N__18800));
    Odrv4 I__2037 (
            .O(N__18800),
            .I(\c0.n17797 ));
    InMux I__2036 (
            .O(N__18797),
            .I(N__18794));
    LocalMux I__2035 (
            .O(N__18794),
            .I(N__18790));
    InMux I__2034 (
            .O(N__18793),
            .I(N__18786));
    Span4Mux_v I__2033 (
            .O(N__18790),
            .I(N__18783));
    InMux I__2032 (
            .O(N__18789),
            .I(N__18780));
    LocalMux I__2031 (
            .O(N__18786),
            .I(\c0.n25_adj_2491 ));
    Odrv4 I__2030 (
            .O(N__18783),
            .I(\c0.n25_adj_2491 ));
    LocalMux I__2029 (
            .O(N__18780),
            .I(\c0.n25_adj_2491 ));
    InMux I__2028 (
            .O(N__18773),
            .I(N__18770));
    LocalMux I__2027 (
            .O(N__18770),
            .I(N__18764));
    InMux I__2026 (
            .O(N__18769),
            .I(N__18761));
    InMux I__2025 (
            .O(N__18768),
            .I(N__18758));
    InMux I__2024 (
            .O(N__18767),
            .I(N__18755));
    Span4Mux_s2_h I__2023 (
            .O(N__18764),
            .I(N__18750));
    LocalMux I__2022 (
            .O(N__18761),
            .I(N__18750));
    LocalMux I__2021 (
            .O(N__18758),
            .I(data_in_frame_5_5));
    LocalMux I__2020 (
            .O(N__18755),
            .I(data_in_frame_5_5));
    Odrv4 I__2019 (
            .O(N__18750),
            .I(data_in_frame_5_5));
    CascadeMux I__2018 (
            .O(N__18743),
            .I(N__18740));
    InMux I__2017 (
            .O(N__18740),
            .I(N__18736));
    CascadeMux I__2016 (
            .O(N__18739),
            .I(N__18732));
    LocalMux I__2015 (
            .O(N__18736),
            .I(N__18728));
    InMux I__2014 (
            .O(N__18735),
            .I(N__18725));
    InMux I__2013 (
            .O(N__18732),
            .I(N__18722));
    InMux I__2012 (
            .O(N__18731),
            .I(N__18719));
    Span4Mux_v I__2011 (
            .O(N__18728),
            .I(N__18714));
    LocalMux I__2010 (
            .O(N__18725),
            .I(N__18714));
    LocalMux I__2009 (
            .O(N__18722),
            .I(\c0.data_in_frame_2_4 ));
    LocalMux I__2008 (
            .O(N__18719),
            .I(\c0.data_in_frame_2_4 ));
    Odrv4 I__2007 (
            .O(N__18714),
            .I(\c0.data_in_frame_2_4 ));
    InMux I__2006 (
            .O(N__18707),
            .I(N__18700));
    InMux I__2005 (
            .O(N__18706),
            .I(N__18700));
    InMux I__2004 (
            .O(N__18705),
            .I(N__18697));
    LocalMux I__2003 (
            .O(N__18700),
            .I(N__18694));
    LocalMux I__2002 (
            .O(N__18697),
            .I(\c0.data_in_frame_1_5 ));
    Odrv12 I__2001 (
            .O(N__18694),
            .I(\c0.data_in_frame_1_5 ));
    CascadeMux I__2000 (
            .O(N__18689),
            .I(n9419_cascade_));
    InMux I__1999 (
            .O(N__18686),
            .I(N__18683));
    LocalMux I__1998 (
            .O(N__18683),
            .I(\c0.n12_adj_2492 ));
    InMux I__1997 (
            .O(N__18680),
            .I(N__18675));
    InMux I__1996 (
            .O(N__18679),
            .I(N__18672));
    InMux I__1995 (
            .O(N__18678),
            .I(N__18669));
    LocalMux I__1994 (
            .O(N__18675),
            .I(\c0.data_in_frame_0_7 ));
    LocalMux I__1993 (
            .O(N__18672),
            .I(\c0.data_in_frame_0_7 ));
    LocalMux I__1992 (
            .O(N__18669),
            .I(\c0.data_in_frame_0_7 ));
    CascadeMux I__1991 (
            .O(N__18662),
            .I(N__18659));
    InMux I__1990 (
            .O(N__18659),
            .I(N__18654));
    InMux I__1989 (
            .O(N__18658),
            .I(N__18649));
    InMux I__1988 (
            .O(N__18657),
            .I(N__18649));
    LocalMux I__1987 (
            .O(N__18654),
            .I(\c0.data_in_frame_2_0 ));
    LocalMux I__1986 (
            .O(N__18649),
            .I(\c0.data_in_frame_2_0 ));
    CascadeMux I__1985 (
            .O(N__18644),
            .I(\c0.n17553_cascade_ ));
    InMux I__1984 (
            .O(N__18641),
            .I(N__18635));
    InMux I__1983 (
            .O(N__18640),
            .I(N__18632));
    InMux I__1982 (
            .O(N__18639),
            .I(N__18629));
    InMux I__1981 (
            .O(N__18638),
            .I(N__18626));
    LocalMux I__1980 (
            .O(N__18635),
            .I(\c0.data_in_frame_3_7 ));
    LocalMux I__1979 (
            .O(N__18632),
            .I(\c0.data_in_frame_3_7 ));
    LocalMux I__1978 (
            .O(N__18629),
            .I(\c0.data_in_frame_3_7 ));
    LocalMux I__1977 (
            .O(N__18626),
            .I(\c0.data_in_frame_3_7 ));
    CascadeMux I__1976 (
            .O(N__18617),
            .I(\c0.n17406_cascade_ ));
    InMux I__1975 (
            .O(N__18614),
            .I(N__18611));
    LocalMux I__1974 (
            .O(N__18611),
            .I(\c0.tx2.o_Tx_Serial_N_2354 ));
    CascadeMux I__1973 (
            .O(N__18608),
            .I(\c0.tx2.n12306_cascade_ ));
    InMux I__1972 (
            .O(N__18605),
            .I(N__18600));
    InMux I__1971 (
            .O(N__18604),
            .I(N__18595));
    InMux I__1970 (
            .O(N__18603),
            .I(N__18595));
    LocalMux I__1969 (
            .O(N__18600),
            .I(r_Clock_Count_0_adj_2634));
    LocalMux I__1968 (
            .O(N__18595),
            .I(r_Clock_Count_0_adj_2634));
    InMux I__1967 (
            .O(N__18590),
            .I(N__18585));
    InMux I__1966 (
            .O(N__18589),
            .I(N__18582));
    InMux I__1965 (
            .O(N__18588),
            .I(N__18579));
    LocalMux I__1964 (
            .O(N__18585),
            .I(r_Clock_Count_2_adj_2632));
    LocalMux I__1963 (
            .O(N__18582),
            .I(r_Clock_Count_2_adj_2632));
    LocalMux I__1962 (
            .O(N__18579),
            .I(r_Clock_Count_2_adj_2632));
    CascadeMux I__1961 (
            .O(N__18572),
            .I(N__18567));
    InMux I__1960 (
            .O(N__18571),
            .I(N__18564));
    InMux I__1959 (
            .O(N__18570),
            .I(N__18559));
    InMux I__1958 (
            .O(N__18567),
            .I(N__18559));
    LocalMux I__1957 (
            .O(N__18564),
            .I(r_Clock_Count_4_adj_2630));
    LocalMux I__1956 (
            .O(N__18559),
            .I(r_Clock_Count_4_adj_2630));
    InMux I__1955 (
            .O(N__18554),
            .I(N__18549));
    InMux I__1954 (
            .O(N__18553),
            .I(N__18544));
    InMux I__1953 (
            .O(N__18552),
            .I(N__18544));
    LocalMux I__1952 (
            .O(N__18549),
            .I(r_Clock_Count_3_adj_2631));
    LocalMux I__1951 (
            .O(N__18544),
            .I(r_Clock_Count_3_adj_2631));
    InMux I__1950 (
            .O(N__18539),
            .I(N__18534));
    InMux I__1949 (
            .O(N__18538),
            .I(N__18531));
    InMux I__1948 (
            .O(N__18537),
            .I(N__18528));
    LocalMux I__1947 (
            .O(N__18534),
            .I(r_Clock_Count_5_adj_2629));
    LocalMux I__1946 (
            .O(N__18531),
            .I(r_Clock_Count_5_adj_2629));
    LocalMux I__1945 (
            .O(N__18528),
            .I(r_Clock_Count_5_adj_2629));
    CascadeMux I__1944 (
            .O(N__18521),
            .I(\c0.tx2.n10_cascade_ ));
    InMux I__1943 (
            .O(N__18518),
            .I(N__18513));
    InMux I__1942 (
            .O(N__18517),
            .I(N__18510));
    InMux I__1941 (
            .O(N__18516),
            .I(N__18507));
    LocalMux I__1940 (
            .O(N__18513),
            .I(\c0.tx2.r_Clock_Count_7 ));
    LocalMux I__1939 (
            .O(N__18510),
            .I(\c0.tx2.r_Clock_Count_7 ));
    LocalMux I__1938 (
            .O(N__18507),
            .I(\c0.tx2.r_Clock_Count_7 ));
    InMux I__1937 (
            .O(N__18500),
            .I(N__18495));
    InMux I__1936 (
            .O(N__18499),
            .I(N__18492));
    InMux I__1935 (
            .O(N__18498),
            .I(N__18489));
    LocalMux I__1934 (
            .O(N__18495),
            .I(\c0.tx2.r_Clock_Count_6 ));
    LocalMux I__1933 (
            .O(N__18492),
            .I(\c0.tx2.r_Clock_Count_6 ));
    LocalMux I__1932 (
            .O(N__18489),
            .I(\c0.tx2.r_Clock_Count_6 ));
    CascadeMux I__1931 (
            .O(N__18482),
            .I(N__18479));
    InMux I__1930 (
            .O(N__18479),
            .I(N__18474));
    InMux I__1929 (
            .O(N__18478),
            .I(N__18469));
    InMux I__1928 (
            .O(N__18477),
            .I(N__18469));
    LocalMux I__1927 (
            .O(N__18474),
            .I(N__18466));
    LocalMux I__1926 (
            .O(N__18469),
            .I(\c0.tx2.r_Clock_Count_8 ));
    Odrv4 I__1925 (
            .O(N__18466),
            .I(\c0.tx2.r_Clock_Count_8 ));
    InMux I__1924 (
            .O(N__18461),
            .I(N__18458));
    LocalMux I__1923 (
            .O(N__18458),
            .I(\c0.tx2.n16452 ));
    CascadeMux I__1922 (
            .O(N__18455),
            .I(\c0.tx2.r_SM_Main_2_N_2323_1_cascade_ ));
    InMux I__1921 (
            .O(N__18452),
            .I(N__18449));
    LocalMux I__1920 (
            .O(N__18449),
            .I(n320));
    InMux I__1919 (
            .O(N__18446),
            .I(N__18435));
    InMux I__1918 (
            .O(N__18445),
            .I(N__18432));
    InMux I__1917 (
            .O(N__18444),
            .I(N__18423));
    InMux I__1916 (
            .O(N__18443),
            .I(N__18423));
    InMux I__1915 (
            .O(N__18442),
            .I(N__18423));
    InMux I__1914 (
            .O(N__18441),
            .I(N__18423));
    InMux I__1913 (
            .O(N__18440),
            .I(N__18420));
    InMux I__1912 (
            .O(N__18439),
            .I(N__18417));
    InMux I__1911 (
            .O(N__18438),
            .I(N__18414));
    LocalMux I__1910 (
            .O(N__18435),
            .I(n10244));
    LocalMux I__1909 (
            .O(N__18432),
            .I(n10244));
    LocalMux I__1908 (
            .O(N__18423),
            .I(n10244));
    LocalMux I__1907 (
            .O(N__18420),
            .I(n10244));
    LocalMux I__1906 (
            .O(N__18417),
            .I(n10244));
    LocalMux I__1905 (
            .O(N__18414),
            .I(n10244));
    CascadeMux I__1904 (
            .O(N__18401),
            .I(N__18398));
    InMux I__1903 (
            .O(N__18398),
            .I(N__18393));
    InMux I__1902 (
            .O(N__18397),
            .I(N__18390));
    InMux I__1901 (
            .O(N__18396),
            .I(N__18387));
    LocalMux I__1900 (
            .O(N__18393),
            .I(r_Clock_Count_1_adj_2633));
    LocalMux I__1899 (
            .O(N__18390),
            .I(r_Clock_Count_1_adj_2633));
    LocalMux I__1898 (
            .O(N__18387),
            .I(r_Clock_Count_1_adj_2633));
    CascadeMux I__1897 (
            .O(N__18380),
            .I(\c0.n18411_cascade_ ));
    InMux I__1896 (
            .O(N__18377),
            .I(N__18373));
    InMux I__1895 (
            .O(N__18376),
            .I(N__18370));
    LocalMux I__1894 (
            .O(N__18373),
            .I(data_out_frame2_18_6));
    LocalMux I__1893 (
            .O(N__18370),
            .I(data_out_frame2_18_6));
    CascadeMux I__1892 (
            .O(N__18365),
            .I(\c0.n18552_cascade_ ));
    CascadeMux I__1891 (
            .O(N__18362),
            .I(\c0.n18555_cascade_ ));
    InMux I__1890 (
            .O(N__18359),
            .I(N__18356));
    LocalMux I__1889 (
            .O(N__18356),
            .I(\c0.n22_adj_2521 ));
    CascadeMux I__1888 (
            .O(N__18353),
            .I(N__18350));
    InMux I__1887 (
            .O(N__18350),
            .I(N__18347));
    LocalMux I__1886 (
            .O(N__18347),
            .I(n317));
    CascadeMux I__1885 (
            .O(N__18344),
            .I(N__18341));
    InMux I__1884 (
            .O(N__18341),
            .I(N__18338));
    LocalMux I__1883 (
            .O(N__18338),
            .I(n318));
    CascadeMux I__1882 (
            .O(N__18335),
            .I(N__18332));
    InMux I__1881 (
            .O(N__18332),
            .I(N__18329));
    LocalMux I__1880 (
            .O(N__18329),
            .I(N__18326));
    Odrv4 I__1879 (
            .O(N__18326),
            .I(n319));
    CascadeMux I__1878 (
            .O(N__18323),
            .I(N__18320));
    InMux I__1877 (
            .O(N__18320),
            .I(N__18317));
    LocalMux I__1876 (
            .O(N__18317),
            .I(n321));
    InMux I__1875 (
            .O(N__18314),
            .I(N__18311));
    LocalMux I__1874 (
            .O(N__18311),
            .I(N__18307));
    InMux I__1873 (
            .O(N__18310),
            .I(N__18304));
    Span4Mux_v I__1872 (
            .O(N__18307),
            .I(N__18301));
    LocalMux I__1871 (
            .O(N__18304),
            .I(data_out_frame2_5_0));
    Odrv4 I__1870 (
            .O(N__18301),
            .I(data_out_frame2_5_0));
    CascadeMux I__1869 (
            .O(N__18296),
            .I(\c0.n5_adj_2477_cascade_ ));
    InMux I__1868 (
            .O(N__18293),
            .I(N__18290));
    LocalMux I__1867 (
            .O(N__18290),
            .I(N__18287));
    Odrv4 I__1866 (
            .O(N__18287),
            .I(\c0.n6_adj_2436 ));
    InMux I__1865 (
            .O(N__18284),
            .I(N__18280));
    InMux I__1864 (
            .O(N__18283),
            .I(N__18277));
    LocalMux I__1863 (
            .O(N__18280),
            .I(N__18274));
    LocalMux I__1862 (
            .O(N__18277),
            .I(data_out_frame2_18_1));
    Odrv4 I__1861 (
            .O(N__18274),
            .I(data_out_frame2_18_1));
    InMux I__1860 (
            .O(N__18269),
            .I(N__18266));
    LocalMux I__1859 (
            .O(N__18266),
            .I(\c0.n18468 ));
    InMux I__1858 (
            .O(N__18263),
            .I(N__18259));
    InMux I__1857 (
            .O(N__18262),
            .I(N__18256));
    LocalMux I__1856 (
            .O(N__18259),
            .I(data_out_frame2_5_1));
    LocalMux I__1855 (
            .O(N__18256),
            .I(data_out_frame2_5_1));
    InMux I__1854 (
            .O(N__18251),
            .I(N__18247));
    InMux I__1853 (
            .O(N__18250),
            .I(N__18244));
    LocalMux I__1852 (
            .O(N__18247),
            .I(N__18241));
    LocalMux I__1851 (
            .O(N__18244),
            .I(data_out_frame2_10_2));
    Odrv4 I__1850 (
            .O(N__18241),
            .I(data_out_frame2_10_2));
    CascadeMux I__1849 (
            .O(N__18236),
            .I(N__18233));
    InMux I__1848 (
            .O(N__18233),
            .I(N__18230));
    LocalMux I__1847 (
            .O(N__18230),
            .I(N__18227));
    Span4Mux_h I__1846 (
            .O(N__18227),
            .I(N__18223));
    InMux I__1845 (
            .O(N__18226),
            .I(N__18220));
    Span4Mux_v I__1844 (
            .O(N__18223),
            .I(N__18217));
    LocalMux I__1843 (
            .O(N__18220),
            .I(data_out_frame2_11_2));
    Odrv4 I__1842 (
            .O(N__18217),
            .I(data_out_frame2_11_2));
    InMux I__1841 (
            .O(N__18212),
            .I(N__18208));
    InMux I__1840 (
            .O(N__18211),
            .I(N__18205));
    LocalMux I__1839 (
            .O(N__18208),
            .I(data_out_frame2_12_0));
    LocalMux I__1838 (
            .O(N__18205),
            .I(data_out_frame2_12_0));
    InMux I__1837 (
            .O(N__18200),
            .I(N__18197));
    LocalMux I__1836 (
            .O(N__18197),
            .I(N__18194));
    Odrv12 I__1835 (
            .O(N__18194),
            .I(\c0.n17794 ));
    InMux I__1834 (
            .O(N__18191),
            .I(N__18188));
    LocalMux I__1833 (
            .O(N__18188),
            .I(N__18185));
    Span4Mux_h I__1832 (
            .O(N__18185),
            .I(N__18182));
    Span4Mux_v I__1831 (
            .O(N__18182),
            .I(N__18179));
    Odrv4 I__1830 (
            .O(N__18179),
            .I(\c0.n18078 ));
    CascadeMux I__1829 (
            .O(N__18176),
            .I(\c0.n18408_cascade_ ));
    InMux I__1828 (
            .O(N__18173),
            .I(N__18170));
    LocalMux I__1827 (
            .O(N__18170),
            .I(N__18167));
    Span12Mux_v I__1826 (
            .O(N__18167),
            .I(N__18164));
    Odrv12 I__1825 (
            .O(N__18164),
            .I(\c0.n6_adj_2506 ));
    InMux I__1824 (
            .O(N__18161),
            .I(N__18158));
    LocalMux I__1823 (
            .O(N__18158),
            .I(\c0.n5_adj_2495 ));
    CascadeMux I__1822 (
            .O(N__18155),
            .I(N__18152));
    InMux I__1821 (
            .O(N__18152),
            .I(N__18149));
    LocalMux I__1820 (
            .O(N__18149),
            .I(N__18145));
    InMux I__1819 (
            .O(N__18148),
            .I(N__18142));
    Span4Mux_v I__1818 (
            .O(N__18145),
            .I(N__18139));
    LocalMux I__1817 (
            .O(N__18142),
            .I(data_out_frame2_5_5));
    Odrv4 I__1816 (
            .O(N__18139),
            .I(data_out_frame2_5_5));
    InMux I__1815 (
            .O(N__18134),
            .I(N__18131));
    LocalMux I__1814 (
            .O(N__18131),
            .I(N__18128));
    Span4Mux_s1_h I__1813 (
            .O(N__18128),
            .I(N__18125));
    Odrv4 I__1812 (
            .O(N__18125),
            .I(\c0.n6_adj_2496 ));
    CascadeMux I__1811 (
            .O(N__18122),
            .I(N__18118));
    InMux I__1810 (
            .O(N__18121),
            .I(N__18115));
    InMux I__1809 (
            .O(N__18118),
            .I(N__18112));
    LocalMux I__1808 (
            .O(N__18115),
            .I(data_out_frame2_11_3));
    LocalMux I__1807 (
            .O(N__18112),
            .I(data_out_frame2_11_3));
    InMux I__1806 (
            .O(N__18107),
            .I(N__18104));
    LocalMux I__1805 (
            .O(N__18104),
            .I(N__18101));
    Odrv12 I__1804 (
            .O(N__18101),
            .I(\c0.n17629 ));
    InMux I__1803 (
            .O(N__18098),
            .I(N__18095));
    LocalMux I__1802 (
            .O(N__18095),
            .I(N__18092));
    Span4Mux_h I__1801 (
            .O(N__18092),
            .I(N__18089));
    Span4Mux_v I__1800 (
            .O(N__18089),
            .I(N__18086));
    Span4Mux_v I__1799 (
            .O(N__18086),
            .I(N__18083));
    Odrv4 I__1798 (
            .O(N__18083),
            .I(\c0.n8725 ));
    InMux I__1797 (
            .O(N__18080),
            .I(N__18076));
    InMux I__1796 (
            .O(N__18079),
            .I(N__18073));
    LocalMux I__1795 (
            .O(N__18076),
            .I(data_out_frame2_10_0));
    LocalMux I__1794 (
            .O(N__18073),
            .I(data_out_frame2_10_0));
    InMux I__1793 (
            .O(N__18068),
            .I(N__18065));
    LocalMux I__1792 (
            .O(N__18065),
            .I(N__18061));
    InMux I__1791 (
            .O(N__18064),
            .I(N__18058));
    Span4Mux_v I__1790 (
            .O(N__18061),
            .I(N__18055));
    LocalMux I__1789 (
            .O(N__18058),
            .I(data_out_frame2_17_0));
    Odrv4 I__1788 (
            .O(N__18055),
            .I(data_out_frame2_17_0));
    CascadeMux I__1787 (
            .O(N__18050),
            .I(N__18047));
    InMux I__1786 (
            .O(N__18047),
            .I(N__18043));
    InMux I__1785 (
            .O(N__18046),
            .I(N__18040));
    LocalMux I__1784 (
            .O(N__18043),
            .I(N__18037));
    LocalMux I__1783 (
            .O(N__18040),
            .I(data_out_frame2_16_0));
    Odrv4 I__1782 (
            .O(N__18037),
            .I(data_out_frame2_16_0));
    InMux I__1781 (
            .O(N__18032),
            .I(N__18029));
    LocalMux I__1780 (
            .O(N__18029),
            .I(\c0.n18600 ));
    CascadeMux I__1779 (
            .O(N__18026),
            .I(N__18022));
    InMux I__1778 (
            .O(N__18025),
            .I(N__18017));
    InMux I__1777 (
            .O(N__18022),
            .I(N__18017));
    LocalMux I__1776 (
            .O(N__18017),
            .I(data_out_frame2_8_6));
    InMux I__1775 (
            .O(N__18014),
            .I(N__18011));
    LocalMux I__1774 (
            .O(N__18011),
            .I(N__18008));
    Span12Mux_s7_v I__1773 (
            .O(N__18008),
            .I(N__18005));
    Odrv12 I__1772 (
            .O(N__18005),
            .I(\c0.n18564 ));
    CascadeMux I__1771 (
            .O(N__18002),
            .I(N__17999));
    InMux I__1770 (
            .O(N__17999),
            .I(N__17995));
    InMux I__1769 (
            .O(N__17998),
            .I(N__17992));
    LocalMux I__1768 (
            .O(N__17995),
            .I(N__17989));
    LocalMux I__1767 (
            .O(N__17992),
            .I(N__17984));
    Span4Mux_v I__1766 (
            .O(N__17989),
            .I(N__17984));
    Odrv4 I__1765 (
            .O(N__17984),
            .I(data_out_frame2_16_1));
    InMux I__1764 (
            .O(N__17981),
            .I(N__17978));
    LocalMux I__1763 (
            .O(N__17978),
            .I(N__17974));
    InMux I__1762 (
            .O(N__17977),
            .I(N__17971));
    Span4Mux_s1_h I__1761 (
            .O(N__17974),
            .I(N__17968));
    LocalMux I__1760 (
            .O(N__17971),
            .I(data_out_frame2_17_1));
    Odrv4 I__1759 (
            .O(N__17968),
            .I(data_out_frame2_17_1));
    InMux I__1758 (
            .O(N__17963),
            .I(N__17959));
    InMux I__1757 (
            .O(N__17962),
            .I(N__17956));
    LocalMux I__1756 (
            .O(N__17959),
            .I(data_out_frame2_18_0));
    LocalMux I__1755 (
            .O(N__17956),
            .I(data_out_frame2_18_0));
    InMux I__1754 (
            .O(N__17951),
            .I(N__17947));
    InMux I__1753 (
            .O(N__17950),
            .I(N__17944));
    LocalMux I__1752 (
            .O(N__17947),
            .I(data_out_frame2_10_3));
    LocalMux I__1751 (
            .O(N__17944),
            .I(data_out_frame2_10_3));
    InMux I__1750 (
            .O(N__17939),
            .I(N__17935));
    InMux I__1749 (
            .O(N__17938),
            .I(N__17932));
    LocalMux I__1748 (
            .O(N__17935),
            .I(data_out_frame2_14_4));
    LocalMux I__1747 (
            .O(N__17932),
            .I(data_out_frame2_14_4));
    InMux I__1746 (
            .O(N__17927),
            .I(N__17924));
    LocalMux I__1745 (
            .O(N__17924),
            .I(N__17921));
    Span4Mux_h I__1744 (
            .O(N__17921),
            .I(N__17917));
    InMux I__1743 (
            .O(N__17920),
            .I(N__17914));
    Span4Mux_v I__1742 (
            .O(N__17917),
            .I(N__17911));
    LocalMux I__1741 (
            .O(N__17914),
            .I(data_out_frame2_7_6));
    Odrv4 I__1740 (
            .O(N__17911),
            .I(data_out_frame2_7_6));
    InMux I__1739 (
            .O(N__17906),
            .I(N__17902));
    InMux I__1738 (
            .O(N__17905),
            .I(N__17899));
    LocalMux I__1737 (
            .O(N__17902),
            .I(data_out_frame2_8_5));
    LocalMux I__1736 (
            .O(N__17899),
            .I(data_out_frame2_8_5));
    InMux I__1735 (
            .O(N__17894),
            .I(N__17890));
    InMux I__1734 (
            .O(N__17893),
            .I(N__17887));
    LocalMux I__1733 (
            .O(N__17890),
            .I(N__17884));
    LocalMux I__1732 (
            .O(N__17887),
            .I(data_out_frame2_15_1));
    Odrv4 I__1731 (
            .O(N__17884),
            .I(data_out_frame2_15_1));
    CascadeMux I__1730 (
            .O(N__17879),
            .I(N__17876));
    InMux I__1729 (
            .O(N__17876),
            .I(N__17872));
    InMux I__1728 (
            .O(N__17875),
            .I(N__17869));
    LocalMux I__1727 (
            .O(N__17872),
            .I(N__17866));
    LocalMux I__1726 (
            .O(N__17869),
            .I(data_out_frame2_11_6));
    Odrv12 I__1725 (
            .O(N__17866),
            .I(data_out_frame2_11_6));
    InMux I__1724 (
            .O(N__17861),
            .I(N__17857));
    InMux I__1723 (
            .O(N__17860),
            .I(N__17854));
    LocalMux I__1722 (
            .O(N__17857),
            .I(N__17851));
    LocalMux I__1721 (
            .O(N__17854),
            .I(data_out_frame2_15_6));
    Odrv12 I__1720 (
            .O(N__17851),
            .I(data_out_frame2_15_6));
    CascadeMux I__1719 (
            .O(N__17846),
            .I(N__17843));
    InMux I__1718 (
            .O(N__17843),
            .I(N__17839));
    InMux I__1717 (
            .O(N__17842),
            .I(N__17836));
    LocalMux I__1716 (
            .O(N__17839),
            .I(N__17833));
    LocalMux I__1715 (
            .O(N__17836),
            .I(data_out_frame2_5_2));
    Odrv4 I__1714 (
            .O(N__17833),
            .I(data_out_frame2_5_2));
    CascadeMux I__1713 (
            .O(N__17828),
            .I(N__17825));
    InMux I__1712 (
            .O(N__17825),
            .I(N__17821));
    InMux I__1711 (
            .O(N__17824),
            .I(N__17818));
    LocalMux I__1710 (
            .O(N__17821),
            .I(N__17815));
    LocalMux I__1709 (
            .O(N__17818),
            .I(data_out_frame2_15_2));
    Odrv4 I__1708 (
            .O(N__17815),
            .I(data_out_frame2_15_2));
    CascadeMux I__1707 (
            .O(N__17810),
            .I(N__17807));
    InMux I__1706 (
            .O(N__17807),
            .I(N__17803));
    InMux I__1705 (
            .O(N__17806),
            .I(N__17800));
    LocalMux I__1704 (
            .O(N__17803),
            .I(N__17797));
    LocalMux I__1703 (
            .O(N__17800),
            .I(data_out_frame2_15_0));
    Odrv4 I__1702 (
            .O(N__17797),
            .I(data_out_frame2_15_0));
    CascadeMux I__1701 (
            .O(N__17792),
            .I(N__17789));
    InMux I__1700 (
            .O(N__17789),
            .I(N__17783));
    InMux I__1699 (
            .O(N__17788),
            .I(N__17783));
    LocalMux I__1698 (
            .O(N__17783),
            .I(data_out_frame2_13_2));
    InMux I__1697 (
            .O(N__17780),
            .I(N__17777));
    LocalMux I__1696 (
            .O(N__17777),
            .I(N__17774));
    Span4Mux_h I__1695 (
            .O(N__17774),
            .I(N__17771));
    Odrv4 I__1694 (
            .O(N__17771),
            .I(\c0.n18492 ));
    InMux I__1693 (
            .O(N__17768),
            .I(N__17765));
    LocalMux I__1692 (
            .O(N__17765),
            .I(N__17762));
    Odrv4 I__1691 (
            .O(N__17762),
            .I(\c0.n17827 ));
    InMux I__1690 (
            .O(N__17759),
            .I(N__17753));
    InMux I__1689 (
            .O(N__17758),
            .I(N__17753));
    LocalMux I__1688 (
            .O(N__17753),
            .I(data_out_frame2_12_5));
    CascadeMux I__1687 (
            .O(N__17750),
            .I(\c0.n9043_cascade_ ));
    InMux I__1686 (
            .O(N__17747),
            .I(N__17744));
    LocalMux I__1685 (
            .O(N__17744),
            .I(N__17740));
    InMux I__1684 (
            .O(N__17743),
            .I(N__17737));
    Span12Mux_v I__1683 (
            .O(N__17740),
            .I(N__17734));
    LocalMux I__1682 (
            .O(N__17737),
            .I(data_out_frame2_14_6));
    Odrv12 I__1681 (
            .O(N__17734),
            .I(data_out_frame2_14_6));
    InMux I__1680 (
            .O(N__17729),
            .I(N__17726));
    LocalMux I__1679 (
            .O(N__17726),
            .I(N__17722));
    InMux I__1678 (
            .O(N__17725),
            .I(N__17719));
    Sp12to4 I__1677 (
            .O(N__17722),
            .I(N__17716));
    LocalMux I__1676 (
            .O(N__17719),
            .I(data_out_frame2_10_6));
    Odrv12 I__1675 (
            .O(N__17716),
            .I(data_out_frame2_10_6));
    CascadeMux I__1674 (
            .O(N__17711),
            .I(N__17708));
    InMux I__1673 (
            .O(N__17708),
            .I(N__17705));
    LocalMux I__1672 (
            .O(N__17705),
            .I(N__17701));
    InMux I__1671 (
            .O(N__17704),
            .I(N__17698));
    Span4Mux_v I__1670 (
            .O(N__17701),
            .I(N__17695));
    LocalMux I__1669 (
            .O(N__17698),
            .I(data_out_frame2_11_0));
    Odrv4 I__1668 (
            .O(N__17695),
            .I(data_out_frame2_11_0));
    InMux I__1667 (
            .O(N__17690),
            .I(N__17687));
    LocalMux I__1666 (
            .O(N__17687),
            .I(N__17684));
    Span4Mux_v I__1665 (
            .O(N__17684),
            .I(N__17681));
    Span4Mux_v I__1664 (
            .O(N__17681),
            .I(N__17677));
    InMux I__1663 (
            .O(N__17680),
            .I(N__17674));
    Span4Mux_v I__1662 (
            .O(N__17677),
            .I(N__17671));
    LocalMux I__1661 (
            .O(N__17674),
            .I(data_out_frame2_6_6));
    Odrv4 I__1660 (
            .O(N__17671),
            .I(data_out_frame2_6_6));
    InMux I__1659 (
            .O(N__17666),
            .I(N__17663));
    LocalMux I__1658 (
            .O(N__17663),
            .I(N__17660));
    Odrv12 I__1657 (
            .O(N__17660),
            .I(\c0.n9_adj_2507 ));
    CascadeMux I__1656 (
            .O(N__17657),
            .I(\c0.n17325_cascade_ ));
    CascadeMux I__1655 (
            .O(N__17654),
            .I(\c0.n8_adj_2459_cascade_ ));
    InMux I__1654 (
            .O(N__17651),
            .I(N__17648));
    LocalMux I__1653 (
            .O(N__17648),
            .I(\c0.n2604 ));
    InMux I__1652 (
            .O(N__17645),
            .I(N__17642));
    LocalMux I__1651 (
            .O(N__17642),
            .I(\c0.n11_adj_2460 ));
    CEMux I__1650 (
            .O(N__17639),
            .I(N__17636));
    LocalMux I__1649 (
            .O(N__17636),
            .I(N__17633));
    Span4Mux_s2_h I__1648 (
            .O(N__17633),
            .I(N__17630));
    Odrv4 I__1647 (
            .O(N__17630),
            .I(\c0.n9605 ));
    SRMux I__1646 (
            .O(N__17627),
            .I(N__17624));
    LocalMux I__1645 (
            .O(N__17624),
            .I(\c0.n9900 ));
    InMux I__1644 (
            .O(N__17621),
            .I(N__17618));
    LocalMux I__1643 (
            .O(N__17618),
            .I(\c0.n17806 ));
    InMux I__1642 (
            .O(N__17615),
            .I(N__17611));
    InMux I__1641 (
            .O(N__17614),
            .I(N__17608));
    LocalMux I__1640 (
            .O(N__17611),
            .I(data_out_frame2_18_5));
    LocalMux I__1639 (
            .O(N__17608),
            .I(data_out_frame2_18_5));
    InMux I__1638 (
            .O(N__17603),
            .I(N__17600));
    LocalMux I__1637 (
            .O(N__17600),
            .I(\c0.n2607 ));
    CascadeMux I__1636 (
            .O(N__17597),
            .I(N__17594));
    InMux I__1635 (
            .O(N__17594),
            .I(N__17591));
    LocalMux I__1634 (
            .O(N__17591),
            .I(\c0.n17513 ));
    InMux I__1633 (
            .O(N__17588),
            .I(N__17585));
    LocalMux I__1632 (
            .O(N__17585),
            .I(\c0.n2602 ));
    CascadeMux I__1631 (
            .O(N__17582),
            .I(N__17579));
    InMux I__1630 (
            .O(N__17579),
            .I(N__17569));
    InMux I__1629 (
            .O(N__17578),
            .I(N__17569));
    InMux I__1628 (
            .O(N__17577),
            .I(N__17569));
    InMux I__1627 (
            .O(N__17576),
            .I(N__17566));
    LocalMux I__1626 (
            .O(N__17569),
            .I(N__17563));
    LocalMux I__1625 (
            .O(N__17566),
            .I(\c0.data_in_frame_3_2 ));
    Odrv4 I__1624 (
            .O(N__17563),
            .I(\c0.data_in_frame_3_2 ));
    CascadeMux I__1623 (
            .O(N__17558),
            .I(N__17555));
    InMux I__1622 (
            .O(N__17555),
            .I(N__17552));
    LocalMux I__1621 (
            .O(N__17552),
            .I(\c0.n9_adj_2500 ));
    InMux I__1620 (
            .O(N__17549),
            .I(N__17545));
    InMux I__1619 (
            .O(N__17548),
            .I(N__17542));
    LocalMux I__1618 (
            .O(N__17545),
            .I(\c0.data_out_frame2_0_5 ));
    LocalMux I__1617 (
            .O(N__17542),
            .I(\c0.data_out_frame2_0_5 ));
    CascadeMux I__1616 (
            .O(N__17537),
            .I(N__17533));
    CascadeMux I__1615 (
            .O(N__17536),
            .I(N__17530));
    InMux I__1614 (
            .O(N__17533),
            .I(N__17527));
    InMux I__1613 (
            .O(N__17530),
            .I(N__17524));
    LocalMux I__1612 (
            .O(N__17527),
            .I(\c0.data_in_frame_3_3 ));
    LocalMux I__1611 (
            .O(N__17524),
            .I(\c0.data_in_frame_3_3 ));
    CascadeMux I__1610 (
            .O(N__17519),
            .I(\c0.n17629_cascade_ ));
    InMux I__1609 (
            .O(N__17516),
            .I(N__17513));
    LocalMux I__1608 (
            .O(N__17513),
            .I(\c0.n16_adj_2546 ));
    InMux I__1607 (
            .O(N__17510),
            .I(N__17507));
    LocalMux I__1606 (
            .O(N__17507),
            .I(\c0.n9254 ));
    CascadeMux I__1605 (
            .O(N__17504),
            .I(\c0.n9254_cascade_ ));
    InMux I__1604 (
            .O(N__17501),
            .I(N__17495));
    InMux I__1603 (
            .O(N__17500),
            .I(N__17489));
    InMux I__1602 (
            .O(N__17499),
            .I(N__17489));
    InMux I__1601 (
            .O(N__17498),
            .I(N__17486));
    LocalMux I__1600 (
            .O(N__17495),
            .I(N__17483));
    InMux I__1599 (
            .O(N__17494),
            .I(N__17480));
    LocalMux I__1598 (
            .O(N__17489),
            .I(\c0.data_in_frame_2_5 ));
    LocalMux I__1597 (
            .O(N__17486),
            .I(\c0.data_in_frame_2_5 ));
    Odrv4 I__1596 (
            .O(N__17483),
            .I(\c0.data_in_frame_2_5 ));
    LocalMux I__1595 (
            .O(N__17480),
            .I(\c0.data_in_frame_2_5 ));
    InMux I__1594 (
            .O(N__17471),
            .I(N__17467));
    InMux I__1593 (
            .O(N__17470),
            .I(N__17464));
    LocalMux I__1592 (
            .O(N__17467),
            .I(\c0.n8976 ));
    LocalMux I__1591 (
            .O(N__17464),
            .I(\c0.n8976 ));
    CascadeMux I__1590 (
            .O(N__17459),
            .I(N__17456));
    InMux I__1589 (
            .O(N__17456),
            .I(N__17453));
    LocalMux I__1588 (
            .O(N__17453),
            .I(N__17448));
    InMux I__1587 (
            .O(N__17452),
            .I(N__17443));
    InMux I__1586 (
            .O(N__17451),
            .I(N__17443));
    Odrv12 I__1585 (
            .O(N__17448),
            .I(\c0.data_in_frame_1_3 ));
    LocalMux I__1584 (
            .O(N__17443),
            .I(\c0.data_in_frame_1_3 ));
    CascadeMux I__1583 (
            .O(N__17438),
            .I(N__17435));
    InMux I__1582 (
            .O(N__17435),
            .I(N__17432));
    LocalMux I__1581 (
            .O(N__17432),
            .I(N__17429));
    Span4Mux_v I__1580 (
            .O(N__17429),
            .I(N__17426));
    Odrv4 I__1579 (
            .O(N__17426),
            .I(\c0.n5_adj_2515 ));
    InMux I__1578 (
            .O(N__17423),
            .I(N__17420));
    LocalMux I__1577 (
            .O(N__17420),
            .I(\c0.n17507 ));
    CascadeMux I__1576 (
            .O(N__17417),
            .I(\c0.n17476_cascade_ ));
    InMux I__1575 (
            .O(N__17414),
            .I(N__17411));
    LocalMux I__1574 (
            .O(N__17411),
            .I(\c0.n17476 ));
    CascadeMux I__1573 (
            .O(N__17408),
            .I(\c0.n17478_cascade_ ));
    InMux I__1572 (
            .O(N__17405),
            .I(N__17402));
    LocalMux I__1571 (
            .O(N__17402),
            .I(n316));
    CascadeMux I__1570 (
            .O(N__17399),
            .I(\c0.n17507_cascade_ ));
    CascadeMux I__1569 (
            .O(N__17396),
            .I(N__17393));
    InMux I__1568 (
            .O(N__17393),
            .I(N__17385));
    InMux I__1567 (
            .O(N__17392),
            .I(N__17385));
    InMux I__1566 (
            .O(N__17391),
            .I(N__17382));
    InMux I__1565 (
            .O(N__17390),
            .I(N__17379));
    LocalMux I__1564 (
            .O(N__17385),
            .I(\c0.data_in_frame_0_4 ));
    LocalMux I__1563 (
            .O(N__17382),
            .I(\c0.data_in_frame_0_4 ));
    LocalMux I__1562 (
            .O(N__17379),
            .I(\c0.data_in_frame_0_4 ));
    InMux I__1561 (
            .O(N__17372),
            .I(\c0.tx2.n16374 ));
    InMux I__1560 (
            .O(N__17369),
            .I(\c0.tx2.n16375 ));
    InMux I__1559 (
            .O(N__17366),
            .I(\c0.tx2.n16376 ));
    InMux I__1558 (
            .O(N__17363),
            .I(\c0.tx2.n16377 ));
    InMux I__1557 (
            .O(N__17360),
            .I(\c0.tx2.n16378 ));
    InMux I__1556 (
            .O(N__17357),
            .I(bfn_1_32_0_));
    InMux I__1555 (
            .O(N__17354),
            .I(N__17351));
    LocalMux I__1554 (
            .O(N__17351),
            .I(\c0.tx2.n17953 ));
    InMux I__1553 (
            .O(N__17348),
            .I(N__17345));
    LocalMux I__1552 (
            .O(N__17345),
            .I(\c0.tx2.n18013 ));
    InMux I__1551 (
            .O(N__17342),
            .I(N__17339));
    LocalMux I__1550 (
            .O(N__17339),
            .I(\c0.tx2.n17939 ));
    CascadeMux I__1549 (
            .O(N__17336),
            .I(\c0.n18435_cascade_ ));
    CascadeMux I__1548 (
            .O(N__17333),
            .I(N__17330));
    InMux I__1547 (
            .O(N__17330),
            .I(N__17327));
    LocalMux I__1546 (
            .O(N__17327),
            .I(N__17324));
    Span12Mux_s3_v I__1545 (
            .O(N__17324),
            .I(N__17321));
    Odrv12 I__1544 (
            .O(N__17321),
            .I(\c0.n17836 ));
    CascadeMux I__1543 (
            .O(N__17318),
            .I(\c0.n18360_cascade_ ));
    InMux I__1542 (
            .O(N__17315),
            .I(N__17312));
    LocalMux I__1541 (
            .O(N__17312),
            .I(N__17309));
    Odrv4 I__1540 (
            .O(N__17309),
            .I(\c0.n6_adj_2504 ));
    CascadeMux I__1539 (
            .O(N__17306),
            .I(\c0.n18471_cascade_ ));
    InMux I__1538 (
            .O(N__17303),
            .I(N__17300));
    LocalMux I__1537 (
            .O(N__17300),
            .I(\c0.n18363 ));
    CascadeMux I__1536 (
            .O(N__17297),
            .I(\c0.n22_adj_2530_cascade_ ));
    InMux I__1535 (
            .O(N__17294),
            .I(bfn_1_31_0_));
    InMux I__1534 (
            .O(N__17291),
            .I(\c0.tx2.n16372 ));
    InMux I__1533 (
            .O(N__17288),
            .I(\c0.tx2.n16373 ));
    CascadeMux I__1532 (
            .O(N__17285),
            .I(\c0.n5_adj_2503_cascade_ ));
    InMux I__1531 (
            .O(N__17282),
            .I(N__17276));
    InMux I__1530 (
            .O(N__17281),
            .I(N__17276));
    LocalMux I__1529 (
            .O(N__17276),
            .I(data_out_frame2_14_2));
    CascadeMux I__1528 (
            .O(N__17273),
            .I(\c0.n18606_cascade_ ));
    CascadeMux I__1527 (
            .O(N__17270),
            .I(\c0.n18570_cascade_ ));
    InMux I__1526 (
            .O(N__17267),
            .I(N__17264));
    LocalMux I__1525 (
            .O(N__17264),
            .I(\c0.n17779 ));
    CascadeMux I__1524 (
            .O(N__17261),
            .I(\c0.n17773_cascade_ ));
    InMux I__1523 (
            .O(N__17258),
            .I(N__17255));
    LocalMux I__1522 (
            .O(N__17255),
            .I(N__17252));
    Odrv12 I__1521 (
            .O(N__17252),
            .I(\c0.n18074 ));
    CascadeMux I__1520 (
            .O(N__17249),
            .I(\c0.n18432_cascade_ ));
    InMux I__1519 (
            .O(N__17246),
            .I(N__17242));
    InMux I__1518 (
            .O(N__17245),
            .I(N__17239));
    LocalMux I__1517 (
            .O(N__17242),
            .I(N__17236));
    LocalMux I__1516 (
            .O(N__17239),
            .I(data_out_frame2_16_2));
    Odrv12 I__1515 (
            .O(N__17236),
            .I(data_out_frame2_16_2));
    CascadeMux I__1514 (
            .O(N__17231),
            .I(\c0.n18486_cascade_ ));
    CascadeMux I__1513 (
            .O(N__17228),
            .I(\c0.n18489_cascade_ ));
    InMux I__1512 (
            .O(N__17225),
            .I(N__17222));
    LocalMux I__1511 (
            .O(N__17222),
            .I(\c0.n18084 ));
    CascadeMux I__1510 (
            .O(N__17219),
            .I(\c0.n18366_cascade_ ));
    InMux I__1509 (
            .O(N__17216),
            .I(N__17213));
    LocalMux I__1508 (
            .O(N__17213),
            .I(N__17210));
    Odrv4 I__1507 (
            .O(N__17210),
            .I(\c0.n6_adj_2466 ));
    InMux I__1506 (
            .O(N__17207),
            .I(N__17204));
    LocalMux I__1505 (
            .O(N__17204),
            .I(\c0.n22_adj_2529 ));
    CascadeMux I__1504 (
            .O(N__17201),
            .I(\c0.n18369_cascade_ ));
    InMux I__1503 (
            .O(N__17198),
            .I(N__17194));
    InMux I__1502 (
            .O(N__17197),
            .I(N__17191));
    LocalMux I__1501 (
            .O(N__17194),
            .I(N__17188));
    LocalMux I__1500 (
            .O(N__17191),
            .I(data_out_frame2_7_5));
    Odrv4 I__1499 (
            .O(N__17188),
            .I(data_out_frame2_7_5));
    CascadeMux I__1498 (
            .O(N__17183),
            .I(\c0.n18387_cascade_ ));
    InMux I__1497 (
            .O(N__17180),
            .I(N__17177));
    LocalMux I__1496 (
            .O(N__17177),
            .I(N__17174));
    Odrv4 I__1495 (
            .O(N__17174),
            .I(\c0.n5_adj_2463 ));
    InMux I__1494 (
            .O(N__17171),
            .I(N__17167));
    InMux I__1493 (
            .O(N__17170),
            .I(N__17164));
    LocalMux I__1492 (
            .O(N__17167),
            .I(data_out_frame2_16_5));
    LocalMux I__1491 (
            .O(N__17164),
            .I(data_out_frame2_16_5));
    InMux I__1490 (
            .O(N__17159),
            .I(N__17155));
    InMux I__1489 (
            .O(N__17158),
            .I(N__17152));
    LocalMux I__1488 (
            .O(N__17155),
            .I(N__17149));
    LocalMux I__1487 (
            .O(N__17152),
            .I(data_out_frame2_9_5));
    Odrv4 I__1486 (
            .O(N__17149),
            .I(data_out_frame2_9_5));
    InMux I__1485 (
            .O(N__17144),
            .I(N__17141));
    LocalMux I__1484 (
            .O(N__17141),
            .I(N__17137));
    InMux I__1483 (
            .O(N__17140),
            .I(N__17134));
    Span4Mux_s1_h I__1482 (
            .O(N__17137),
            .I(N__17131));
    LocalMux I__1481 (
            .O(N__17134),
            .I(data_out_frame2_6_2));
    Odrv4 I__1480 (
            .O(N__17131),
            .I(data_out_frame2_6_2));
    InMux I__1479 (
            .O(N__17126),
            .I(N__17123));
    LocalMux I__1478 (
            .O(N__17123),
            .I(\c0.n18474 ));
    CascadeMux I__1477 (
            .O(N__17120),
            .I(\c0.n18534_cascade_ ));
    InMux I__1476 (
            .O(N__17117),
            .I(N__17113));
    InMux I__1475 (
            .O(N__17116),
            .I(N__17110));
    LocalMux I__1474 (
            .O(N__17113),
            .I(data_out_frame2_17_5));
    LocalMux I__1473 (
            .O(N__17110),
            .I(data_out_frame2_17_5));
    CascadeMux I__1472 (
            .O(N__17105),
            .I(\c0.n18537_cascade_ ));
    InMux I__1471 (
            .O(N__17102),
            .I(N__17099));
    LocalMux I__1470 (
            .O(N__17099),
            .I(\c0.n17803 ));
    InMux I__1469 (
            .O(N__17096),
            .I(N__17093));
    LocalMux I__1468 (
            .O(N__17093),
            .I(N__17090));
    Odrv12 I__1467 (
            .O(N__17090),
            .I(\c0.n18080 ));
    CascadeMux I__1466 (
            .O(N__17087),
            .I(\c0.n18384_cascade_ ));
    InMux I__1465 (
            .O(N__17084),
            .I(N__17081));
    LocalMux I__1464 (
            .O(N__17081),
            .I(\c0.n22_adj_2523 ));
    InMux I__1463 (
            .O(N__17078),
            .I(N__17072));
    InMux I__1462 (
            .O(N__17077),
            .I(N__17072));
    LocalMux I__1461 (
            .O(N__17072),
            .I(\c0.data_out_frame2_0_0 ));
    InMux I__1460 (
            .O(N__17069),
            .I(N__17063));
    InMux I__1459 (
            .O(N__17068),
            .I(N__17063));
    LocalMux I__1458 (
            .O(N__17063),
            .I(data_out_frame2_7_2));
    InMux I__1457 (
            .O(N__17060),
            .I(N__17056));
    InMux I__1456 (
            .O(N__17059),
            .I(N__17053));
    LocalMux I__1455 (
            .O(N__17056),
            .I(N__17050));
    LocalMux I__1454 (
            .O(N__17053),
            .I(\c0.data_out_frame2_0_6 ));
    Odrv12 I__1453 (
            .O(N__17050),
            .I(\c0.data_out_frame2_0_6 ));
    CascadeMux I__1452 (
            .O(N__17045),
            .I(\c0.n18546_cascade_ ));
    CascadeMux I__1451 (
            .O(N__17042),
            .I(N__17038));
    InMux I__1450 (
            .O(N__17041),
            .I(N__17033));
    InMux I__1449 (
            .O(N__17038),
            .I(N__17033));
    LocalMux I__1448 (
            .O(N__17033),
            .I(data_out_frame2_11_5));
    InMux I__1447 (
            .O(N__17030),
            .I(\c0.n16405 ));
    InMux I__1446 (
            .O(N__17027),
            .I(\c0.n16406 ));
    InMux I__1445 (
            .O(N__17024),
            .I(\c0.n16407 ));
    InMux I__1444 (
            .O(N__17021),
            .I(\c0.n16408 ));
    InMux I__1443 (
            .O(N__17018),
            .I(\c0.n16409 ));
    InMux I__1442 (
            .O(N__17015),
            .I(\c0.n16410 ));
    InMux I__1441 (
            .O(N__17012),
            .I(\c0.n16411 ));
    CascadeMux I__1440 (
            .O(N__17009),
            .I(\c0.n20_adj_2547_cascade_ ));
    InMux I__1439 (
            .O(N__17006),
            .I(N__17003));
    LocalMux I__1438 (
            .O(N__17003),
            .I(N__16999));
    InMux I__1437 (
            .O(N__17002),
            .I(N__16996));
    Odrv4 I__1436 (
            .O(N__16999),
            .I(\c0.n9317 ));
    LocalMux I__1435 (
            .O(N__16996),
            .I(\c0.n9317 ));
    InMux I__1434 (
            .O(N__16991),
            .I(N__16988));
    LocalMux I__1433 (
            .O(N__16988),
            .I(\c0.n8063 ));
    InMux I__1432 (
            .O(N__16985),
            .I(N__16982));
    LocalMux I__1431 (
            .O(N__16982),
            .I(\c0.n17650 ));
    CascadeMux I__1430 (
            .O(N__16979),
            .I(\c0.n8645_cascade_ ));
    InMux I__1429 (
            .O(N__16976),
            .I(N__16973));
    LocalMux I__1428 (
            .O(N__16973),
            .I(N__16970));
    Odrv4 I__1427 (
            .O(N__16970),
            .I(\c0.n9186 ));
    CascadeMux I__1426 (
            .O(N__16967),
            .I(\c0.n30_adj_2489_cascade_ ));
    InMux I__1425 (
            .O(N__16964),
            .I(N__16961));
    LocalMux I__1424 (
            .O(N__16961),
            .I(\c0.n18_adj_2545 ));
    CascadeMux I__1423 (
            .O(N__16958),
            .I(\c0.n9186_cascade_ ));
    CascadeMux I__1422 (
            .O(N__16955),
            .I(\c0.n8857_cascade_ ));
    CascadeMux I__1421 (
            .O(N__16952),
            .I(\c0.n8725_cascade_ ));
    CascadeMux I__1420 (
            .O(N__16949),
            .I(\c0.n8063_cascade_ ));
    CascadeMux I__1419 (
            .O(N__16946),
            .I(N__16942));
    CascadeMux I__1418 (
            .O(N__16945),
            .I(N__16938));
    InMux I__1417 (
            .O(N__16942),
            .I(N__16928));
    InMux I__1416 (
            .O(N__16941),
            .I(N__16928));
    InMux I__1415 (
            .O(N__16938),
            .I(N__16928));
    InMux I__1414 (
            .O(N__16937),
            .I(N__16928));
    LocalMux I__1413 (
            .O(N__16928),
            .I(\c0.data_in_frame_0_3 ));
    IoInMux I__1412 (
            .O(N__16925),
            .I(N__16922));
    LocalMux I__1411 (
            .O(N__16922),
            .I(N__16919));
    IoSpan4Mux I__1410 (
            .O(N__16919),
            .I(N__16916));
    IoSpan4Mux I__1409 (
            .O(N__16916),
            .I(N__16913));
    IoSpan4Mux I__1408 (
            .O(N__16913),
            .I(N__16910));
    Odrv4 I__1407 (
            .O(N__16910),
            .I(CLK_pad_gb_input));
    defparam IN_MUX_bfv_9_29_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_29_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_29_0_));
    defparam IN_MUX_bfv_9_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_30_0_ (
            .carryinitin(n16419),
            .carryinitout(bfn_9_30_0_));
    defparam IN_MUX_bfv_9_31_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_31_0_ (
            .carryinitin(n16427),
            .carryinitout(bfn_9_31_0_));
    defparam IN_MUX_bfv_9_32_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_32_0_ (
            .carryinitin(n16435),
            .carryinitout(bfn_9_32_0_));
    defparam IN_MUX_bfv_5_29_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_29_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_29_0_));
    defparam IN_MUX_bfv_5_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_30_0_ (
            .carryinitin(n16326),
            .carryinitout(bfn_5_30_0_));
    defparam IN_MUX_bfv_5_31_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_31_0_ (
            .carryinitin(n16334),
            .carryinitout(bfn_5_31_0_));
    defparam IN_MUX_bfv_5_32_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_32_0_ (
            .carryinitin(n16342),
            .carryinitout(bfn_5_32_0_));
    defparam IN_MUX_bfv_1_31_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_31_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_31_0_));
    defparam IN_MUX_bfv_1_32_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_32_0_ (
            .carryinitin(\c0.tx2.n16379 ),
            .carryinitout(bfn_1_32_0_));
    defparam IN_MUX_bfv_5_25_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_25_0_));
    defparam IN_MUX_bfv_5_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_26_0_ (
            .carryinitin(\c0.tx.n16364 ),
            .carryinitout(bfn_5_26_0_));
    defparam IN_MUX_bfv_6_30_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_30_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_30_0_));
    defparam IN_MUX_bfv_1_22_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_22_0_));
    defparam IN_MUX_bfv_12_24_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_24_0_));
    defparam IN_MUX_bfv_12_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_25_0_ (
            .carryinitin(\c0.n16312 ),
            .carryinitout(bfn_12_25_0_));
    defparam IN_MUX_bfv_13_26_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_26_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_26_0_));
    defparam IN_MUX_bfv_16_29_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_29_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_29_0_));
    defparam IN_MUX_bfv_16_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_30_0_ (
            .carryinitin(n16387),
            .carryinitout(bfn_16_30_0_));
    defparam IN_MUX_bfv_16_31_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_31_0_ (
            .carryinitin(n16395),
            .carryinitout(bfn_16_31_0_));
    defparam IN_MUX_bfv_16_32_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_32_0_ (
            .carryinitin(n16403),
            .carryinitout(bfn_16_32_0_));
    ICE_GB CLK_pad_gb (
            .USERSIGNALTOGLOBALBUFFER(N__16925),
            .GLOBALBUFFEROUTPUT(CLK_c));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_998_LC_1_17_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_998_LC_1_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_998_LC_1_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_998_LC_1_17_0  (
            .in0(N__29030),
            .in1(N__21728),
            .in2(_gnd_net_),
            .in3(N__17501),
            .lcout(\c0.n17602 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_995_LC_1_17_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_995_LC_1_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_995_LC_1_17_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_995_LC_1_17_1  (
            .in0(N__29011),
            .in1(_gnd_net_),
            .in2(N__16945),
            .in3(N__22168),
            .lcout(\c0.n9163 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i15_LC_1_17_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i15_LC_1_17_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i15_LC_1_17_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i15_LC_1_17_2  (
            .in0(N__45511),
            .in1(N__27778),
            .in2(_gnd_net_),
            .in3(N__27719),
            .lcout(data_in_1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50251),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i33_LC_1_17_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i33_LC_1_17_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i33_LC_1_17_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_0___i33_LC_1_17_3  (
            .in0(N__22103),
            .in1(N__27850),
            .in2(_gnd_net_),
            .in3(N__45512),
            .lcout(data_in_4_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50251),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_945_LC_1_17_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_945_LC_1_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_945_LC_1_17_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_945_LC_1_17_4  (
            .in0(_gnd_net_),
            .in1(N__16937),
            .in2(_gnd_net_),
            .in3(N__29010),
            .lcout(\c0.n17550 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i4_LC_1_17_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i4_LC_1_17_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i4_LC_1_17_5 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \c0.data_in_frame_0___i4_LC_1_17_5  (
            .in0(N__27611),
            .in1(N__24272),
            .in2(N__16946),
            .in3(N__31976),
            .lcout(\c0.data_in_frame_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50251),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_987_LC_1_17_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_987_LC_1_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_987_LC_1_17_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_987_LC_1_17_6  (
            .in0(_gnd_net_),
            .in1(N__17392),
            .in2(_gnd_net_),
            .in3(N__16941),
            .lcout(\c0.n22_adj_2508 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i5_LC_1_17_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i5_LC_1_17_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i5_LC_1_17_7 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \c0.data_in_frame_0___i5_LC_1_17_7  (
            .in0(N__21629),
            .in1(N__24273),
            .in2(N__17396),
            .in3(N__31977),
            .lcout(\c0.data_in_frame_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50251),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i18_LC_1_18_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i18_LC_1_18_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i18_LC_1_18_1 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \c0.data_in_frame_0___i18_LC_1_18_1  (
            .in0(N__24271),
            .in1(N__31418),
            .in2(N__29040),
            .in3(N__31975),
            .lcout(\c0.data_in_frame_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50253),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_988_LC_1_18_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_988_LC_1_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_988_LC_1_18_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_988_LC_1_18_2  (
            .in0(_gnd_net_),
            .in1(N__29031),
            .in2(_gnd_net_),
            .in3(N__21718),
            .lcout(\c0.n9186 ),
            .ltout(\c0.n9186_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1015_LC_1_18_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1015_LC_1_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1015_LC_1_18_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1015_LC_1_18_3  (
            .in0(N__20556),
            .in1(N__18797),
            .in2(N__16958),
            .in3(N__18773),
            .lcout(\c0.n8857 ),
            .ltout(\c0.n8857_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_931_LC_1_18_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_931_LC_1_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_931_LC_1_18_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_931_LC_1_18_4  (
            .in0(N__20072),
            .in1(N__23022),
            .in2(N__16955),
            .in3(N__22229),
            .lcout(\c0.n17541 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_996_LC_1_18_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_996_LC_1_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_996_LC_1_18_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_996_LC_1_18_5  (
            .in0(N__20482),
            .in1(N__20071),
            .in2(N__25589),
            .in3(N__20425),
            .lcout(\c0.n8725 ),
            .ltout(\c0.n8725_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_864_LC_1_18_6 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_864_LC_1_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_864_LC_1_18_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_864_LC_1_18_6  (
            .in0(N__17510),
            .in1(N__25025),
            .in2(N__16952),
            .in3(N__17006),
            .lcout(\c0.n17594 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1024_LC_1_18_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1024_LC_1_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1024_LC_1_18_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1024_LC_1_18_7  (
            .in0(N__17494),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20424),
            .lcout(\c0.n9176 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_960_LC_1_19_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_960_LC_1_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_960_LC_1_19_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_960_LC_1_19_0  (
            .in0(N__22755),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24673),
            .lcout(\c0.n8063 ),
            .ltout(\c0.n8063_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_1115_LC_1_19_1 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_1115_LC_1_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_1115_LC_1_19_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_1115_LC_1_19_1  (
            .in0(N__16985),
            .in1(N__22450),
            .in2(N__16949),
            .in3(N__16964),
            .lcout(),
            .ltout(\c0.n20_adj_2547_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_1116_LC_1_19_2 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_1116_LC_1_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_1116_LC_1_19_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_adj_1116_LC_1_19_2  (
            .in0(N__17002),
            .in1(N__20600),
            .in2(N__17009),
            .in3(N__17516),
            .lcout(\c0.n8056 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i49_LC_1_19_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i49_LC_1_19_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i49_LC_1_19_3 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \c0.data_in_0___i49_LC_1_19_3  (
            .in0(N__23823),
            .in1(_gnd_net_),
            .in2(N__24605),
            .in3(N__45481),
            .lcout(data_in_6_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50255),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_857_LC_1_19_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_857_LC_1_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_857_LC_1_19_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_857_LC_1_19_4  (
            .in0(N__22002),
            .in1(N__28759),
            .in2(_gnd_net_),
            .in3(N__17498),
            .lcout(\c0.n9317 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_958_LC_1_19_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_958_LC_1_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_958_LC_1_19_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_958_LC_1_19_5  (
            .in0(N__28760),
            .in1(N__22406),
            .in2(N__27518),
            .in3(N__16991),
            .lcout(\c0.n17544 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_952_LC_1_19_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_952_LC_1_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_952_LC_1_19_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_952_LC_1_19_7  (
            .in0(_gnd_net_),
            .in1(N__25583),
            .in2(_gnd_net_),
            .in3(N__20073),
            .lcout(\c0.n17650 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_830_LC_1_20_1 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_830_LC_1_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_830_LC_1_20_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_830_LC_1_20_1  (
            .in0(N__19958),
            .in1(N__17452),
            .in2(N__17536),
            .in3(N__19859),
            .lcout(\c0.n8645 ),
            .ltout(\c0.n8645_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1089_LC_1_20_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1089_LC_1_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1089_LC_1_20_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1089_LC_1_20_2  (
            .in0(N__18706),
            .in1(N__17577),
            .in2(N__16979),
            .in3(N__19871),
            .lcout(\c0.n30_adj_2489 ),
            .ltout(\c0.n30_adj_2489_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1108_LC_1_20_3 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1108_LC_1_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1108_LC_1_20_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_1108_LC_1_20_3  (
            .in0(N__16976),
            .in1(N__22333),
            .in2(N__16967),
            .in3(N__17470),
            .lcout(\c0.n18_adj_2545 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_2_lut_LC_1_20_5 .C_ON=1'b0;
    defparam \c0.i15_2_lut_LC_1_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i15_2_lut_LC_1_20_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i15_2_lut_LC_1_20_5  (
            .in0(N__17578),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17451),
            .lcout(\c0.n9365 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i7_LC_1_20_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i7_LC_1_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i7_LC_1_20_6 .LUT_INIT=16'b0000110010101110;
    LogicCell40 \c0.data_out_frame2_0___i7_LC_1_20_6  (
            .in0(N__33170),
            .in1(N__17059),
            .in2(N__33678),
            .in3(N__23873),
            .lcout(\c0.data_out_frame2_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50257),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1090_LC_1_20_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1090_LC_1_20_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1090_LC_1_20_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1090_LC_1_20_7  (
            .in0(N__19959),
            .in1(N__22139),
            .in2(N__17582),
            .in3(N__18707),
            .lcout(\c0.n17516 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1074_LC_1_21_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1074_LC_1_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1074_LC_1_21_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1074_LC_1_21_0  (
            .in0(N__22225),
            .in1(N__23793),
            .in2(N__20074),
            .in3(N__22831),
            .lcout(\c0.n9204 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1034_LC_1_21_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1034_LC_1_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1034_LC_1_21_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1034_LC_1_21_1  (
            .in0(_gnd_net_),
            .in1(N__24955),
            .in2(_gnd_net_),
            .in3(N__21582),
            .lcout(\c0.n9328 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15831_3_lut_LC_1_21_2 .C_ON=1'b0;
    defparam \c0.i15831_3_lut_LC_1_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i15831_3_lut_LC_1_21_2 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \c0.i15831_3_lut_LC_1_21_2  (
            .in0(N__17548),
            .in1(N__30985),
            .in2(_gnd_net_),
            .in3(N__30564),
            .lcout(\c0.n18080 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i43_LC_1_21_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i43_LC_1_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i43_LC_1_21_3 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \c0.data_in_frame_0___i43_LC_1_21_3  (
            .in0(N__24721),
            .in1(N__24274),
            .in2(N__33038),
            .in3(N__31918),
            .lcout(data_in_frame_5_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50261),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i81_LC_1_21_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i81_LC_1_21_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i81_LC_1_21_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.data_in_frame_0___i81_LC_1_21_4  (
            .in0(_gnd_net_),
            .in1(N__24415),
            .in2(_gnd_net_),
            .in3(N__31917),
            .lcout(\c0.data_in_frame_10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50261),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1051_LC_1_21_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1051_LC_1_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1051_LC_1_21_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1051_LC_1_21_5  (
            .in0(N__24720),
            .in1(N__24956),
            .in2(_gnd_net_),
            .in3(N__21583),
            .lcout(\c0.n8976 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_832_LC_1_21_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_832_LC_1_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_832_LC_1_21_6 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \c0.i1_2_lut_adj_832_LC_1_21_6  (
            .in0(N__22553),
            .in1(_gnd_net_),
            .in2(N__21946),
            .in3(_gnd_net_),
            .lcout(\c0.n17513 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2272__i0_LC_1_22_0 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter2_2272__i0_LC_1_22_0 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_2272__i0_LC_1_22_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter2_2272__i0_LC_1_22_0  (
            .in0(_gnd_net_),
            .in1(N__19619),
            .in2(N__30625),
            .in3(_gnd_net_),
            .lcout(\c0.byte_transmit_counter2_0 ),
            .ltout(),
            .carryin(bfn_1_22_0_),
            .carryout(\c0.n16405 ),
            .clk(N__50266),
            .ce(N__17639),
            .sr(N__17627));
    defparam \c0.byte_transmit_counter2_2272__i1_LC_1_22_1 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter2_2272__i1_LC_1_22_1 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_2272__i1_LC_1_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter2_2272__i1_LC_1_22_1  (
            .in0(_gnd_net_),
            .in1(N__30930),
            .in2(_gnd_net_),
            .in3(N__17030),
            .lcout(\c0.byte_transmit_counter2_1 ),
            .ltout(),
            .carryin(\c0.n16405 ),
            .carryout(\c0.n16406 ),
            .clk(N__50266),
            .ce(N__17639),
            .sr(N__17627));
    defparam \c0.byte_transmit_counter2_2272__i2_LC_1_22_2 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter2_2272__i2_LC_1_22_2 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_2272__i2_LC_1_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter2_2272__i2_LC_1_22_2  (
            .in0(_gnd_net_),
            .in1(N__26758),
            .in2(_gnd_net_),
            .in3(N__17027),
            .lcout(\c0.byte_transmit_counter2_2 ),
            .ltout(),
            .carryin(\c0.n16406 ),
            .carryout(\c0.n16407 ),
            .clk(N__50266),
            .ce(N__17639),
            .sr(N__17627));
    defparam \c0.byte_transmit_counter2_2272__i3_LC_1_22_3 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter2_2272__i3_LC_1_22_3 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_2272__i3_LC_1_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter2_2272__i3_LC_1_22_3  (
            .in0(_gnd_net_),
            .in1(N__26602),
            .in2(_gnd_net_),
            .in3(N__17024),
            .lcout(\c0.byte_transmit_counter2_3 ),
            .ltout(),
            .carryin(\c0.n16407 ),
            .carryout(\c0.n16408 ),
            .clk(N__50266),
            .ce(N__17639),
            .sr(N__17627));
    defparam \c0.byte_transmit_counter2_2272__i4_LC_1_22_4 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter2_2272__i4_LC_1_22_4 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_2272__i4_LC_1_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter2_2272__i4_LC_1_22_4  (
            .in0(_gnd_net_),
            .in1(N__26455),
            .in2(_gnd_net_),
            .in3(N__17021),
            .lcout(\c0.byte_transmit_counter2_4 ),
            .ltout(),
            .carryin(\c0.n16408 ),
            .carryout(\c0.n16409 ),
            .clk(N__50266),
            .ce(N__17639),
            .sr(N__17627));
    defparam \c0.byte_transmit_counter2_2272__i5_LC_1_22_5 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter2_2272__i5_LC_1_22_5 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_2272__i5_LC_1_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter2_2272__i5_LC_1_22_5  (
            .in0(_gnd_net_),
            .in1(N__19687),
            .in2(_gnd_net_),
            .in3(N__17018),
            .lcout(\c0.byte_transmit_counter2_5 ),
            .ltout(),
            .carryin(\c0.n16409 ),
            .carryout(\c0.n16410 ),
            .clk(N__50266),
            .ce(N__17639),
            .sr(N__17627));
    defparam \c0.byte_transmit_counter2_2272__i6_LC_1_22_6 .C_ON=1'b1;
    defparam \c0.byte_transmit_counter2_2272__i6_LC_1_22_6 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_2272__i6_LC_1_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter2_2272__i6_LC_1_22_6  (
            .in0(_gnd_net_),
            .in1(N__19663),
            .in2(_gnd_net_),
            .in3(N__17015),
            .lcout(\c0.byte_transmit_counter2_6 ),
            .ltout(),
            .carryin(\c0.n16410 ),
            .carryout(\c0.n16411 ),
            .clk(N__50266),
            .ce(N__17639),
            .sr(N__17627));
    defparam \c0.byte_transmit_counter2_2272__i7_LC_1_22_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2272__i7_LC_1_22_7 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter2_2272__i7_LC_1_22_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.byte_transmit_counter2_2272__i7_LC_1_22_7  (
            .in0(_gnd_net_),
            .in1(N__19636),
            .in2(_gnd_net_),
            .in3(N__17012),
            .lcout(\c0.byte_transmit_counter2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50266),
            .ce(N__17639),
            .sr(N__17627));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16006_LC_1_23_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16006_LC_1_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16006_LC_1_23_0 .LUT_INIT=16'b1010111111000000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_16006_LC_1_23_0  (
            .in0(N__17894),
            .in1(N__25316),
            .in2(N__30964),
            .in3(N__30560),
            .lcout(\c0.n18474 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i131_LC_1_23_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i131_LC_1_23_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i131_LC_1_23_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i131_LC_1_23_1  (
            .in0(N__32816),
            .in1(N__34112),
            .in2(_gnd_net_),
            .in3(N__17245),
            .lcout(data_out_frame2_16_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50273),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15805_3_lut_LC_1_23_2 .C_ON=1'b0;
    defparam \c0.i15805_3_lut_LC_1_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i15805_3_lut_LC_1_23_2 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \c0.i15805_3_lut_LC_1_23_2  (
            .in0(N__30875),
            .in1(N__17077),
            .in2(_gnd_net_),
            .in3(N__30563),
            .lcout(\c0.n18074 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i1_LC_1_23_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i1_LC_1_23_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i1_LC_1_23_3 .LUT_INIT=16'b0000101011001110;
    LogicCell40 \c0.data_out_frame2_0___i1_LC_1_23_3  (
            .in0(N__17078),
            .in1(N__33159),
            .in2(N__33692),
            .in3(N__23881),
            .lcout(\c0.data_out_frame2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50273),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1080_LC_1_23_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1080_LC_1_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1080_LC_1_23_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1080_LC_1_23_4  (
            .in0(N__20380),
            .in1(N__18936),
            .in2(_gnd_net_),
            .in3(N__22960),
            .lcout(n9380),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i59_LC_1_23_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i59_LC_1_23_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i59_LC_1_23_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i59_LC_1_23_5  (
            .in0(N__32817),
            .in1(N__34769),
            .in2(_gnd_net_),
            .in3(N__17069),
            .lcout(data_out_frame2_7_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50273),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_2_i5_3_lut_LC_1_23_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_2_i5_3_lut_LC_1_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_2_i5_3_lut_LC_1_23_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_2_i5_3_lut_LC_1_23_6  (
            .in0(N__17068),
            .in1(N__17144),
            .in2(_gnd_net_),
            .in3(N__30561),
            .lcout(\c0.n5_adj_2463 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15818_3_lut_LC_1_23_7 .C_ON=1'b0;
    defparam \c0.i15818_3_lut_LC_1_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.i15818_3_lut_LC_1_23_7 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \c0.i15818_3_lut_LC_1_23_7  (
            .in0(N__30562),
            .in1(N__17060),
            .in2(_gnd_net_),
            .in3(N__30874),
            .lcout(\c0.n18078 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16066_LC_1_24_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16066_LC_1_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16066_LC_1_24_0 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_16066_LC_1_24_0  (
            .in0(N__19118),
            .in1(N__30979),
            .in2(N__17042),
            .in3(N__30669),
            .lcout(),
            .ltout(\c0.n18546_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18546_bdd_4_lut_LC_1_24_1 .C_ON=1'b0;
    defparam \c0.n18546_bdd_4_lut_LC_1_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.n18546_bdd_4_lut_LC_1_24_1 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n18546_bdd_4_lut_LC_1_24_1  (
            .in0(N__30980),
            .in1(N__17905),
            .in2(N__17045),
            .in3(N__17159),
            .lcout(\c0.n17803 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i91_LC_1_24_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i91_LC_1_24_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i91_LC_1_24_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i91_LC_1_24_2  (
            .in0(N__34765),
            .in1(N__18226),
            .in2(_gnd_net_),
            .in3(N__32821),
            .lcout(data_out_frame2_11_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50280),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i94_LC_1_24_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i94_LC_1_24_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i94_LC_1_24_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i94_LC_1_24_3  (
            .in0(N__32819),
            .in1(N__35603),
            .in2(_gnd_net_),
            .in3(N__17041),
            .lcout(data_out_frame2_11_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50280),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3957_3_lut_4_lut_LC_1_24_4 .C_ON=1'b0;
    defparam \c0.i3957_3_lut_4_lut_LC_1_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3957_3_lut_4_lut_LC_1_24_4 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \c0.i3957_3_lut_4_lut_LC_1_24_4  (
            .in0(N__20143),
            .in1(N__34684),
            .in2(N__23702),
            .in3(N__28066),
            .lcout(\c0.n2604 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18474_bdd_4_lut_LC_1_24_5 .C_ON=1'b0;
    defparam \c0.n18474_bdd_4_lut_LC_1_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.n18474_bdd_4_lut_LC_1_24_5 .LUT_INIT=16'b1101110010011000;
    LogicCell40 \c0.n18474_bdd_4_lut_LC_1_24_5  (
            .in0(N__30978),
            .in1(N__17126),
            .in2(N__19160),
            .in3(N__18998),
            .lcout(\c0.n17836 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i109_LC_1_24_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i109_LC_1_24_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i109_LC_1_24_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_out_frame2_0___i109_LC_1_24_6  (
            .in0(N__19540),
            .in1(N__36463),
            .in2(_gnd_net_),
            .in3(N__32820),
            .lcout(data_out_frame2_13_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50280),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i142_LC_1_24_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i142_LC_1_24_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i142_LC_1_24_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i142_LC_1_24_7  (
            .in0(N__32818),
            .in1(N__35602),
            .in2(_gnd_net_),
            .in3(N__17117),
            .lcout(data_out_frame2_17_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50280),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16056_LC_1_25_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16056_LC_1_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16056_LC_1_25_0 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_16056_LC_1_25_0  (
            .in0(N__17614),
            .in1(N__30986),
            .in2(N__20849),
            .in3(N__30670),
            .lcout(),
            .ltout(\c0.n18534_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18534_bdd_4_lut_LC_1_25_1 .C_ON=1'b0;
    defparam \c0.n18534_bdd_4_lut_LC_1_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.n18534_bdd_4_lut_LC_1_25_1 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n18534_bdd_4_lut_LC_1_25_1  (
            .in0(N__30987),
            .in1(N__17170),
            .in2(N__17120),
            .in3(N__17116),
            .lcout(),
            .ltout(\c0.n18537_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_5_i22_4_lut_LC_1_25_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_5_i22_4_lut_LC_1_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_5_i22_4_lut_LC_1_25_2 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_5_i22_4_lut_LC_1_25_2  (
            .in0(N__26782),
            .in1(N__19025),
            .in2(N__17105),
            .in3(N__26942),
            .lcout(\c0.n22_adj_2523 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15950_LC_1_25_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15950_LC_1_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15950_LC_1_25_3 .LUT_INIT=16'b1011110010001100;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_15950_LC_1_25_3  (
            .in0(N__17621),
            .in1(N__26783),
            .in2(N__26667),
            .in3(N__17102),
            .lcout(),
            .ltout(\c0.n18384_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18384_bdd_4_lut_LC_1_25_4 .C_ON=1'b0;
    defparam \c0.n18384_bdd_4_lut_LC_1_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.n18384_bdd_4_lut_LC_1_25_4 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n18384_bdd_4_lut_LC_1_25_4  (
            .in0(N__26624),
            .in1(N__17096),
            .in2(N__17087),
            .in3(N__18134),
            .lcout(),
            .ltout(\c0.n18387_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i5_LC_1_25_5 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i5_LC_1_25_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i5_LC_1_25_5 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \c0.tx2.r_Tx_Data_i5_LC_1_25_5  (
            .in0(N__17084),
            .in1(N__26625),
            .in2(N__17183),
            .in3(N__26476),
            .lcout(\c0.tx2.r_Tx_Data_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50285),
            .ce(N__26400),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_2_i6_4_lut_LC_1_26_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_2_i6_4_lut_LC_1_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_2_i6_4_lut_LC_1_26_0 .LUT_INIT=16'b1101100010001000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_2_i6_4_lut_LC_1_26_0  (
            .in0(N__30988),
            .in1(N__17180),
            .in2(N__17846),
            .in3(N__30672),
            .lcout(\c0.n6_adj_2466 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15824_3_lut_LC_1_26_1 .C_ON=1'b0;
    defparam \c0.i15824_3_lut_LC_1_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.i15824_3_lut_LC_1_26_1 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \c0.i15824_3_lut_LC_1_26_1  (
            .in0(N__30673),
            .in1(_gnd_net_),
            .in2(N__23249),
            .in3(N__30989),
            .lcout(\c0.n18084 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i46_LC_1_26_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i46_LC_1_26_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i46_LC_1_26_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i46_LC_1_26_2  (
            .in0(N__36409),
            .in1(N__18148),
            .in2(_gnd_net_),
            .in3(N__32651),
            .lcout(data_out_frame2_5_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50290),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i62_LC_1_26_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i62_LC_1_26_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i62_LC_1_26_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i62_LC_1_26_3  (
            .in0(N__32648),
            .in1(N__35595),
            .in2(_gnd_net_),
            .in3(N__17197),
            .lcout(data_out_frame2_7_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50290),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i134_LC_1_26_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i134_LC_1_26_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i134_LC_1_26_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i134_LC_1_26_4  (
            .in0(N__35099),
            .in1(N__17171),
            .in2(_gnd_net_),
            .in3(N__32650),
            .lcout(data_out_frame2_16_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50290),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i78_LC_1_26_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i78_LC_1_26_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i78_LC_1_26_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i78_LC_1_26_5  (
            .in0(N__32649),
            .in1(N__36410),
            .in2(_gnd_net_),
            .in3(N__17158),
            .lcout(data_out_frame2_9_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50290),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1128_LC_1_26_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1128_LC_1_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1128_LC_1_26_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1128_LC_1_26_6  (
            .in0(_gnd_net_),
            .in1(N__36547),
            .in2(_gnd_net_),
            .in3(N__25835),
            .lcout(\c0.n6_adj_2550 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i51_LC_1_26_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i51_LC_1_26_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i51_LC_1_26_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i51_LC_1_26_7  (
            .in0(N__32647),
            .in1(N__35306),
            .in2(_gnd_net_),
            .in3(N__17140),
            .lcout(data_out_frame2_6_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50290),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16016_LC_1_27_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16016_LC_1_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16016_LC_1_27_0 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_16016_LC_1_27_0  (
            .in0(N__20816),
            .in1(N__31033),
            .in2(N__29156),
            .in3(N__30671),
            .lcout(),
            .ltout(\c0.n18486_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18486_bdd_4_lut_LC_1_27_1 .C_ON=1'b0;
    defparam \c0.n18486_bdd_4_lut_LC_1_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.n18486_bdd_4_lut_LC_1_27_1 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n18486_bdd_4_lut_LC_1_27_1  (
            .in0(N__31034),
            .in1(N__17246),
            .in2(N__17231),
            .in3(N__19208),
            .lcout(),
            .ltout(\c0.n18489_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_2_i22_4_lut_LC_1_27_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_2_i22_4_lut_LC_1_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_2_i22_4_lut_LC_1_27_2 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_2_i22_4_lut_LC_1_27_2  (
            .in0(N__26843),
            .in1(N__20861),
            .in2(N__17228),
            .in3(N__26906),
            .lcout(\c0.n22_adj_2529 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15921_LC_1_27_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15921_LC_1_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15921_LC_1_27_3 .LUT_INIT=16'b1100111110100000;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_15921_LC_1_27_3  (
            .in0(N__19352),
            .in1(N__17768),
            .in2(N__26662),
            .in3(N__26844),
            .lcout(),
            .ltout(\c0.n18366_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18366_bdd_4_lut_LC_1_27_4 .C_ON=1'b0;
    defparam \c0.n18366_bdd_4_lut_LC_1_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.n18366_bdd_4_lut_LC_1_27_4 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n18366_bdd_4_lut_LC_1_27_4  (
            .in0(N__26626),
            .in1(N__17225),
            .in2(N__17219),
            .in3(N__17216),
            .lcout(),
            .ltout(\c0.n18369_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i2_LC_1_27_5 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i2_LC_1_27_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i2_LC_1_27_5 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \c0.tx2.r_Tx_Data_i2_LC_1_27_5  (
            .in0(N__17207),
            .in1(N__26627),
            .in2(N__17201),
            .in3(N__26500),
            .lcout(\c0.tx2.r_Tx_Data_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50298),
            .ce(N__26409),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_5_i5_3_lut_LC_1_28_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_5_i5_3_lut_LC_1_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_5_i5_3_lut_LC_1_28_0 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_5_i5_3_lut_LC_1_28_0  (
            .in0(N__30766),
            .in1(_gnd_net_),
            .in2(N__19181),
            .in3(N__17198),
            .lcout(\c0.n5_adj_2495 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i12_3_lut_LC_1_28_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i12_3_lut_LC_1_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i12_3_lut_LC_1_28_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_4_i12_3_lut_LC_1_28_1  (
            .in0(N__20996),
            .in1(N__30761),
            .in2(_gnd_net_),
            .in3(N__17938),
            .lcout(\c0.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16026_LC_1_28_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16026_LC_1_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16026_LC_1_28_2 .LUT_INIT=16'b1110010010101010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_16026_LC_1_28_2  (
            .in0(N__30760),
            .in1(N__17281),
            .in2(N__17828),
            .in3(N__30965),
            .lcout(\c0.n18492 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_1_i5_3_lut_LC_1_28_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_1_i5_3_lut_LC_1_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_1_i5_3_lut_LC_1_28_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_1_i5_3_lut_LC_1_28_3  (
            .in0(N__19310),
            .in1(N__30764),
            .in2(_gnd_net_),
            .in3(N__19229),
            .lcout(),
            .ltout(\c0.n5_adj_2503_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_1_i6_4_lut_LC_1_28_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_1_i6_4_lut_LC_1_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_1_i6_4_lut_LC_1_28_4 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_1_i6_4_lut_LC_1_28_4  (
            .in0(N__30765),
            .in1(N__18262),
            .in2(N__17285),
            .in3(N__30968),
            .lcout(\c0.n6_adj_2504 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16046_LC_1_28_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16046_LC_1_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16046_LC_1_28_5 .LUT_INIT=16'b1110011011000100;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_16046_LC_1_28_5  (
            .in0(N__30967),
            .in1(N__30763),
            .in2(N__18122),
            .in3(N__17950),
            .lcout(\c0.n18522 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16110_LC_1_28_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16110_LC_1_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16110_LC_1_28_6 .LUT_INIT=16'b1110011010100010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_16110_LC_1_28_6  (
            .in0(N__30762),
            .in1(N__30966),
            .in2(N__19484),
            .in3(N__17962),
            .lcout(\c0.n18600 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i115_LC_1_28_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i115_LC_1_28_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i115_LC_1_28_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_out_frame2_0___i115_LC_1_28_7  (
            .in0(N__17282),
            .in1(N__35298),
            .in2(_gnd_net_),
            .in3(N__32796),
            .lcout(data_out_frame2_14_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50306),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_LC_1_29_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_LC_1_29_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_LC_1_29_0 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_LC_1_29_0  (
            .in0(N__20834),
            .in1(N__30981),
            .in2(N__17810),
            .in3(N__30738),
            .lcout(),
            .ltout(\c0.n18606_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18606_bdd_4_lut_LC_1_29_1 .C_ON=1'b0;
    defparam \c0.n18606_bdd_4_lut_LC_1_29_1 .SEQ_MODE=4'b0000;
    defparam \c0.n18606_bdd_4_lut_LC_1_29_1 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n18606_bdd_4_lut_LC_1_29_1  (
            .in0(N__30982),
            .in1(N__18211),
            .in2(N__17273),
            .in3(N__30047),
            .lcout(\c0.n17779 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16086_LC_1_29_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16086_LC_1_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16086_LC_1_29_2 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_16086_LC_1_29_2  (
            .in0(N__18079),
            .in1(N__30983),
            .in2(N__17711),
            .in3(N__30739),
            .lcout(),
            .ltout(\c0.n18570_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18570_bdd_4_lut_LC_1_29_3 .C_ON=1'b0;
    defparam \c0.n18570_bdd_4_lut_LC_1_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.n18570_bdd_4_lut_LC_1_29_3 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n18570_bdd_4_lut_LC_1_29_3  (
            .in0(N__30984),
            .in1(N__20945),
            .in2(N__17270),
            .in3(N__19082),
            .lcout(),
            .ltout(\c0.n17773_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_LC_1_29_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_LC_1_29_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_LC_1_29_4 .LUT_INIT=16'b1011101111000000;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_LC_1_29_4  (
            .in0(N__17267),
            .in1(N__26619),
            .in2(N__17261),
            .in3(N__26784),
            .lcout(),
            .ltout(\c0.n18432_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18432_bdd_4_lut_LC_1_29_5 .C_ON=1'b0;
    defparam \c0.n18432_bdd_4_lut_LC_1_29_5 .SEQ_MODE=4'b0000;
    defparam \c0.n18432_bdd_4_lut_LC_1_29_5 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \c0.n18432_bdd_4_lut_LC_1_29_5  (
            .in0(N__17258),
            .in1(N__26661),
            .in2(N__17249),
            .in3(N__18293),
            .lcout(),
            .ltout(\c0.n18435_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i0_LC_1_29_6 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i0_LC_1_29_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i0_LC_1_29_6 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \c0.tx2.r_Tx_Data_i0_LC_1_29_6  (
            .in0(N__19454),
            .in1(N__26620),
            .in2(N__17336),
            .in3(N__26501),
            .lcout(\c0.tx2.r_Tx_Data_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50314),
            .ce(N__26405),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15916_LC_1_30_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15916_LC_1_30_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15916_LC_1_30_1 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_15916_LC_1_30_1  (
            .in0(N__19241),
            .in1(N__26616),
            .in2(N__17333),
            .in3(N__26780),
            .lcout(),
            .ltout(\c0.n18360_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18360_bdd_4_lut_LC_1_30_2 .C_ON=1'b0;
    defparam \c0.n18360_bdd_4_lut_LC_1_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.n18360_bdd_4_lut_LC_1_30_2 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n18360_bdd_4_lut_LC_1_30_2  (
            .in0(N__26617),
            .in1(N__30488),
            .in2(N__17318),
            .in3(N__17315),
            .lcout(\c0.n18363 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18468_bdd_4_lut_LC_1_30_3 .C_ON=1'b0;
    defparam \c0.n18468_bdd_4_lut_LC_1_30_3 .SEQ_MODE=4'b0000;
    defparam \c0.n18468_bdd_4_lut_LC_1_30_3 .LUT_INIT=16'b1100110010111000;
    LogicCell40 \c0.n18468_bdd_4_lut_LC_1_30_3  (
            .in0(N__17981),
            .in1(N__18269),
            .in2(N__18002),
            .in3(N__30990),
            .lcout(),
            .ltout(\c0.n18471_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_1_i22_4_lut_LC_1_30_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_1_i22_4_lut_LC_1_30_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_1_i22_4_lut_LC_1_30_4 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_1_i22_4_lut_LC_1_30_4  (
            .in0(N__26781),
            .in1(N__21044),
            .in2(N__17306),
            .in3(N__26933),
            .lcout(),
            .ltout(\c0.n22_adj_2530_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i1_LC_1_30_5 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i1_LC_1_30_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i1_LC_1_30_5 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \c0.tx2.r_Tx_Data_i1_LC_1_30_5  (
            .in0(N__17303),
            .in1(N__26618),
            .in2(N__17297),
            .in3(N__26518),
            .lcout(\c0.tx2.r_Tx_Data_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50323),
            .ce(N__26378),
            .sr(_gnd_net_));
    defparam \c0.tx2.add_59_2_lut_LC_1_31_0 .C_ON=1'b1;
    defparam \c0.tx2.add_59_2_lut_LC_1_31_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.add_59_2_lut_LC_1_31_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx2.add_59_2_lut_LC_1_31_0  (
            .in0(_gnd_net_),
            .in1(N__18605),
            .in2(_gnd_net_),
            .in3(N__17294),
            .lcout(n321),
            .ltout(),
            .carryin(bfn_1_31_0_),
            .carryout(\c0.tx2.n16372 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.add_59_3_lut_LC_1_31_1 .C_ON=1'b1;
    defparam \c0.tx2.add_59_3_lut_LC_1_31_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.add_59_3_lut_LC_1_31_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx2.add_59_3_lut_LC_1_31_1  (
            .in0(_gnd_net_),
            .in1(N__18397),
            .in2(_gnd_net_),
            .in3(N__17291),
            .lcout(n320),
            .ltout(),
            .carryin(\c0.tx2.n16372 ),
            .carryout(\c0.tx2.n16373 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.add_59_4_lut_LC_1_31_2 .C_ON=1'b1;
    defparam \c0.tx2.add_59_4_lut_LC_1_31_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.add_59_4_lut_LC_1_31_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx2.add_59_4_lut_LC_1_31_2  (
            .in0(_gnd_net_),
            .in1(N__18589),
            .in2(_gnd_net_),
            .in3(N__17288),
            .lcout(n319),
            .ltout(),
            .carryin(\c0.tx2.n16373 ),
            .carryout(\c0.tx2.n16374 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.add_59_5_lut_LC_1_31_3 .C_ON=1'b1;
    defparam \c0.tx2.add_59_5_lut_LC_1_31_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.add_59_5_lut_LC_1_31_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx2.add_59_5_lut_LC_1_31_3  (
            .in0(_gnd_net_),
            .in1(N__18554),
            .in2(_gnd_net_),
            .in3(N__17372),
            .lcout(n318),
            .ltout(),
            .carryin(\c0.tx2.n16374 ),
            .carryout(\c0.tx2.n16375 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.add_59_6_lut_LC_1_31_4 .C_ON=1'b1;
    defparam \c0.tx2.add_59_6_lut_LC_1_31_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.add_59_6_lut_LC_1_31_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx2.add_59_6_lut_LC_1_31_4  (
            .in0(_gnd_net_),
            .in1(N__18571),
            .in2(_gnd_net_),
            .in3(N__17369),
            .lcout(n317),
            .ltout(),
            .carryin(\c0.tx2.n16375 ),
            .carryout(\c0.tx2.n16376 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.add_59_7_lut_LC_1_31_5 .C_ON=1'b1;
    defparam \c0.tx2.add_59_7_lut_LC_1_31_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.add_59_7_lut_LC_1_31_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx2.add_59_7_lut_LC_1_31_5  (
            .in0(_gnd_net_),
            .in1(N__18538),
            .in2(_gnd_net_),
            .in3(N__17366),
            .lcout(n316),
            .ltout(),
            .carryin(\c0.tx2.n16376 ),
            .carryout(\c0.tx2.n16377 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.add_59_8_lut_LC_1_31_6 .C_ON=1'b1;
    defparam \c0.tx2.add_59_8_lut_LC_1_31_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.add_59_8_lut_LC_1_31_6 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx2.add_59_8_lut_LC_1_31_6  (
            .in0(N__18440),
            .in1(N__18499),
            .in2(_gnd_net_),
            .in3(N__17363),
            .lcout(\c0.tx2.n18013 ),
            .ltout(),
            .carryin(\c0.tx2.n16377 ),
            .carryout(\c0.tx2.n16378 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.add_59_9_lut_LC_1_31_7 .C_ON=1'b1;
    defparam \c0.tx2.add_59_9_lut_LC_1_31_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.add_59_9_lut_LC_1_31_7 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx2.add_59_9_lut_LC_1_31_7  (
            .in0(N__18438),
            .in1(N__18517),
            .in2(_gnd_net_),
            .in3(N__17360),
            .lcout(\c0.tx2.n17953 ),
            .ltout(),
            .carryin(\c0.tx2.n16378 ),
            .carryout(\c0.tx2.n16379 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.add_59_10_lut_LC_1_32_0 .C_ON=1'b0;
    defparam \c0.tx2.add_59_10_lut_LC_1_32_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.add_59_10_lut_LC_1_32_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx2.add_59_10_lut_LC_1_32_0  (
            .in0(N__18439),
            .in1(N__18477),
            .in2(_gnd_net_),
            .in3(N__17357),
            .lcout(\c0.tx2.n17939 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i7_LC_1_32_1 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i7_LC_1_32_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i7_LC_1_32_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.tx2.r_Clock_Count__i7_LC_1_32_1  (
            .in0(N__17354),
            .in1(N__21416),
            .in2(_gnd_net_),
            .in3(N__18518),
            .lcout(\c0.tx2.r_Clock_Count_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50342),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i6_LC_1_32_2 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i6_LC_1_32_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i6_LC_1_32_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.tx2.r_Clock_Count__i6_LC_1_32_2  (
            .in0(N__21415),
            .in1(N__18500),
            .in2(_gnd_net_),
            .in3(N__17348),
            .lcout(\c0.tx2.r_Clock_Count_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50342),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i8_LC_1_32_3 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i8_LC_1_32_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i8_LC_1_32_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.tx2.r_Clock_Count__i8_LC_1_32_3  (
            .in0(N__18478),
            .in1(N__21417),
            .in2(_gnd_net_),
            .in3(N__17342),
            .lcout(\c0.tx2.r_Clock_Count_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50342),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i5_LC_1_32_4 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i5_LC_1_32_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i5_LC_1_32_4 .LUT_INIT=16'b1100101000000000;
    LogicCell40 \c0.tx2.r_Clock_Count__i5_LC_1_32_4  (
            .in0(N__17405),
            .in1(N__18539),
            .in2(N__21432),
            .in3(N__18445),
            .lcout(r_Clock_Count_5_adj_2629),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50342),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i1_4_lut_4_lut_4_lut_LC_1_32_7 .C_ON=1'b0;
    defparam \c0.tx2.i1_4_lut_4_lut_4_lut_LC_1_32_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i1_4_lut_4_lut_4_lut_LC_1_32_7 .LUT_INIT=16'b1111000011111110;
    LogicCell40 \c0.tx2.i1_4_lut_4_lut_4_lut_LC_1_32_7  (
            .in0(N__21340),
            .in1(N__21266),
            .in2(N__21431),
            .in3(N__21470),
            .lcout(n10244),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16081_LC_2_17_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16081_LC_2_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16081_LC_2_17_0 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_16081_LC_2_17_0  (
            .in0(N__31030),
            .in1(N__17729),
            .in2(N__17879),
            .in3(N__30645),
            .lcout(\c0.n18564 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_991_LC_2_17_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_991_LC_2_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_991_LC_2_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_991_LC_2_17_2  (
            .in0(N__17391),
            .in1(N__21858),
            .in2(_gnd_net_),
            .in3(N__20426),
            .lcout(\c0.n17507 ),
            .ltout(\c0.n17507_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_914_LC_2_17_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_914_LC_2_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_914_LC_2_17_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_914_LC_2_17_3  (
            .in0(N__21772),
            .in1(N__19784),
            .in2(N__17399),
            .in3(N__18735),
            .lcout(\c0.n8687 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_6_i5_3_lut_LC_2_17_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_6_i5_3_lut_LC_2_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_6_i5_3_lut_LC_2_17_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_6_i5_3_lut_LC_2_17_4  (
            .in0(N__17927),
            .in1(N__17690),
            .in2(_gnd_net_),
            .in3(N__30644),
            .lcout(\c0.n5_adj_2515 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i36_LC_2_17_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i36_LC_2_17_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i36_LC_2_17_5 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \c0.data_in_frame_0___i36_LC_2_17_5  (
            .in0(N__20427),
            .in1(N__24218),
            .in2(N__27578),
            .in3(N__31979),
            .lcout(\c0.data_in_frame_4_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50252),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1047_LC_2_17_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1047_LC_2_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1047_LC_2_17_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1047_LC_2_17_6  (
            .in0(_gnd_net_),
            .in1(N__17390),
            .in2(_gnd_net_),
            .in3(N__21857),
            .lcout(\c0.n20_adj_2427 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16076_LC_2_17_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16076_LC_2_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16076_LC_2_17_7 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_16076_LC_2_17_7  (
            .in0(N__30643),
            .in1(N__17747),
            .in2(N__31084),
            .in3(N__17861),
            .lcout(\c0.n18558 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1098_LC_2_18_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1098_LC_2_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1098_LC_2_18_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1098_LC_2_18_0  (
            .in0(N__22548),
            .in1(N__21895),
            .in2(_gnd_net_),
            .in3(N__22637),
            .lcout(\c0.n2839 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_964_LC_2_18_1 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_964_LC_2_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_964_LC_2_18_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_964_LC_2_18_1  (
            .in0(N__17423),
            .in1(N__20611),
            .in2(N__20689),
            .in3(N__18789),
            .lcout(\c0.n12_adj_2492 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_973_LC_2_18_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_973_LC_2_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_973_LC_2_18_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_973_LC_2_18_2  (
            .in0(N__21907),
            .in1(N__18679),
            .in2(_gnd_net_),
            .in3(N__21839),
            .lcout(\c0.n9058 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_962_LC_2_18_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_962_LC_2_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_962_LC_2_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_962_LC_2_18_3  (
            .in0(N__28217),
            .in1(N__20668),
            .in2(_gnd_net_),
            .in3(N__19937),
            .lcout(\c0.n17476 ),
            .ltout(\c0.n17476_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_977_LC_2_18_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_977_LC_2_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_977_LC_2_18_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_977_LC_2_18_4  (
            .in0(N__25445),
            .in1(N__24884),
            .in2(N__17417),
            .in3(N__23773),
            .lcout(),
            .ltout(\c0.n17478_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_983_LC_2_18_5 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_983_LC_2_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_983_LC_2_18_5 .LUT_INIT=16'b1111100111110110;
    LogicCell40 \c0.i1_4_lut_adj_983_LC_2_18_5  (
            .in0(N__19880),
            .in1(N__17414),
            .in2(N__17408),
            .in3(N__20178),
            .lcout(\c0.n9_adj_2507 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i17_LC_2_19_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i17_LC_2_19_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i17_LC_2_19_0 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \c0.data_in_frame_0___i17_LC_2_19_0  (
            .in0(N__27122),
            .in1(N__24246),
            .in2(N__18662),
            .in3(N__31950),
            .lcout(\c0.data_in_frame_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50258),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i8_LC_2_19_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i8_LC_2_19_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i8_LC_2_19_1 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \c0.data_in_frame_0___i8_LC_2_19_1  (
            .in0(N__24245),
            .in1(N__18680),
            .in2(N__31981),
            .in3(N__21653),
            .lcout(\c0.data_in_frame_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50258),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i22_LC_2_19_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i22_LC_2_19_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i22_LC_2_19_2 .LUT_INIT=16'b0000000011001010;
    LogicCell40 \c0.data_in_frame_0___i22_LC_2_19_2  (
            .in0(N__26996),
            .in1(N__17500),
            .in2(N__24278),
            .in3(N__31951),
            .lcout(\c0.data_in_frame_2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50258),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1076_LC_2_19_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1076_LC_2_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1076_LC_2_19_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1076_LC_2_19_3  (
            .in0(N__23794),
            .in1(N__22952),
            .in2(N__18938),
            .in3(N__22839),
            .lcout(\c0.n17629 ),
            .ltout(\c0.n17629_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_2_lut_LC_2_19_4 .C_ON=1'b0;
    defparam \c0.i5_2_lut_LC_2_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i5_2_lut_LC_2_19_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i5_2_lut_LC_2_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17519),
            .in3(N__20402),
            .lcout(\c0.n16_adj_2546 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1020_LC_2_19_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1020_LC_2_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1020_LC_2_19_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1020_LC_2_19_5  (
            .in0(N__22670),
            .in1(N__22627),
            .in2(_gnd_net_),
            .in3(N__20099),
            .lcout(\c0.n9254 ),
            .ltout(\c0.n9254_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1002_LC_2_19_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1002_LC_2_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1002_LC_2_19_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1002_LC_2_19_6  (
            .in0(N__20437),
            .in1(N__20481),
            .in2(N__17504),
            .in3(N__17499),
            .lcout(\c0.n17522 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i20_LC_2_19_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i20_LC_2_19_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i20_LC_2_19_7 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \c0.data_in_frame_0___i20_LC_2_19_7  (
            .in0(N__24244),
            .in1(N__21723),
            .in2(N__31980),
            .in3(N__37573),
            .lcout(\c0.data_in_frame_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50258),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_939_LC_2_20_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_939_LC_2_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_939_LC_2_20_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_939_LC_2_20_0  (
            .in0(N__24931),
            .in1(N__20144),
            .in2(_gnd_net_),
            .in3(N__17471),
            .lcout(\c0.n8886 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i12_LC_2_20_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i12_LC_2_20_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i12_LC_2_20_1 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \c0.data_in_frame_0___i12_LC_2_20_1  (
            .in0(N__24275),
            .in1(N__27643),
            .in2(N__17459),
            .in3(N__31808),
            .lcout(\c0.data_in_frame_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50262),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i50_LC_2_20_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i50_LC_2_20_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i50_LC_2_20_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \c0.data_in_frame_0___i50_LC_2_20_2  (
            .in0(N__31806),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20186),
            .lcout(\c0.data_in_frame_6_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50262),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i65_LC_2_20_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i65_LC_2_20_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i65_LC_2_20_3 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \c0.data_in_frame_0___i65_LC_2_20_3  (
            .in0(N__28767),
            .in1(N__31804),
            .in2(N__23918),
            .in3(N__20261),
            .lcout(data_in_frame_8_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50262),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_6_i6_4_lut_LC_2_20_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_6_i6_4_lut_LC_2_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_6_i6_4_lut_LC_2_20_4 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_6_i6_4_lut_LC_2_20_4  (
            .in0(N__30758),
            .in1(N__20798),
            .in2(N__17438),
            .in3(N__31031),
            .lcout(\c0.n6_adj_2506 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i38_LC_2_20_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i38_LC_2_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i38_LC_2_20_5 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \c0.data_in_frame_0___i38_LC_2_20_5  (
            .in0(N__24276),
            .in1(N__21905),
            .in2(N__27215),
            .in3(N__31809),
            .lcout(\c0.data_in_frame_4_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50262),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i49_LC_2_20_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i49_LC_2_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i49_LC_2_20_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \c0.data_in_frame_0___i49_LC_2_20_6  (
            .in0(N__31805),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23777),
            .lcout(\c0.data_in_frame_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50262),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i42_LC_2_20_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i42_LC_2_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i42_LC_2_20_7 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \c0.data_in_frame_0___i42_LC_2_20_7  (
            .in0(N__24277),
            .in1(N__24963),
            .in2(N__39899),
            .in3(N__31807),
            .lcout(data_in_frame_5_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50262),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_913_LC_2_21_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_913_LC_2_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_913_LC_2_21_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_913_LC_2_21_0  (
            .in0(N__21773),
            .in1(N__22172),
            .in2(N__18743),
            .in3(N__22480),
            .lcout(\c0.n17467 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3963_3_lut_4_lut_LC_2_21_1 .C_ON=1'b0;
    defparam \c0.i3963_3_lut_4_lut_LC_2_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3963_3_lut_4_lut_LC_2_21_1 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \c0.i3963_3_lut_4_lut_LC_2_21_1  (
            .in0(N__21592),
            .in1(N__34673),
            .in2(N__22102),
            .in3(N__28062),
            .lcout(\c0.n2607 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3953_3_lut_4_lut_LC_2_21_2 .C_ON=1'b0;
    defparam \c0.i3953_3_lut_4_lut_LC_2_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3953_3_lut_4_lut_LC_2_21_2 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \c0.i3953_3_lut_4_lut_LC_2_21_2  (
            .in0(N__34674),
            .in1(N__29563),
            .in2(N__28067),
            .in3(N__18767),
            .lcout(\c0.n2602 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i6_LC_2_21_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i6_LC_2_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i6_LC_2_21_3 .LUT_INIT=16'b0000110010101110;
    LogicCell40 \c0.data_out_frame2_0___i6_LC_2_21_3  (
            .in0(N__33166),
            .in1(N__17549),
            .in2(N__33697),
            .in3(N__23866),
            .lcout(\c0.data_out_frame2_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50267),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i28_LC_2_21_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i28_LC_2_21_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i28_LC_2_21_4 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \c0.data_in_frame_0___i28_LC_2_21_4  (
            .in0(N__24259),
            .in1(N__27548),
            .in2(N__17537),
            .in3(N__31817),
            .lcout(\c0.data_in_frame_3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50267),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i13_LC_2_21_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i13_LC_2_21_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i13_LC_2_21_5 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \c0.data_in_frame_0___i13_LC_2_21_5  (
            .in0(N__19963),
            .in1(N__37661),
            .in2(N__31923),
            .in3(N__24261),
            .lcout(\c0.data_in_frame_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50267),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i41_LC_2_21_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i41_LC_2_21_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i41_LC_2_21_6 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \c0.data_in_frame_0___i41_LC_2_21_6  (
            .in0(N__24260),
            .in1(N__22098),
            .in2(N__21605),
            .in3(N__31816),
            .lcout(data_in_frame_5_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50267),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i46_LC_2_21_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i46_LC_2_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i46_LC_2_21_7 .LUT_INIT=16'b0000110000001010;
    LogicCell40 \c0.data_in_frame_0___i46_LC_2_21_7  (
            .in0(N__29564),
            .in1(N__18768),
            .in2(N__31922),
            .in3(N__24262),
            .lcout(data_in_frame_5_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50267),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_972_LC_2_22_0 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_972_LC_2_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_972_LC_2_22_0 .LUT_INIT=16'b1111011001101111;
    LogicCell40 \c0.i2_4_lut_adj_972_LC_2_22_0  (
            .in0(N__24556),
            .in1(N__17603),
            .in2(N__17597),
            .in3(N__17588),
            .lcout(\c0.n9_adj_2500 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i64_LC_2_22_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i64_LC_2_22_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i64_LC_2_22_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \c0.data_in_frame_0___i64_LC_2_22_1  (
            .in0(N__31831),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20033),
            .lcout(\c0.data_in_frame_7_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50274),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i48_LC_2_22_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i48_LC_2_22_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i48_LC_2_22_2 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \c0.data_in_frame_0___i48_LC_2_22_2  (
            .in0(N__24264),
            .in1(N__28315),
            .in2(N__36923),
            .in3(N__31838),
            .lcout(data_in_frame_5_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50274),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i52_LC_2_22_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i52_LC_2_22_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i52_LC_2_22_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \c0.data_in_frame_0___i52_LC_2_22_3  (
            .in0(N__31830),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22280),
            .lcout(\c0.data_in_frame_6_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50274),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i56_LC_2_22_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i56_LC_2_22_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i56_LC_2_22_4 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \c0.data_in_frame_0___i56_LC_2_22_4  (
            .in0(N__24263),
            .in1(N__36962),
            .in2(N__25107),
            .in3(N__31840),
            .lcout(\c0.data_in_frame_6_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50274),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i27_LC_2_22_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i27_LC_2_22_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i27_LC_2_22_5 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \c0.data_in_frame_0___i27_LC_2_22_5  (
            .in0(N__17576),
            .in1(N__37523),
            .in2(N__31926),
            .in3(N__24266),
            .lcout(\c0.data_in_frame_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50274),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i63_LC_2_22_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i63_LC_2_22_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i63_LC_2_22_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.data_in_frame_0___i63_LC_2_22_6  (
            .in0(_gnd_net_),
            .in1(N__22736),
            .in2(_gnd_net_),
            .in3(N__31839),
            .lcout(\c0.data_in_frame_7_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50274),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i25_LC_2_22_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i25_LC_2_22_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i25_LC_2_22_7 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \c0.data_in_frame_0___i25_LC_2_22_7  (
            .in0(N__22580),
            .in1(N__27839),
            .in2(N__31925),
            .in3(N__24265),
            .lcout(\c0.data_in_frame_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50274),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_982_LC_2_23_0 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_982_LC_2_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_982_LC_2_23_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i1_4_lut_adj_982_LC_2_23_0  (
            .in0(N__22241),
            .in1(N__22190),
            .in2(N__17558),
            .in3(N__17645),
            .lcout(),
            .ltout(\c0.n17325_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_984_LC_2_23_1 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_984_LC_2_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_984_LC_2_23_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i1_4_lut_adj_984_LC_2_23_1  (
            .in0(N__17666),
            .in1(N__24806),
            .in2(N__17657),
            .in3(N__18953),
            .lcout(\c0.n31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_970_LC_2_23_2 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_970_LC_2_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_970_LC_2_23_2 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \c0.i1_4_lut_adj_970_LC_2_23_2  (
            .in0(N__22767),
            .in1(N__20306),
            .in2(N__18907),
            .in3(N__22379),
            .lcout(),
            .ltout(\c0.n8_adj_2459_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_3_lut_4_lut_LC_2_23_3 .C_ON=1'b0;
    defparam \c0.i4_3_lut_4_lut_LC_2_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4_3_lut_4_lut_LC_2_23_3 .LUT_INIT=16'b1111100111110110;
    LogicCell40 \c0.i4_3_lut_4_lut_LC_2_23_3  (
            .in0(N__18863),
            .in1(N__19997),
            .in2(N__17654),
            .in3(N__17651),
            .lcout(\c0.n11_adj_2460 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15860_3_lut_4_lut_LC_2_23_4 .C_ON=1'b0;
    defparam \c0.i15860_3_lut_4_lut_LC_2_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i15860_3_lut_4_lut_LC_2_23_4 .LUT_INIT=16'b0000000000110100;
    LogicCell40 \c0.i15860_3_lut_4_lut_LC_2_23_4  (
            .in0(N__23198),
            .in1(N__33522),
            .in2(N__33379),
            .in3(N__33242),
            .lcout(\c0.n9605 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1086_LC_2_23_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1086_LC_2_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1086_LC_2_23_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1086_LC_2_23_5  (
            .in0(N__33241),
            .in1(N__33363),
            .in2(N__33529),
            .in3(N__23199),
            .lcout(\c0.n9900 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i107_LC_2_24_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i107_LC_2_24_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i107_LC_2_24_0 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \c0.data_out_frame2_0___i107_LC_2_24_0  (
            .in0(_gnd_net_),
            .in1(N__35828),
            .in2(N__17792),
            .in3(N__32764),
            .lcout(data_out_frame2_13_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50286),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18540_bdd_4_lut_LC_2_24_1 .C_ON=1'b0;
    defparam \c0.n18540_bdd_4_lut_LC_2_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.n18540_bdd_4_lut_LC_2_24_1 .LUT_INIT=16'b1111101001000100;
    LogicCell40 \c0.n18540_bdd_4_lut_LC_2_24_1  (
            .in0(N__30963),
            .in1(N__17758),
            .in2(N__19100),
            .in3(N__23627),
            .lcout(\c0.n17806 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i57_LC_2_24_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i57_LC_2_24_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i57_LC_2_24_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \c0.data_in_frame_0___i57_LC_2_24_2  (
            .in0(N__31919),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24575),
            .lcout(data_in_frame_7_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50286),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i150_LC_2_24_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i150_LC_2_24_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i150_LC_2_24_3 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \c0.data_out_frame2_0___i150_LC_2_24_3  (
            .in0(_gnd_net_),
            .in1(N__17615),
            .in2(N__32825),
            .in3(N__35098),
            .lcout(data_out_frame2_18_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50286),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18492_bdd_4_lut_LC_2_24_4 .C_ON=1'b0;
    defparam \c0.n18492_bdd_4_lut_LC_2_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.n18492_bdd_4_lut_LC_2_24_4 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \c0.n18492_bdd_4_lut_LC_2_24_4  (
            .in0(N__17788),
            .in1(N__30962),
            .in2(N__19013),
            .in3(N__17780),
            .lcout(\c0.n17827 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i102_LC_2_24_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i102_LC_2_24_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i102_LC_2_24_5 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \c0.data_out_frame2_0___i102_LC_2_24_5  (
            .in0(_gnd_net_),
            .in1(N__17759),
            .in2(N__32824),
            .in3(N__35097),
            .lcout(data_out_frame2_12_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50286),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_853_LC_2_24_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_853_LC_2_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_853_LC_2_24_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_853_LC_2_24_6  (
            .in0(N__25062),
            .in1(N__23050),
            .in2(_gnd_net_),
            .in3(N__19058),
            .lcout(\c0.n9043 ),
            .ltout(\c0.n9043_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_1120_LC_2_24_7 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_1120_LC_2_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_1120_LC_2_24_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_4_lut_adj_1120_LC_2_24_7  (
            .in0(N__22893),
            .in1(N__28316),
            .in2(N__17750),
            .in3(N__25073),
            .lcout(\c0.n17562 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i119_LC_2_25_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i119_LC_2_25_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i119_LC_2_25_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i119_LC_2_25_0  (
            .in0(N__36042),
            .in1(N__17743),
            .in2(_gnd_net_),
            .in3(N__32620),
            .lcout(data_out_frame2_14_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50291),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i41_LC_2_25_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i41_LC_2_25_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i41_LC_2_25_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i41_LC_2_25_1  (
            .in0(N__32617),
            .in1(N__35951),
            .in2(_gnd_net_),
            .in3(N__18310),
            .lcout(data_out_frame2_5_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50291),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i87_LC_2_25_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i87_LC_2_25_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i87_LC_2_25_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i87_LC_2_25_2  (
            .in0(N__36044),
            .in1(N__17725),
            .in2(_gnd_net_),
            .in3(N__32623),
            .lcout(data_out_frame2_10_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50291),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i89_LC_2_25_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i89_LC_2_25_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i89_LC_2_25_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i89_LC_2_25_3  (
            .in0(N__32619),
            .in1(N__34886),
            .in2(_gnd_net_),
            .in3(N__17704),
            .lcout(data_out_frame2_11_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50291),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i55_LC_2_25_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i55_LC_2_25_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i55_LC_2_25_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i55_LC_2_25_4  (
            .in0(N__36043),
            .in1(N__17680),
            .in2(_gnd_net_),
            .in3(N__32621),
            .lcout(data_out_frame2_6_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50291),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i63_LC_2_25_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i63_LC_2_25_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i63_LC_2_25_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i63_LC_2_25_5  (
            .in0(N__32618),
            .in1(N__35534),
            .in2(_gnd_net_),
            .in3(N__17920),
            .lcout(data_out_frame2_7_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50291),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i70_LC_2_25_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i70_LC_2_25_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i70_LC_2_25_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_out_frame2_0___i70_LC_2_25_6  (
            .in0(N__17906),
            .in1(N__35093),
            .in2(_gnd_net_),
            .in3(N__32622),
            .lcout(data_out_frame2_8_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50291),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i122_LC_2_25_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i122_LC_2_25_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i122_LC_2_25_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i122_LC_2_25_7  (
            .in0(N__32616),
            .in1(N__34829),
            .in2(_gnd_net_),
            .in3(N__17893),
            .lcout(data_out_frame2_15_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50291),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i95_LC_2_26_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i95_LC_2_26_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i95_LC_2_26_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i95_LC_2_26_0  (
            .in0(N__32757),
            .in1(N__35533),
            .in2(_gnd_net_),
            .in3(N__17875),
            .lcout(data_out_frame2_11_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50299),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i127_LC_2_26_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i127_LC_2_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i127_LC_2_26_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i127_LC_2_26_1  (
            .in0(N__35532),
            .in1(N__17860),
            .in2(_gnd_net_),
            .in3(N__32760),
            .lcout(data_out_frame2_15_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50299),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i43_LC_2_26_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i43_LC_2_26_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i43_LC_2_26_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i43_LC_2_26_2  (
            .in0(N__32754),
            .in1(N__35821),
            .in2(_gnd_net_),
            .in3(N__17842),
            .lcout(data_out_frame2_5_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50299),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i123_LC_2_26_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i123_LC_2_26_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i123_LC_2_26_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i123_LC_2_26_3  (
            .in0(N__34764),
            .in1(N__17824),
            .in2(_gnd_net_),
            .in3(N__32759),
            .lcout(data_out_frame2_15_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50299),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i71_LC_2_26_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i71_LC_2_26_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i71_LC_2_26_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i71_LC_2_26_4  (
            .in0(N__32755),
            .in1(N__35042),
            .in2(_gnd_net_),
            .in3(N__18025),
            .lcout(data_out_frame2_8_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50299),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i121_LC_2_26_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i121_LC_2_26_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i121_LC_2_26_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i121_LC_2_26_5  (
            .in0(N__34885),
            .in1(N__17806),
            .in2(_gnd_net_),
            .in3(N__32758),
            .lcout(data_out_frame2_15_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50299),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i83_LC_2_26_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i83_LC_2_26_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i83_LC_2_26_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i83_LC_2_26_6  (
            .in0(N__32756),
            .in1(N__35305),
            .in2(_gnd_net_),
            .in3(N__18250),
            .lcout(data_out_frame2_10_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50299),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18564_bdd_4_lut_LC_2_26_7 .C_ON=1'b0;
    defparam \c0.n18564_bdd_4_lut_LC_2_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.n18564_bdd_4_lut_LC_2_26_7 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \c0.n18564_bdd_4_lut_LC_2_26_7  (
            .in0(N__23378),
            .in1(N__31032),
            .in2(N__18026),
            .in3(N__18014),
            .lcout(\c0.n17794 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i146_LC_2_27_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i146_LC_2_27_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i146_LC_2_27_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i146_LC_2_27_0  (
            .in0(N__32626),
            .in1(N__34165),
            .in2(_gnd_net_),
            .in3(N__18283),
            .lcout(data_out_frame2_18_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50307),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i130_LC_2_27_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i130_LC_2_27_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i130_LC_2_27_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i130_LC_2_27_1  (
            .in0(N__34164),
            .in1(N__17998),
            .in2(_gnd_net_),
            .in3(N__32629),
            .lcout(data_out_frame2_16_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50307),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i137_LC_2_27_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i137_LC_2_27_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i137_LC_2_27_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i137_LC_2_27_2  (
            .in0(N__32625),
            .in1(N__34880),
            .in2(_gnd_net_),
            .in3(N__18064),
            .lcout(data_out_frame2_17_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50307),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i138_LC_2_27_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i138_LC_2_27_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i138_LC_2_27_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i138_LC_2_27_3  (
            .in0(N__34825),
            .in1(N__17977),
            .in2(_gnd_net_),
            .in3(N__32630),
            .lcout(data_out_frame2_17_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50307),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i129_LC_2_27_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i129_LC_2_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i129_LC_2_27_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i129_LC_2_27_4  (
            .in0(N__32624),
            .in1(N__34220),
            .in2(_gnd_net_),
            .in3(N__18046),
            .lcout(data_out_frame2_16_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50307),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i145_LC_2_27_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i145_LC_2_27_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i145_LC_2_27_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i145_LC_2_27_5  (
            .in0(N__34219),
            .in1(N__17963),
            .in2(_gnd_net_),
            .in3(N__32631),
            .lcout(data_out_frame2_18_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50307),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i84_LC_2_27_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i84_LC_2_27_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i84_LC_2_27_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i84_LC_2_27_6  (
            .in0(N__32627),
            .in1(N__35260),
            .in2(_gnd_net_),
            .in3(N__17951),
            .lcout(data_out_frame2_10_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50307),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i117_LC_2_27_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i117_LC_2_27_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i117_LC_2_27_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i117_LC_2_27_7  (
            .in0(N__36155),
            .in1(N__17939),
            .in2(_gnd_net_),
            .in3(N__32628),
            .lcout(data_out_frame2_14_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50307),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_5_i6_4_lut_LC_2_28_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_5_i6_4_lut_LC_2_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_5_i6_4_lut_LC_2_28_0 .LUT_INIT=16'b1010101011000000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_5_i6_4_lut_LC_2_28_0  (
            .in0(N__18161),
            .in1(N__30768),
            .in2(N__18155),
            .in3(N__31122),
            .lcout(\c0.n6_adj_2496 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i92_LC_2_28_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i92_LC_2_28_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i92_LC_2_28_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i92_LC_2_28_1  (
            .in0(N__35706),
            .in1(N__18121),
            .in2(_gnd_net_),
            .in3(N__32723),
            .lcout(data_out_frame2_11_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50315),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_954_LC_2_28_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_954_LC_2_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_954_LC_2_28_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_954_LC_2_28_2  (
            .in0(N__20461),
            .in1(N__18107),
            .in2(_gnd_net_),
            .in3(N__18098),
            .lcout(\c0.n8890 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i64_LC_2_28_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i64_LC_2_28_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i64_LC_2_28_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i64_LC_2_28_3  (
            .in0(N__45291),
            .in1(N__29800),
            .in2(_gnd_net_),
            .in3(N__32140),
            .lcout(data_in_7_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50315),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_993_LC_2_28_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_993_LC_2_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_993_LC_2_28_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i1_2_lut_adj_993_LC_2_28_4  (
            .in0(_gnd_net_),
            .in1(N__30767),
            .in2(_gnd_net_),
            .in3(N__31118),
            .lcout(\c0.n134 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i81_LC_2_28_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i81_LC_2_28_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i81_LC_2_28_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i81_LC_2_28_5  (
            .in0(N__35407),
            .in1(N__18080),
            .in2(_gnd_net_),
            .in3(N__32722),
            .lcout(data_out_frame2_10_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50315),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i53_LC_2_28_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i53_LC_2_28_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i53_LC_2_28_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i53_LC_2_28_6  (
            .in0(N__32721),
            .in1(N__36151),
            .in2(_gnd_net_),
            .in3(N__30214),
            .lcout(data_out_frame2_6_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50315),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_7_i6_4_lut_LC_2_28_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_7_i6_4_lut_LC_2_28_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_7_i6_4_lut_LC_2_28_7 .LUT_INIT=16'b1010110010100000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_7_i6_4_lut_LC_2_28_7  (
            .in0(N__20327),
            .in1(N__19192),
            .in2(N__31142),
            .in3(N__30769),
            .lcout(\c0.n6_adj_2464 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18600_bdd_4_lut_LC_2_29_0 .C_ON=1'b0;
    defparam \c0.n18600_bdd_4_lut_LC_2_29_0 .SEQ_MODE=4'b0000;
    defparam \c0.n18600_bdd_4_lut_LC_2_29_0 .LUT_INIT=16'b1110111001010000;
    LogicCell40 \c0.n18600_bdd_4_lut_LC_2_29_0  (
            .in0(N__31132),
            .in1(N__18068),
            .in2(N__18050),
            .in3(N__18032),
            .lcout(\c0.n18603 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_0_i5_3_lut_LC_2_29_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_0_i5_3_lut_LC_2_29_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_0_i5_3_lut_LC_2_29_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_0_i5_3_lut_LC_2_29_1  (
            .in0(N__30735),
            .in1(_gnd_net_),
            .in2(N__19328),
            .in3(N__19139),
            .lcout(),
            .ltout(\c0.n5_adj_2477_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_0_i6_4_lut_LC_2_29_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_0_i6_4_lut_LC_2_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_0_i6_4_lut_LC_2_29_2 .LUT_INIT=16'b1110010010100000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_0_i6_4_lut_LC_2_29_2  (
            .in0(N__31134),
            .in1(N__18314),
            .in2(N__18296),
            .in3(N__30737),
            .lcout(\c0.n6_adj_2436 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i151_LC_2_29_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i151_LC_2_29_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i151_LC_2_29_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i151_LC_2_29_3  (
            .in0(N__35029),
            .in1(N__18377),
            .in2(_gnd_net_),
            .in3(N__32810),
            .lcout(data_out_frame2_18_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50324),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16001_LC_2_29_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16001_LC_2_29_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16001_LC_2_29_4 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_16001_LC_2_29_4  (
            .in0(N__31133),
            .in1(N__18284),
            .in2(N__21032),
            .in3(N__30736),
            .lcout(\c0.n18468 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i42_LC_2_29_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i42_LC_2_29_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i42_LC_2_29_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i42_LC_2_29_5  (
            .in0(N__35886),
            .in1(N__18263),
            .in2(_gnd_net_),
            .in3(N__32811),
            .lcout(data_out_frame2_5_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50324),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16031_LC_2_29_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16031_LC_2_29_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16031_LC_2_29_6 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_16031_LC_2_29_6  (
            .in0(N__31131),
            .in1(N__18251),
            .in2(N__18236),
            .in3(N__30734),
            .lcout(\c0.n18504 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i97_LC_2_29_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i97_LC_2_29_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i97_LC_2_29_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i97_LC_2_29_7  (
            .in0(N__34213),
            .in1(N__18212),
            .in2(_gnd_net_),
            .in3(N__32812),
            .lcout(data_out_frame2_12_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50324),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15960_LC_2_30_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15960_LC_2_30_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15960_LC_2_30_1 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_15960_LC_2_30_1  (
            .in0(N__18200),
            .in1(N__26675),
            .in2(N__18815),
            .in3(N__26827),
            .lcout(),
            .ltout(\c0.n18408_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18408_bdd_4_lut_LC_2_30_2 .C_ON=1'b0;
    defparam \c0.n18408_bdd_4_lut_LC_2_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.n18408_bdd_4_lut_LC_2_30_2 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n18408_bdd_4_lut_LC_2_30_2  (
            .in0(N__26676),
            .in1(N__18191),
            .in2(N__18176),
            .in3(N__18173),
            .lcout(),
            .ltout(\c0.n18411_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i6_LC_2_30_3 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i6_LC_2_30_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i6_LC_2_30_3 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \c0.tx2.r_Tx_Data_i6_LC_2_30_3  (
            .in0(N__18359),
            .in1(N__26677),
            .in2(N__18380),
            .in3(N__26508),
            .lcout(\c0.tx2.r_Tx_Data_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50333),
            .ce(N__26377),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16071_LC_2_30_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16071_LC_2_30_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16071_LC_2_30_4 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_16071_LC_2_30_4  (
            .in0(N__31140),
            .in1(N__18376),
            .in2(N__21101),
            .in3(N__30733),
            .lcout(),
            .ltout(\c0.n18552_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18552_bdd_4_lut_LC_2_30_5 .C_ON=1'b0;
    defparam \c0.n18552_bdd_4_lut_LC_2_30_5 .SEQ_MODE=4'b0000;
    defparam \c0.n18552_bdd_4_lut_LC_2_30_5 .LUT_INIT=16'b1111000010101100;
    LogicCell40 \c0.n18552_bdd_4_lut_LC_2_30_5  (
            .in0(N__19555),
            .in1(N__19295),
            .in2(N__18365),
            .in3(N__31141),
            .lcout(),
            .ltout(\c0.n18555_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_6_i22_4_lut_LC_2_30_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_6_i22_4_lut_LC_2_30_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_6_i22_4_lut_LC_2_30_6 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_6_i22_4_lut_LC_2_30_6  (
            .in0(N__26826),
            .in1(N__20636),
            .in2(N__18362),
            .in3(N__26929),
            .lcout(\c0.n22_adj_2521 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i4_LC_2_31_0 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i4_LC_2_31_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i4_LC_2_31_0 .LUT_INIT=16'b1101100000000000;
    LogicCell40 \c0.tx2.r_Clock_Count__i4_LC_2_31_0  (
            .in0(N__21411),
            .in1(N__18570),
            .in2(N__18353),
            .in3(N__18444),
            .lcout(r_Clock_Count_4_adj_2630),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50343),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i3_LC_2_31_1 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i3_LC_2_31_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i3_LC_2_31_1 .LUT_INIT=16'b1010100000100000;
    LogicCell40 \c0.tx2.r_Clock_Count__i3_LC_2_31_1  (
            .in0(N__18441),
            .in1(N__21413),
            .in2(N__18344),
            .in3(N__18553),
            .lcout(r_Clock_Count_3_adj_2631),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50343),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i2_LC_2_31_2 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i2_LC_2_31_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i2_LC_2_31_2 .LUT_INIT=16'b1101100000000000;
    LogicCell40 \c0.tx2.r_Clock_Count__i2_LC_2_31_2  (
            .in0(N__21412),
            .in1(N__18590),
            .in2(N__18335),
            .in3(N__18443),
            .lcout(r_Clock_Count_2_adj_2632),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50343),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i2_3_lut_4_lut_LC_2_31_3 .C_ON=1'b0;
    defparam \c0.tx2.i2_3_lut_4_lut_LC_2_31_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i2_3_lut_4_lut_LC_2_31_3 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \c0.tx2.i2_3_lut_4_lut_LC_2_31_3  (
            .in0(N__21505),
            .in1(N__21347),
            .in2(N__21294),
            .in3(N__21409),
            .lcout(\c0.tx2.n7727 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i0_LC_2_31_4 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i0_LC_2_31_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i0_LC_2_31_4 .LUT_INIT=16'b1100100001000000;
    LogicCell40 \c0.tx2.r_Clock_Count__i0_LC_2_31_4  (
            .in0(N__21410),
            .in1(N__18442),
            .in2(N__18323),
            .in3(N__18604),
            .lcout(r_Clock_Count_0_adj_2634),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50343),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i4_4_lut_LC_2_31_5 .C_ON=1'b0;
    defparam \c0.tx2.i4_4_lut_LC_2_31_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i4_4_lut_LC_2_31_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.tx2.i4_4_lut_LC_2_31_5  (
            .in0(N__18603),
            .in1(N__18588),
            .in2(N__18572),
            .in3(N__18552),
            .lcout(),
            .ltout(\c0.tx2.n10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i5_3_lut_LC_2_31_6 .C_ON=1'b0;
    defparam \c0.tx2.i5_3_lut_LC_2_31_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i5_3_lut_LC_2_31_6 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \c0.tx2.i5_3_lut_LC_2_31_6  (
            .in0(N__18537),
            .in1(_gnd_net_),
            .in2(N__18521),
            .in3(N__18396),
            .lcout(\c0.tx2.n16452 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i11588211_i1_3_lut_LC_2_31_7 .C_ON=1'b0;
    defparam \c0.tx2.i11588211_i1_3_lut_LC_2_31_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i11588211_i1_3_lut_LC_2_31_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.tx2.i11588211_i1_3_lut_LC_2_31_7  (
            .in0(N__25889),
            .in1(N__19568),
            .in2(_gnd_net_),
            .in3(N__19490),
            .lcout(\c0.tx2.o_Tx_Serial_N_2354 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i15730_2_lut_3_lut_LC_2_32_0 .C_ON=1'b0;
    defparam \c0.tx2.i15730_2_lut_3_lut_LC_2_32_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i15730_2_lut_3_lut_LC_2_32_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.tx2.i15730_2_lut_3_lut_LC_2_32_0  (
            .in0(N__25884),
            .in1(N__26181),
            .in2(_gnd_net_),
            .in3(N__21465),
            .lcout(\c0.tx2.n17990 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i2_4_lut_LC_2_32_1 .C_ON=1'b0;
    defparam \c0.tx2.i2_4_lut_LC_2_32_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i2_4_lut_LC_2_32_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.tx2.i2_4_lut_LC_2_32_1  (
            .in0(N__18516),
            .in1(N__18498),
            .in2(N__18482),
            .in3(N__18461),
            .lcout(\c0.tx2.r_SM_Main_2_N_2323_1 ),
            .ltout(\c0.tx2.r_SM_Main_2_N_2323_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_i1_LC_2_32_2 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_i1_LC_2_32_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_SM_Main_i1_LC_2_32_2 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \c0.tx2.r_SM_Main_i1_LC_2_32_2  (
            .in0(N__21284),
            .in1(N__21342),
            .in2(N__18455),
            .in3(N__21425),
            .lcout(\c0.tx2.r_SM_Main_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50353),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_i2_LC_2_32_3 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_i2_LC_2_32_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_SM_Main_i2_LC_2_32_3 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \c0.tx2.r_SM_Main_i2_LC_2_32_3  (
            .in0(N__21343),
            .in1(N__21466),
            .in2(N__21433),
            .in3(N__21283),
            .lcout(r_SM_Main_2_adj_2628),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50353),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i1_LC_2_32_4 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i1_LC_2_32_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i1_LC_2_32_4 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \c0.tx2.r_Clock_Count__i1_LC_2_32_4  (
            .in0(N__18452),
            .in1(N__21421),
            .in2(N__18401),
            .in3(N__18446),
            .lcout(r_Clock_Count_1_adj_2633),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50353),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i9901_3_lut_LC_2_32_6 .C_ON=1'b0;
    defparam \c0.tx2.i9901_3_lut_LC_2_32_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i9901_3_lut_LC_2_32_6 .LUT_INIT=16'b1100110010111011;
    LogicCell40 \c0.tx2.i9901_3_lut_LC_2_32_6  (
            .in0(N__18614),
            .in1(N__21279),
            .in2(_gnd_net_),
            .in3(N__21341),
            .lcout(),
            .ltout(\c0.tx2.n12306_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.o_Tx_Serial_45_LC_2_32_7 .C_ON=1'b0;
    defparam \c0.tx2.o_Tx_Serial_45_LC_2_32_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.o_Tx_Serial_45_LC_2_32_7 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \c0.tx2.o_Tx_Serial_45_LC_2_32_7  (
            .in0(_gnd_net_),
            .in1(N__21414),
            .in2(N__18608),
            .in3(N__21135),
            .lcout(tx2_o),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50353),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i1_LC_3_17_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i1_LC_3_17_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i1_LC_3_17_0 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i1_LC_3_17_0  (
            .in0(N__33378),
            .in1(N__33515),
            .in2(N__33698),
            .in3(N__33229),
            .lcout(\c0.FRAME_MATCHER_state_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50254),
            .ce(),
            .sr(N__33413));
    defparam \c0.i3945_3_lut_LC_3_17_1 .C_ON=1'b0;
    defparam \c0.i3945_3_lut_LC_3_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3945_3_lut_LC_3_17_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.i3945_3_lut_LC_3_17_1  (
            .in0(N__39932),
            .in1(N__22009),
            .in2(_gnd_net_),
            .in3(N__24217),
            .lcout(n2598),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_859_LC_3_17_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_859_LC_3_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_859_LC_3_17_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_859_LC_3_17_2  (
            .in0(_gnd_net_),
            .in1(N__47648),
            .in2(_gnd_net_),
            .in3(N__41807),
            .lcout(\c0.n8600 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_894_LC_3_17_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_894_LC_3_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_894_LC_3_17_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_894_LC_3_17_3  (
            .in0(_gnd_net_),
            .in1(N__21552),
            .in2(_gnd_net_),
            .in3(N__22046),
            .lcout(\c0.n17424 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_986_LC_3_17_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_986_LC_3_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_986_LC_3_17_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_986_LC_3_17_4  (
            .in0(_gnd_net_),
            .in1(N__19753),
            .in2(_gnd_net_),
            .in3(N__18640),
            .lcout(\c0.n17614 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.equal_100_i4_2_lut_LC_3_17_6 .C_ON=1'b0;
    defparam \c0.rx.equal_100_i4_2_lut_LC_3_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.equal_100_i4_2_lut_LC_3_17_6 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \c0.rx.equal_100_i4_2_lut_LC_3_17_6  (
            .in0(N__39241),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39313),
            .lcout(n4_adj_2582),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.equal_102_i4_2_lut_LC_3_17_7 .C_ON=1'b0;
    defparam \c0.rx.equal_102_i4_2_lut_LC_3_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.equal_102_i4_2_lut_LC_3_17_7 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \c0.rx.equal_102_i4_2_lut_LC_3_17_7  (
            .in0(N__39314),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39240),
            .lcout(n4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i62_LC_3_18_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i62_LC_3_18_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i62_LC_3_18_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i62_LC_3_18_0  (
            .in0(N__20729),
            .in1(N__45482),
            .in2(_gnd_net_),
            .in3(N__36210),
            .lcout(data_in_7_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50259),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_965_LC_3_18_1 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_965_LC_3_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_965_LC_3_18_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_965_LC_3_18_1  (
            .in0(N__19807),
            .in1(N__18686),
            .in2(N__29133),
            .in3(N__20528),
            .lcout(\c0.n9334 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i6_LC_3_18_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i6_LC_3_18_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i6_LC_3_18_2 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \c0.data_in_frame_0___i6_LC_3_18_2  (
            .in0(N__37616),
            .in1(N__24270),
            .in2(N__21868),
            .in3(N__31876),
            .lcout(\c0.data_in_frame_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50259),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_961_LC_3_18_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_961_LC_3_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_961_LC_3_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_961_LC_3_18_3  (
            .in0(N__18678),
            .in1(N__18731),
            .in2(_gnd_net_),
            .in3(N__18657),
            .lcout(\c0.n9349 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i15_LC_3_18_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i15_LC_3_18_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i15_LC_3_18_4 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \c0.data_in_frame_0___i15_LC_3_18_4  (
            .in0(N__27797),
            .in1(N__24269),
            .in2(N__19904),
            .in3(N__31875),
            .lcout(\c0.data_in_frame_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50259),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i32_LC_3_18_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i32_LC_3_18_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i32_LC_3_18_5 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \c0.data_in_frame_0___i32_LC_3_18_5  (
            .in0(N__24268),
            .in1(N__18641),
            .in2(N__31943),
            .in3(N__23954),
            .lcout(\c0.data_in_frame_3_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50259),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1026_LC_3_18_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1026_LC_3_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1026_LC_3_18_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1026_LC_3_18_6  (
            .in0(N__18658),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18638),
            .lcout(\c0.n17553 ),
            .ltout(\c0.n17553_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_994_LC_3_18_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_994_LC_3_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_994_LC_3_18_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_994_LC_3_18_7  (
            .in0(N__22134),
            .in1(N__29122),
            .in2(N__18644),
            .in3(N__19898),
            .lcout(\c0.n8658 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1033_LC_3_19_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1033_LC_3_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1033_LC_3_19_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1033_LC_3_19_0  (
            .in0(N__21685),
            .in1(N__19754),
            .in2(N__21764),
            .in3(N__18639),
            .lcout(\c0.n25_adj_2491 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_933_LC_3_19_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_933_LC_3_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_933_LC_3_19_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_933_LC_3_19_1  (
            .in0(_gnd_net_),
            .in1(N__22485),
            .in2(_gnd_net_),
            .in3(N__22669),
            .lcout(\c0.n17406 ),
            .ltout(\c0.n17406_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_936_LC_3_19_2 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_936_LC_3_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_936_LC_3_19_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_4_lut_adj_936_LC_3_19_2  (
            .in0(N__18855),
            .in1(N__22591),
            .in2(N__18617),
            .in3(N__21837),
            .lcout(\c0.n17656 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i2_LC_3_19_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i2_LC_3_19_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i2_LC_3_19_3 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \c0.data_in_frame_0___i2_LC_3_19_3  (
            .in0(N__24240),
            .in1(N__29126),
            .in2(N__31941),
            .in3(N__27077),
            .lcout(\c0.data_in_frame_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50263),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i1_LC_3_19_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i1_LC_3_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i1_LC_3_19_4 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \c0.data_in_frame_0___i1_LC_3_19_4  (
            .in0(N__23984),
            .in1(N__24242),
            .in2(N__18883),
            .in3(N__31870),
            .lcout(\c0.data_in_frame_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50263),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_846_LC_3_19_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_846_LC_3_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_846_LC_3_19_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_846_LC_3_19_5  (
            .in0(_gnd_net_),
            .in1(N__18876),
            .in2(_gnd_net_),
            .in3(N__18769),
            .lcout(\c0.n23_adj_2426 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i21_LC_3_19_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i21_LC_3_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i21_LC_3_19_6 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \c0.data_in_frame_0___i21_LC_3_19_6  (
            .in0(N__27325),
            .in1(N__24243),
            .in2(N__18739),
            .in3(N__31871),
            .lcout(\c0.data_in_frame_2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50263),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i35_LC_3_19_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i35_LC_3_19_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i35_LC_3_19_7 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \c0.data_in_frame_0___i35_LC_3_19_7  (
            .in0(N__24241),
            .in1(N__29858),
            .in2(N__31942),
            .in3(N__21754),
            .lcout(\c0.data_in_frame_4_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50263),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i14_LC_3_20_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i14_LC_3_20_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i14_LC_3_20_0 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \c0.data_in_frame_0___i14_LC_3_20_0  (
            .in0(N__18705),
            .in1(N__36259),
            .in2(N__31850),
            .in3(N__24213),
            .lcout(\c0.data_in_frame_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50268),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_942_LC_3_20_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_942_LC_3_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_942_LC_3_20_1 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_942_LC_3_20_1  (
            .in0(N__34660),
            .in1(N__34452),
            .in2(_gnd_net_),
            .in3(N__31712),
            .lcout(n9419),
            .ltout(n9419_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i67_LC_3_20_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i67_LC_3_20_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i67_LC_3_20_2 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \c0.data_in_frame_0___i67_LC_3_20_2  (
            .in0(N__31713),
            .in1(N__33941),
            .in2(N__18689),
            .in3(N__22953),
            .lcout(data_in_frame_8_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50268),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i47_LC_3_20_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i47_LC_3_20_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i47_LC_3_20_3 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \c0.data_in_frame_0___i47_LC_3_20_3  (
            .in0(N__24212),
            .in1(N__31271),
            .in2(N__24677),
            .in3(N__31723),
            .lcout(data_in_frame_5_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50268),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i23_LC_3_20_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i23_LC_3_20_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i23_LC_3_20_4 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \c0.data_in_frame_0___i23_LC_3_20_4  (
            .in0(N__22484),
            .in1(N__27718),
            .in2(N__31851),
            .in3(N__24214),
            .lcout(\c0.data_in_frame_2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50268),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1087_LC_3_20_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1087_LC_3_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1087_LC_3_20_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1087_LC_3_20_5  (
            .in0(N__29056),
            .in1(N__18793),
            .in2(N__20570),
            .in3(N__21722),
            .lcout(\c0.n17569 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i39_LC_3_20_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i39_LC_3_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i39_LC_3_20_6 .LUT_INIT=16'b0000110000001010;
    LogicCell40 \c0.data_in_frame_0___i39_LC_3_20_6  (
            .in0(N__28384),
            .in1(N__22628),
            .in2(N__31852),
            .in3(N__24215),
            .lcout(\c0.data_in_frame_4_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50268),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12308_3_lut_LC_3_20_7 .C_ON=1'b0;
    defparam \c0.i12308_3_lut_LC_3_20_7 .SEQ_MODE=4'b0000;
    defparam \c0.i12308_3_lut_LC_3_20_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.i12308_3_lut_LC_3_20_7  (
            .in0(N__33508),
            .in1(N__25133),
            .in2(_gnd_net_),
            .in3(N__23263),
            .lcout(\c0.n81 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i70_LC_3_21_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i70_LC_3_21_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i70_LC_3_21_0 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \c0.data_in_frame_0___i70_LC_3_21_0  (
            .in0(N__31790),
            .in1(N__20728),
            .in2(N__20276),
            .in3(N__19053),
            .lcout(data_in_frame_8_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50275),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i61_LC_3_21_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i61_LC_3_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i61_LC_3_21_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.data_in_frame_0___i61_LC_3_21_1  (
            .in0(_gnd_net_),
            .in1(N__27473),
            .in2(_gnd_net_),
            .in3(N__31796),
            .lcout(\c0.data_in_frame_7_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50275),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i30_LC_3_21_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i30_LC_3_21_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i30_LC_3_21_2 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \c0.data_in_frame_0___i30_LC_3_21_2  (
            .in0(N__25385),
            .in1(N__27182),
            .in2(N__31920),
            .in3(N__24267),
            .lcout(\c0.data_in_frame_3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50275),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i71_LC_3_21_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i71_LC_3_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i71_LC_3_21_3 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \c0.data_in_frame_0___i71_LC_3_21_3  (
            .in0(N__28438),
            .in1(N__31791),
            .in2(N__38768),
            .in3(N__20273),
            .lcout(data_in_frame_8_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50275),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i69_LC_3_21_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i69_LC_3_21_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i69_LC_3_21_4 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \c0.data_in_frame_0___i69_LC_3_21_4  (
            .in0(N__31789),
            .in1(N__38384),
            .in2(N__20275),
            .in3(N__25052),
            .lcout(data_in_frame_8_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50275),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1017_LC_3_21_5 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1017_LC_3_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1017_LC_3_21_5 .LUT_INIT=16'b1111000011110100;
    LogicCell40 \c0.i1_4_lut_adj_1017_LC_3_21_5  (
            .in0(N__33387),
            .in1(N__33217),
            .in2(N__32826),
            .in3(N__23859),
            .lcout(n1396),
            .ltout(n1396_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i88_LC_3_21_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i88_LC_3_21_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i88_LC_3_21_6 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \c0.data_in_frame_0___i88_LC_3_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18839),
            .in3(N__23156),
            .lcout(\c0.data_in_frame_10_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50275),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i53_LC_3_21_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i53_LC_3_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i53_LC_3_21_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.data_in_frame_0___i53_LC_3_21_7  (
            .in0(_gnd_net_),
            .in1(N__18908),
            .in2(_gnd_net_),
            .in3(N__31795),
            .lcout(\c0.data_in_frame_6_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50275),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3927_3_lut_4_lut_LC_3_22_0 .C_ON=1'b0;
    defparam \c0.i3927_3_lut_4_lut_LC_3_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3927_3_lut_4_lut_LC_3_22_0 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \c0.i3927_3_lut_4_lut_LC_3_22_0  (
            .in0(N__33764),
            .in1(N__34675),
            .in2(N__28631),
            .in3(N__28058),
            .lcout(n2589),
            .ltout(n2589_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_899_LC_3_22_1 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_899_LC_3_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_899_LC_3_22_1 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \c0.i7_4_lut_adj_899_LC_3_22_1  (
            .in0(N__25502),
            .in1(N__24782),
            .in2(N__18836),
            .in3(N__18903),
            .lcout(\c0.n23_adj_2462 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i74_LC_3_22_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i74_LC_3_22_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i74_LC_3_22_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.data_in_frame_0___i74_LC_3_22_2  (
            .in0(_gnd_net_),
            .in1(N__28826),
            .in2(_gnd_net_),
            .in3(N__31822),
            .lcout(\c0.data_in_frame_9_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50281),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i54_LC_3_22_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i54_LC_3_22_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i54_LC_3_22_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \c0.data_in_frame_0___i54_LC_3_22_3  (
            .in0(N__31818),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27947),
            .lcout(data_in_frame_6_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50281),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i59_LC_3_22_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i59_LC_3_22_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i59_LC_3_22_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.data_in_frame_0___i59_LC_3_22_4  (
            .in0(_gnd_net_),
            .in1(N__18833),
            .in2(_gnd_net_),
            .in3(N__31821),
            .lcout(\c0.data_in_frame_7_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50281),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i62_LC_3_22_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i62_LC_3_22_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i62_LC_3_22_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \c0.data_in_frame_0___i62_LC_3_22_5  (
            .in0(N__31819),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22352),
            .lcout(\c0.data_in_frame_7_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50281),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i51_LC_3_22_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i51_LC_3_22_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i51_LC_3_22_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.data_in_frame_0___i51_LC_3_22_6  (
            .in0(_gnd_net_),
            .in1(N__24908),
            .in2(_gnd_net_),
            .in3(N__31820),
            .lcout(\c0.data_in_frame_6_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50281),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18558_bdd_4_lut_LC_3_22_7 .C_ON=1'b0;
    defparam \c0.n18558_bdd_4_lut_LC_3_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.n18558_bdd_4_lut_LC_3_22_7 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \c0.n18558_bdd_4_lut_LC_3_22_7  (
            .in0(N__20966),
            .in1(N__30991),
            .in2(N__20759),
            .in3(N__18827),
            .lcout(\c0.n17797 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1095_LC_3_23_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1095_LC_3_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1095_LC_3_23_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1095_LC_3_23_0  (
            .in0(N__28477),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22832),
            .lcout(\c0.n9028 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_979_LC_3_23_1 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_979_LC_3_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_979_LC_3_23_1 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \c0.i2_4_lut_adj_979_LC_3_23_1  (
            .in0(N__18980),
            .in1(N__25232),
            .in2(N__18965),
            .in3(N__27946),
            .lcout(\c0.n10_adj_2505 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1092_LC_3_23_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1092_LC_3_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1092_LC_3_23_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1092_LC_3_23_3  (
            .in0(N__28340),
            .in1(N__25345),
            .in2(_gnd_net_),
            .in3(N__20136),
            .lcout(\c0.n8061 ),
            .ltout(\c0.n8061_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1099_LC_3_23_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1099_LC_3_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1099_LC_3_23_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1099_LC_3_23_4  (
            .in0(N__18947),
            .in1(N__28621),
            .in2(N__18941),
            .in3(N__20579),
            .lcout(\c0.n17538 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3939_3_lut_4_lut_LC_3_23_5 .C_ON=1'b0;
    defparam \c0.i3939_3_lut_4_lut_LC_3_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3939_3_lut_4_lut_LC_3_23_5 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \c0.i3939_3_lut_4_lut_LC_3_23_5  (
            .in0(N__18937),
            .in1(N__34672),
            .in2(N__27437),
            .in3(N__28052),
            .lcout(n2595),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_896_LC_3_23_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_896_LC_3_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_896_LC_3_23_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_896_LC_3_23_6  (
            .in0(_gnd_net_),
            .in1(N__29084),
            .in2(_gnd_net_),
            .in3(N__18884),
            .lcout(\c0.n9039 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_967_LC_3_23_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_967_LC_3_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_967_LC_3_23_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_967_LC_3_23_7  (
            .in0(N__28432),
            .in1(N__28476),
            .in2(_gnd_net_),
            .in3(N__25461),
            .lcout(\c0.n9279 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i164_LC_3_24_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i164_LC_3_24_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i164_LC_3_24_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_frame2_0___i164_LC_3_24_0  (
            .in0(N__24315),
            .in1(N__32985),
            .in2(N__36557),
            .in3(N__25207),
            .lcout(\c0.data_out_frame2_20_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50292),
            .ce(N__32771),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_903_LC_3_24_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_903_LC_3_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_903_LC_3_24_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_903_LC_3_24_1  (
            .in0(N__19996),
            .in1(N__21608),
            .in2(_gnd_net_),
            .in3(N__18862),
            .lcout(\c0.n9151 ),
            .ltout(\c0.n9151_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_850_LC_3_24_2 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_850_LC_3_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_850_LC_3_24_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_850_LC_3_24_2  (
            .in0(N__19031),
            .in1(N__25106),
            .in2(N__19064),
            .in3(N__22805),
            .lcout(\c0.n17588 ),
            .ltout(\c0.n17588_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i156_LC_3_24_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i156_LC_3_24_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i156_LC_3_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_out_frame2_0___i156_LC_3_24_3  (
            .in0(_gnd_net_),
            .in1(N__32984),
            .in2(N__19061),
            .in3(N__32213),
            .lcout(\c0.data_out_frame2_19_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50292),
            .ce(N__32771),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_849_LC_3_24_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_849_LC_3_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_849_LC_3_24_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_849_LC_3_24_4  (
            .in0(_gnd_net_),
            .in1(N__28433),
            .in2(_gnd_net_),
            .in3(N__19057),
            .lcout(\c0.n6_adj_2429 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i166_LC_3_24_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i166_LC_3_24_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i166_LC_3_24_6 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.data_out_frame2_0___i166_LC_3_24_6  (
            .in0(N__36556),
            .in1(N__32256),
            .in2(_gnd_net_),
            .in3(N__25175),
            .lcout(\c0.data_out_frame2_20_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50292),
            .ce(N__32771),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i157_LC_3_24_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i157_LC_3_24_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i157_LC_3_24_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_out_frame2_0___i157_LC_3_24_7  (
            .in0(N__28808),
            .in1(N__29197),
            .in2(_gnd_net_),
            .in3(N__24316),
            .lcout(\c0.data_out_frame2_19_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50292),
            .ce(N__32771),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i99_LC_3_25_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i99_LC_3_25_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i99_LC_3_25_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_out_frame2_0___i99_LC_3_25_0  (
            .in0(N__34108),
            .in1(N__32607),
            .in2(_gnd_net_),
            .in3(N__19012),
            .lcout(data_out_frame2_12_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50300),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i120_LC_3_25_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i120_LC_3_25_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i120_LC_3_25_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i120_LC_3_25_1  (
            .in0(N__32601),
            .in1(N__36003),
            .in2(_gnd_net_),
            .in3(N__19444),
            .lcout(data_out_frame2_14_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50300),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i106_LC_3_25_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i106_LC_3_25_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i106_LC_3_25_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_out_frame2_0___i106_LC_3_25_2  (
            .in0(N__18994),
            .in1(N__32605),
            .in2(_gnd_net_),
            .in3(N__35888),
            .lcout(data_out_frame2_13_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50300),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i56_LC_3_25_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i56_LC_3_25_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i56_LC_3_25_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i56_LC_3_25_3  (
            .in0(N__32603),
            .in1(N__36004),
            .in2(_gnd_net_),
            .in3(N__20341),
            .lcout(data_out_frame2_6_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50300),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i126_LC_3_25_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i126_LC_3_25_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i126_LC_3_25_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_out_frame2_0___i126_LC_3_25_4  (
            .in0(N__35601),
            .in1(N__32606),
            .in2(_gnd_net_),
            .in3(N__23641),
            .lcout(data_out_frame2_15_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50300),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i128_LC_3_25_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i128_LC_3_25_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i128_LC_3_25_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i128_LC_3_25_5  (
            .in0(N__32602),
            .in1(N__35467),
            .in2(_gnd_net_),
            .in3(N__19429),
            .lcout(data_out_frame2_15_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50300),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i8_LC_3_25_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i8_LC_3_25_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i8_LC_3_25_6 .LUT_INIT=16'b0000110010101110;
    LogicCell40 \c0.data_out_frame2_0___i8_LC_3_25_6  (
            .in0(N__33149),
            .in1(N__23464),
            .in2(N__33677),
            .in3(N__23877),
            .lcout(\c0.data_out_frame2_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50300),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i98_LC_3_25_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i98_LC_3_25_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i98_LC_3_25_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i98_LC_3_25_7  (
            .in0(N__32604),
            .in1(N__34166),
            .in2(_gnd_net_),
            .in3(N__19153),
            .lcout(data_out_frame2_12_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50300),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i57_LC_3_26_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i57_LC_3_26_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i57_LC_3_26_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i57_LC_3_26_0  (
            .in0(N__34884),
            .in1(N__19135),
            .in2(_gnd_net_),
            .in3(N__32762),
            .lcout(data_out_frame2_7_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50308),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_adj_1038_LC_3_26_1 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_adj_1038_LC_3_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_adj_1038_LC_3_26_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \c0.i1_3_lut_4_lut_adj_1038_LC_3_26_1  (
            .in0(N__33345),
            .in1(N__33230),
            .in2(N__33530),
            .in3(N__23206),
            .lcout(n9606),
            .ltout(n9606_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i86_LC_3_26_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i86_LC_3_26_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i86_LC_3_26_2 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \c0.data_out_frame2_0___i86_LC_3_26_2  (
            .in0(_gnd_net_),
            .in1(N__36104),
            .in2(N__19121),
            .in3(N__19117),
            .lcout(data_out_frame2_10_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50308),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i110_LC_3_26_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i110_LC_3_26_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i110_LC_3_26_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i110_LC_3_26_3  (
            .in0(N__32598),
            .in1(N__36408),
            .in2(_gnd_net_),
            .in3(N__19096),
            .lcout(data_out_frame2_13_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50308),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i73_LC_3_26_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i73_LC_3_26_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i73_LC_3_26_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i73_LC_3_26_4  (
            .in0(N__35950),
            .in1(N__19078),
            .in2(_gnd_net_),
            .in3(N__32763),
            .lcout(data_out_frame2_9_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50308),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i141_LC_3_26_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i141_LC_3_26_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i141_LC_3_26_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \c0.data_out_frame2_0___i141_LC_3_26_5  (
            .in0(N__32599),
            .in1(_gnd_net_),
            .in2(N__35663),
            .in3(N__26200),
            .lcout(data_out_frame2_17_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50308),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i108_LC_3_26_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i108_LC_3_26_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i108_LC_3_26_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i108_LC_3_26_6  (
            .in0(N__35774),
            .in1(N__23329),
            .in2(_gnd_net_),
            .in3(N__32761),
            .lcout(data_out_frame2_13_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50308),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i74_LC_3_26_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i74_LC_3_26_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i74_LC_3_26_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i74_LC_3_26_7  (
            .in0(N__32600),
            .in1(N__35887),
            .in2(_gnd_net_),
            .in3(N__19267),
            .lcout(data_out_frame2_9_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50308),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i50_LC_3_27_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i50_LC_3_27_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i50_LC_3_27_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_out_frame2_0___i50_LC_3_27_0  (
            .in0(N__19228),
            .in1(N__32614),
            .in2(_gnd_net_),
            .in3(N__35355),
            .lcout(data_out_frame2_6_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50316),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i139_LC_3_27_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i139_LC_3_27_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i139_LC_3_27_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i139_LC_3_27_1  (
            .in0(N__32608),
            .in1(N__34757),
            .in2(_gnd_net_),
            .in3(N__19207),
            .lcout(data_out_frame2_17_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50316),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i48_LC_3_27_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i48_LC_3_27_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i48_LC_3_27_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_out_frame2_0___i48_LC_3_27_2  (
            .in0(N__36308),
            .in1(N__32613),
            .in2(_gnd_net_),
            .in3(N__19193),
            .lcout(data_out_frame2_5_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50316),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i67_LC_3_27_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i67_LC_3_27_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i67_LC_3_27_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i67_LC_3_27_3  (
            .in0(N__32611),
            .in1(N__34101),
            .in2(_gnd_net_),
            .in3(N__19372),
            .lcout(data_out_frame2_8_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50316),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i112_LC_3_27_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i112_LC_3_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i112_LC_3_27_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_out_frame2_0___i112_LC_3_27_4  (
            .in0(N__36307),
            .in1(N__32612),
            .in2(_gnd_net_),
            .in3(N__19402),
            .lcout(data_out_frame2_13_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50316),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i54_LC_3_27_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i54_LC_3_27_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i54_LC_3_27_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i54_LC_3_27_5  (
            .in0(N__32610),
            .in1(N__36100),
            .in2(_gnd_net_),
            .in3(N__19174),
            .lcout(data_out_frame2_6_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50316),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i60_LC_3_27_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i60_LC_3_27_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i60_LC_3_27_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_out_frame2_0___i60_LC_3_27_6  (
            .in0(N__35715),
            .in1(N__32615),
            .in2(_gnd_net_),
            .in3(N__19717),
            .lcout(data_out_frame2_7_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50316),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i49_LC_3_27_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i49_LC_3_27_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i49_LC_3_27_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i49_LC_3_27_7  (
            .in0(N__32609),
            .in1(N__35408),
            .in2(_gnd_net_),
            .in3(N__19324),
            .lcout(data_out_frame2_6_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50316),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i58_LC_3_28_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i58_LC_3_28_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i58_LC_3_28_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i58_LC_3_28_0  (
            .in0(N__32715),
            .in1(N__34824),
            .in2(_gnd_net_),
            .in3(N__19309),
            .lcout(data_out_frame2_7_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50325),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i135_LC_3_28_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i135_LC_3_28_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i135_LC_3_28_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i135_LC_3_28_1  (
            .in0(N__35040),
            .in1(N__19291),
            .in2(_gnd_net_),
            .in3(N__32718),
            .lcout(data_out_frame2_16_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50325),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16105_LC_3_28_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16105_LC_3_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16105_LC_3_28_2 .LUT_INIT=16'b1010111111000000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_16105_LC_3_28_2  (
            .in0(N__19276),
            .in1(N__20923),
            .in2(N__31130),
            .in3(N__30759),
            .lcout(\c0.n18588 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i96_LC_3_28_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i96_LC_3_28_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i96_LC_3_28_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i96_LC_3_28_3  (
            .in0(N__35460),
            .in1(N__19277),
            .in2(_gnd_net_),
            .in3(N__32720),
            .lcout(data_out_frame2_11_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50325),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i76_LC_3_28_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i76_LC_3_28_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i76_LC_3_28_4 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \c0.data_out_frame2_0___i76_LC_3_28_4  (
            .in0(N__32716),
            .in1(_gnd_net_),
            .in2(N__23510),
            .in3(N__35770),
            .lcout(data_out_frame2_9_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50325),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i66_LC_3_28_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i66_LC_3_28_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i66_LC_3_28_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i66_LC_3_28_5  (
            .in0(N__34160),
            .in1(N__19252),
            .in2(_gnd_net_),
            .in3(N__32719),
            .lcout(data_out_frame2_8_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50325),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18480_bdd_4_lut_LC_3_28_6 .C_ON=1'b0;
    defparam \c0.n18480_bdd_4_lut_LC_3_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.n18480_bdd_4_lut_LC_3_28_6 .LUT_INIT=16'b1110111001010000;
    LogicCell40 \c0.n18480_bdd_4_lut_LC_3_28_6  (
            .in0(N__31100),
            .in1(N__19268),
            .in2(N__19253),
            .in3(N__23288),
            .lcout(\c0.n17833 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i132_LC_3_28_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i132_LC_3_28_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i132_LC_3_28_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i132_LC_3_28_7  (
            .in0(N__35210),
            .in1(N__25999),
            .in2(_gnd_net_),
            .in3(N__32717),
            .lcout(data_out_frame2_16_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50325),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i75_LC_3_29_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i75_LC_3_29_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i75_LC_3_29_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i75_LC_3_29_0  (
            .in0(N__35809),
            .in1(N__19388),
            .in2(_gnd_net_),
            .in3(N__32800),
            .lcout(data_out_frame2_9_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50334),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i153_LC_3_29_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i153_LC_3_29_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i153_LC_3_29_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_out_frame2_0___i153_LC_3_29_1  (
            .in0(N__32798),
            .in1(N__19474),
            .in2(_gnd_net_),
            .in3(N__25831),
            .lcout(data_out_frame2_19_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50334),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_i0_LC_3_29_2 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_i0_LC_3_29_2 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_SM_Main_i0_LC_3_29_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \c0.rx.r_SM_Main_i0_LC_3_29_2  (
            .in0(_gnd_net_),
            .in1(N__39778),
            .in2(_gnd_net_),
            .in3(N__30182),
            .lcout(\c0.rx.r_SM_Main_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50334),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i152_LC_3_29_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i152_LC_3_29_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i152_LC_3_29_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i152_LC_3_29_3  (
            .in0(N__32797),
            .in1(N__34956),
            .in2(_gnd_net_),
            .in3(N__21233),
            .lcout(data_out_frame2_18_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50334),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i104_LC_3_29_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i104_LC_3_29_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i104_LC_3_29_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_out_frame2_0___i104_LC_3_29_4  (
            .in0(N__19415),
            .in1(N__34955),
            .in2(_gnd_net_),
            .in3(N__32799),
            .lcout(data_out_frame2_12_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50334),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_0_i22_4_lut_LC_3_29_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_0_i22_4_lut_LC_3_29_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_0_i22_4_lut_LC_3_29_5 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_0_i22_4_lut_LC_3_29_5  (
            .in0(N__26834),
            .in1(N__19460),
            .in2(N__20879),
            .in3(N__26905),
            .lcout(\c0.n22_adj_2510 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16096_LC_3_29_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16096_LC_3_29_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16096_LC_3_29_6 .LUT_INIT=16'b1110110000101100;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_16096_LC_3_29_6  (
            .in0(N__19445),
            .in1(N__30754),
            .in2(N__31143),
            .in3(N__19430),
            .lcout(),
            .ltout(\c0.n18582_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18582_bdd_4_lut_LC_3_29_7 .C_ON=1'b0;
    defparam \c0.n18582_bdd_4_lut_LC_3_29_7 .SEQ_MODE=4'b0000;
    defparam \c0.n18582_bdd_4_lut_LC_3_29_7 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n18582_bdd_4_lut_LC_3_29_7  (
            .in0(N__31128),
            .in1(N__19414),
            .in2(N__19406),
            .in3(N__19403),
            .lcout(\c0.n17788 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18504_bdd_4_lut_LC_3_30_0 .C_ON=1'b0;
    defparam \c0.n18504_bdd_4_lut_LC_3_30_0 .SEQ_MODE=4'b0000;
    defparam \c0.n18504_bdd_4_lut_LC_3_30_0 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \c0.n18504_bdd_4_lut_LC_3_30_0  (
            .in0(N__19387),
            .in1(N__31129),
            .in2(N__19376),
            .in3(N__19358),
            .lcout(\c0.n17824 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Bit_Index_0__bdd_4_lut_LC_3_30_1 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_0__bdd_4_lut_LC_3_30_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_Bit_Index_0__bdd_4_lut_LC_3_30_1 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \c0.tx2.r_Bit_Index_0__bdd_4_lut_LC_3_30_1  (
            .in0(N__26118),
            .in1(N__26051),
            .in2(N__26180),
            .in3(N__19340),
            .lcout(),
            .ltout(\c0.tx2.n18612_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.n18612_bdd_4_lut_LC_3_30_2 .C_ON=1'b0;
    defparam \c0.tx2.n18612_bdd_4_lut_LC_3_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.n18612_bdd_4_lut_LC_3_30_2 .LUT_INIT=16'b1111000011001010;
    LogicCell40 \c0.tx2.n18612_bdd_4_lut_LC_3_30_2  (
            .in0(N__19592),
            .in1(N__19580),
            .in2(N__19571),
            .in3(N__26168),
            .lcout(\c0.tx2.n18615 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Bit_Index_0__bdd_4_lut_16115_LC_3_30_4 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_0__bdd_4_lut_16115_LC_3_30_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_Bit_Index_0__bdd_4_lut_16115_LC_3_30_4 .LUT_INIT=16'b1010110011110000;
    LogicCell40 \c0.tx2.r_Bit_Index_0__bdd_4_lut_16115_LC_3_30_4  (
            .in0(N__21005),
            .in1(N__19562),
            .in2(N__26129),
            .in3(N__26167),
            .lcout(\c0.tx2.n18450 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Bit_Index_i0_LC_3_30_5 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_i0_LC_3_30_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Bit_Index_i0_LC_3_30_5 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \c0.tx2.r_Bit_Index_i0_LC_3_30_5  (
            .in0(N__26119),
            .in1(N__25935),
            .in2(_gnd_net_),
            .in3(N__25905),
            .lcout(r_Bit_Index_0_adj_2637),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50344),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Bit_Index_i1_LC_3_30_6 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_i1_LC_3_30_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Bit_Index_i1_LC_3_30_6 .LUT_INIT=16'b0001010001000100;
    LogicCell40 \c0.tx2.r_Bit_Index_i1_LC_3_30_6  (
            .in0(N__25906),
            .in1(N__26169),
            .in2(N__25942),
            .in3(N__26120),
            .lcout(r_Bit_Index_1_adj_2636),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50344),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i143_LC_3_30_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i143_LC_3_30_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i143_LC_3_30_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_out_frame2_0___i143_LC_3_30_7  (
            .in0(N__19556),
            .in1(N__35523),
            .in2(_gnd_net_),
            .in3(N__32809),
            .lcout(data_out_frame2_17_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50344),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_3_i6_4_lut_LC_3_31_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_3_i6_4_lut_LC_3_31_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_3_i6_4_lut_LC_3_31_0 .LUT_INIT=16'b1100110010100000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_3_i6_4_lut_LC_3_31_0  (
            .in0(N__30773),
            .in1(N__19703),
            .in2(N__19730),
            .in3(N__31043),
            .lcout(\c0.n6_adj_2432 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i11_3_lut_LC_3_31_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i11_3_lut_LC_3_31_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i11_3_lut_LC_3_31_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_4_i11_3_lut_LC_3_31_1  (
            .in0(N__20981),
            .in1(N__19544),
            .in2(_gnd_net_),
            .in3(N__30771),
            .lcout(),
            .ltout(\c0.n11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_1__bdd_4_lut_15987_LC_3_31_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_1__bdd_4_lut_15987_LC_3_31_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_1__bdd_4_lut_15987_LC_3_31_2 .LUT_INIT=16'b1101100010101010;
    LogicCell40 \c0.byte_transmit_counter2_1__bdd_4_lut_15987_LC_3_31_2  (
            .in0(N__31035),
            .in1(N__19526),
            .in2(N__19514),
            .in3(N__26833),
            .lcout(\c0.n18444 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.n18450_bdd_4_lut_LC_3_31_3 .C_ON=1'b0;
    defparam \c0.tx2.n18450_bdd_4_lut_LC_3_31_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.n18450_bdd_4_lut_LC_3_31_3 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \c0.tx2.n18450_bdd_4_lut_LC_3_31_3  (
            .in0(N__19511),
            .in1(N__26170),
            .in2(N__26432),
            .in3(N__19496),
            .lcout(\c0.tx2.n18453 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i44_LC_3_31_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i44_LC_3_31_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i44_LC_3_31_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_out_frame2_0___i44_LC_3_31_4  (
            .in0(N__19729),
            .in1(N__35769),
            .in2(_gnd_net_),
            .in3(N__32813),
            .lcout(data_out_frame2_5_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50354),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_3_i5_3_lut_LC_3_31_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_3_i5_3_lut_LC_3_31_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_3_i5_3_lut_LC_3_31_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_3_i5_3_lut_LC_3_31_7  (
            .in0(N__19718),
            .in1(N__20777),
            .in2(_gnd_net_),
            .in3(N__30772),
            .lcout(\c0.n5_adj_2509 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_adj_1100_LC_3_32_0 .C_ON=1'b0;
    defparam \c0.i1_3_lut_adj_1100_LC_3_32_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_adj_1100_LC_3_32_0 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \c0.i1_3_lut_adj_1100_LC_3_32_0  (
            .in0(N__26668),
            .in1(N__26519),
            .in2(_gnd_net_),
            .in3(N__26785),
            .lcout(),
            .ltout(\c0.n18_adj_2544_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1102_LC_3_32_1 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1102_LC_3_32_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1102_LC_3_32_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i3_4_lut_adj_1102_LC_3_32_1  (
            .in0(N__19697),
            .in1(N__19673),
            .in2(N__19649),
            .in3(N__19646),
            .lcout(\c0.n19_adj_2540 ),
            .ltout(\c0.n19_adj_2540_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15867_2_lut_LC_3_32_2 .C_ON=1'b0;
    defparam \c0.i15867_2_lut_LC_3_32_2 .SEQ_MODE=4'b0000;
    defparam \c0.i15867_2_lut_LC_3_32_2 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \c0.i15867_2_lut_LC_3_32_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19622),
            .in3(N__19822),
            .lcout(\c0.tx2_transmit_N_2287 ),
            .ltout(\c0.tx2_transmit_N_2287_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_transmit_3602_LC_3_32_3 .C_ON=1'b0;
    defparam \c0.tx2_transmit_3602_LC_3_32_3 .SEQ_MODE=4'b1001;
    defparam \c0.tx2_transmit_3602_LC_3_32_3 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \c0.tx2_transmit_3602_LC_3_32_3  (
            .in0(N__33251),
            .in1(N__33322),
            .in2(N__19607),
            .in3(N__33518),
            .lcout(\c0.r_SM_Main_2_N_2326_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50365),
            .ce(),
            .sr(N__33633));
    defparam \c0.i3_3_lut_adj_1105_LC_3_32_4 .C_ON=1'b0;
    defparam \c0.i3_3_lut_adj_1105_LC_3_32_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_3_lut_adj_1105_LC_3_32_4 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \c0.i3_3_lut_adj_1105_LC_3_32_4  (
            .in0(N__33517),
            .in1(N__33249),
            .in2(_gnd_net_),
            .in3(N__33320),
            .lcout(),
            .ltout(\c0.n67_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1071_LC_3_32_5 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1071_LC_3_32_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1071_LC_3_32_5 .LUT_INIT=16'b1111111110110000;
    LogicCell40 \c0.i1_4_lut_adj_1071_LC_3_32_5  (
            .in0(N__19823),
            .in1(N__19604),
            .in2(N__19595),
            .in3(N__32643),
            .lcout(\c0.n4_adj_2480 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i11145_2_lut_LC_3_32_6 .C_ON=1'b0;
    defparam \c0.tx2.i11145_2_lut_LC_3_32_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i11145_2_lut_LC_3_32_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.tx2.i11145_2_lut_LC_3_32_6  (
            .in0(_gnd_net_),
            .in1(N__21500),
            .in2(_gnd_net_),
            .in3(N__21523),
            .lcout(\c0.n13530 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15907_2_lut_3_lut_LC_3_32_7 .C_ON=1'b0;
    defparam \c0.i15907_2_lut_3_lut_LC_3_32_7 .SEQ_MODE=4'b0000;
    defparam \c0.i15907_2_lut_3_lut_LC_3_32_7 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \c0.i15907_2_lut_3_lut_LC_3_32_7  (
            .in0(N__33250),
            .in1(N__33321),
            .in2(_gnd_net_),
            .in3(N__33516),
            .lcout(\c0.n142 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1018_LC_4_17_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1018_LC_4_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1018_LC_4_17_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1018_LC_4_17_0  (
            .in0(N__20290),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25273),
            .lcout(\c0.n8062 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_938_LC_4_17_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_938_LC_4_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_938_LC_4_17_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_938_LC_4_17_1  (
            .in0(_gnd_net_),
            .in1(N__19814),
            .in2(_gnd_net_),
            .in3(N__28716),
            .lcout(\c0.n17529 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_847_LC_4_17_2 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_847_LC_4_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_847_LC_4_17_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_847_LC_4_17_2  (
            .in0(N__29134),
            .in1(N__19922),
            .in2(N__20135),
            .in3(N__19796),
            .lcout(),
            .ltout(\c0.n10_adj_2428_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_848_LC_4_17_3 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_848_LC_4_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_848_LC_4_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i5_3_lut_adj_848_LC_4_17_3  (
            .in0(_gnd_net_),
            .in1(N__25433),
            .in2(N__19787),
            .in3(N__20289),
            .lcout(\c0.n9324 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1050_LC_4_17_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1050_LC_4_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1050_LC_4_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1050_LC_4_17_4  (
            .in0(N__21684),
            .in1(N__20527),
            .in2(_gnd_net_),
            .in3(N__19748),
            .lcout(\c0.n17442 ),
            .ltout(\c0.n17442_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_948_LC_4_17_5 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_948_LC_4_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_948_LC_4_17_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_948_LC_4_17_5  (
            .in0(N__29089),
            .in1(N__19775),
            .in2(N__19766),
            .in3(N__19763),
            .lcout(\c0.n8674 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i10_LC_4_17_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i10_LC_4_17_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i10_LC_4_17_6 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \c0.data_in_frame_0___i10_LC_4_17_6  (
            .in0(N__24256),
            .in1(N__31382),
            .in2(N__28723),
            .in3(N__31937),
            .lcout(data_in_frame_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50256),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i33_LC_4_17_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i33_LC_4_17_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i33_LC_4_17_7 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \c0.data_in_frame_0___i33_LC_4_17_7  (
            .in0(N__19749),
            .in1(N__27865),
            .in2(N__31978),
            .in3(N__24257),
            .lcout(\c0.data_in_frame_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50256),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1079_LC_4_18_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1079_LC_4_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1079_LC_4_18_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1079_LC_4_18_0  (
            .in0(N__28714),
            .in1(N__20093),
            .in2(N__22041),
            .in3(N__19851),
            .lcout(\c0.n8874 ),
            .ltout(\c0.n8874_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_963_LC_4_18_1 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_963_LC_4_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_963_LC_4_18_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_963_LC_4_18_1  (
            .in0(N__19902),
            .in1(N__19967),
            .in2(N__19940),
            .in3(N__19936),
            .lcout(\c0.n9368 ),
            .ltout(\c0.n9368_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_1093_LC_4_18_2 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_1093_LC_4_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_1093_LC_4_18_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_1093_LC_4_18_2  (
            .in0(N__21906),
            .in1(N__21606),
            .in2(N__19925),
            .in3(N__19918),
            .lcout(\c0.n12_adj_2542 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_2_lut_3_lut_4_lut_LC_4_18_3 .C_ON=1'b0;
    defparam \c0.i14_2_lut_3_lut_4_lut_LC_4_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i14_2_lut_3_lut_4_lut_LC_4_18_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i14_2_lut_3_lut_4_lut_LC_4_18_3  (
            .in0(N__22595),
            .in1(N__22635),
            .in2(N__28261),
            .in3(N__22542),
            .lcout(\c0.n9306 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1031_LC_4_18_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1031_LC_4_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1031_LC_4_18_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1031_LC_4_18_4  (
            .in0(_gnd_net_),
            .in1(N__22138),
            .in2(_gnd_net_),
            .in3(N__19903),
            .lcout(\c0.n17632 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_865_LC_4_18_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_865_LC_4_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_865_LC_4_18_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_865_LC_4_18_5  (
            .in0(N__20094),
            .in1(N__22033),
            .in2(_gnd_net_),
            .in3(N__28715),
            .lcout(\c0.n17485 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i40_LC_4_18_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i40_LC_4_18_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i40_LC_4_18_6 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \c0.data_in_frame_0___i40_LC_4_18_6  (
            .in0(N__22543),
            .in1(N__24258),
            .in2(N__27245),
            .in3(N__31877),
            .lcout(\c0.data_in_frame_4_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50264),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i26_LC_4_19_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i26_LC_4_19_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i26_LC_4_19_0 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \c0.data_in_frame_0___i26_LC_4_19_0  (
            .in0(N__24237),
            .in1(N__27689),
            .in2(N__19858),
            .in3(N__31994),
            .lcout(\c0.data_in_frame_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50269),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_884_LC_4_19_1 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_884_LC_4_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_884_LC_4_19_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_884_LC_4_19_1  (
            .in0(N__19832),
            .in1(N__21553),
            .in2(N__24764),
            .in3(N__22183),
            .lcout(),
            .ltout(\c0.n12_adj_2449_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_LC_4_19_2 .C_ON=1'b0;
    defparam \c0.i8_4_lut_LC_4_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_LC_4_19_2 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \c0.i8_4_lut_LC_4_19_2  (
            .in0(N__24838),
            .in1(N__22973),
            .in2(N__20189),
            .in3(N__20182),
            .lcout(),
            .ltout(\c0.n24_adj_2454_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_LC_4_19_3 .C_ON=1'b0;
    defparam \c0.i14_4_lut_LC_4_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_LC_4_19_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i14_4_lut_LC_4_19_3  (
            .in0(N__22358),
            .in1(N__20159),
            .in2(N__20147),
            .in3(N__20003),
            .lcout(\c0.n30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i73_LC_4_19_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i73_LC_4_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i73_LC_4_19_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.data_in_frame_0___i73_LC_4_19_4  (
            .in0(_gnd_net_),
            .in1(N__29351),
            .in2(_gnd_net_),
            .in3(N__31993),
            .lcout(\c0.data_in_frame_9_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50269),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i44_LC_4_19_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i44_LC_4_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i44_LC_4_19_6 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \c0.data_in_frame_0___i44_LC_4_19_6  (
            .in0(N__24238),
            .in1(N__20122),
            .in2(N__23698),
            .in3(N__31992),
            .lcout(data_in_frame_5_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50269),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i24_LC_4_19_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i24_LC_4_19_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i24_LC_4_19_7 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \c0.data_in_frame_0___i24_LC_4_19_7  (
            .in0(N__20098),
            .in1(N__27284),
            .in2(N__31997),
            .in3(N__24239),
            .lcout(\c0.data_in_frame_2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50269),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3917_3_lut_4_lut_LC_4_20_0 .C_ON=1'b0;
    defparam \c0.i3917_3_lut_4_lut_LC_4_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3917_3_lut_4_lut_LC_4_20_0 .LUT_INIT=16'b1010101011100010;
    LogicCell40 \c0.i3917_3_lut_4_lut_LC_4_20_0  (
            .in0(N__20075),
            .in1(N__34659),
            .in2(N__32161),
            .in3(N__28045),
            .lcout(n2584),
            .ltout(n2584_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_901_LC_4_20_1 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_901_LC_4_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_901_LC_4_20_1 .LUT_INIT=16'b1101011111101011;
    LogicCell40 \c0.i5_4_lut_adj_901_LC_4_20_1  (
            .in0(N__20021),
            .in1(N__22783),
            .in2(N__20006),
            .in3(N__22273),
            .lcout(\c0.n21_adj_2465 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i68_LC_4_20_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i68_LC_4_20_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i68_LC_4_20_3 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \c0.data_in_frame_0___i68_LC_4_20_3  (
            .in0(N__25555),
            .in1(N__31798),
            .in2(N__29747),
            .in3(N__20265),
            .lcout(data_in_frame_8_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50276),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i66_LC_4_20_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i66_LC_4_20_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i66_LC_4_20_4 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \c0.data_in_frame_0___i66_LC_4_20_4  (
            .in0(N__31797),
            .in1(N__37042),
            .in2(N__20274),
            .in3(N__22925),
            .lcout(data_in_frame_8_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50276),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i72_LC_4_20_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i72_LC_4_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i72_LC_4_20_5 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \c0.data_in_frame_0___i72_LC_4_20_5  (
            .in0(N__20375),
            .in1(N__31799),
            .in2(N__29807),
            .in3(N__20266),
            .lcout(data_in_frame_8_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50276),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i16_LC_4_20_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i16_LC_4_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i16_LC_4_20_6 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \c0.data_in_frame_0___i16_LC_4_20_6  (
            .in0(N__25432),
            .in1(N__27041),
            .in2(N__31921),
            .in3(N__24216),
            .lcout(\c0.data_in_frame_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50276),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i55_LC_4_20_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i55_LC_4_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i55_LC_4_20_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.data_in_frame_0___i55_LC_4_20_7  (
            .in0(_gnd_net_),
            .in1(N__22375),
            .in2(_gnd_net_),
            .in3(N__31803),
            .lcout(\c0.data_in_frame_6_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50276),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_909_LC_4_21_0 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_909_LC_4_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_909_LC_4_21_0 .LUT_INIT=16'b1111011001101111;
    LogicCell40 \c0.i2_4_lut_adj_909_LC_4_21_0  (
            .in0(N__21928),
            .in1(N__27942),
            .in2(N__20237),
            .in3(N__22201),
            .lcout(\c0.n18_adj_2468 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i60_LC_4_21_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i60_LC_4_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i60_LC_4_21_1 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \c0.data_in_frame_0___i60_LC_4_21_1  (
            .in0(N__22202),
            .in1(_gnd_net_),
            .in2(N__31924),
            .in3(_gnd_net_),
            .lcout(\c0.data_in_frame_7_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50282),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_910_LC_4_21_2 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_910_LC_4_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_910_LC_4_21_2 .LUT_INIT=16'b1111111111011110;
    LogicCell40 \c0.i10_4_lut_adj_910_LC_4_21_2  (
            .in0(N__22345),
            .in1(N__23753),
            .in2(N__20225),
            .in3(N__20312),
            .lcout(),
            .ltout(\c0.n26_adj_2469_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_adj_916_LC_4_21_3 .C_ON=1'b0;
    defparam \c0.i15_4_lut_adj_916_LC_4_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_adj_916_LC_4_21_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i15_4_lut_adj_916_LC_4_21_3  (
            .in0(N__20207),
            .in1(N__22718),
            .in2(N__20201),
            .in3(N__20198),
            .lcout(\c0.n1_adj_2443 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i87_LC_4_21_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i87_LC_4_21_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i87_LC_4_21_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \c0.data_in_frame_0___i87_LC_4_21_4  (
            .in0(_gnd_net_),
            .in1(N__31824),
            .in2(_gnd_net_),
            .in3(N__29450),
            .lcout(data_in_frame_10_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50282),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i85_LC_4_21_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i85_LC_4_21_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i85_LC_4_21_5 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \c0.data_in_frame_0___i85_LC_4_21_5  (
            .in0(N__31829),
            .in1(N__28658),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.data_in_frame_10_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50282),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i80_LC_4_21_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i80_LC_4_21_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i80_LC_4_21_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \c0.data_in_frame_0___i80_LC_4_21_6  (
            .in0(_gnd_net_),
            .in1(N__31823),
            .in2(_gnd_net_),
            .in3(N__25220),
            .lcout(\c0.data_in_frame_9_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50282),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i79_LC_4_21_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i79_LC_4_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i79_LC_4_21_7 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \c0.data_in_frame_0___i79_LC_4_21_7  (
            .in0(N__31828),
            .in1(N__28894),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(data_in_frame_9_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50282),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i9_LC_4_22_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i9_LC_4_22_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i9_LC_4_22_0 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \c0.data_in_frame_0___i9_LC_4_22_0  (
            .in0(N__24251),
            .in1(N__24014),
            .in2(N__22668),
            .in3(N__31849),
            .lcout(\c0.data_in_frame_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50287),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_7_i5_3_lut_LC_4_22_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_7_i5_3_lut_LC_4_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_7_i5_3_lut_LC_4_22_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_7_i5_3_lut_LC_4_22_1  (
            .in0(N__30674),
            .in1(N__32285),
            .in2(_gnd_net_),
            .in3(N__20345),
            .lcout(\c0.n5_adj_2501 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i34_LC_4_22_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i34_LC_4_22_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i34_LC_4_22_2 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \c0.data_in_frame_0___i34_LC_4_22_2  (
            .in0(N__24250),
            .in1(N__21683),
            .in2(N__38513),
            .in3(N__31848),
            .lcout(\c0.data_in_frame_4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50287),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_887_LC_4_22_3 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_887_LC_4_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_887_LC_4_22_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i5_3_lut_adj_887_LC_4_22_3  (
            .in0(N__24523),
            .in1(_gnd_net_),
            .in2(N__20599),
            .in3(N__22310),
            .lcout(\c0.n17534 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i76_LC_4_22_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i76_LC_4_22_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i76_LC_4_22_4 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \c0.data_in_frame_0___i76_LC_4_22_4  (
            .in0(N__23087),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31847),
            .lcout(\c0.data_in_frame_9_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50287),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i31_LC_4_22_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i31_LC_4_22_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i31_LC_4_22_5 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \c0.data_in_frame_0___i31_LC_4_22_5  (
            .in0(N__29088),
            .in1(N__28190),
            .in2(N__31927),
            .in3(N__24252),
            .lcout(\c0.data_in_frame_3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50287),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_978_LC_4_22_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_978_LC_4_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_978_LC_4_22_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_978_LC_4_22_6  (
            .in0(N__28565),
            .in1(N__25270),
            .in2(_gnd_net_),
            .in3(N__20305),
            .lcout(\c0.n17591 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i37_LC_4_22_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i37_LC_4_22_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i37_LC_4_22_7 .LUT_INIT=16'b0000110000001010;
    LogicCell40 \c0.data_in_frame_0___i37_LC_4_22_7  (
            .in0(N__27371),
            .in1(N__21829),
            .in2(N__31928),
            .in3(N__24253),
            .lcout(\c0.data_in_frame_4_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50287),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1045_LC_4_23_0 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1045_LC_4_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1045_LC_4_23_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1045_LC_4_23_0  (
            .in0(N__20491),
            .in1(N__20621),
            .in2(N__25272),
            .in3(N__24995),
            .lcout(\c0.n17470 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_842_LC_4_23_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_842_LC_4_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_842_LC_4_23_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_842_LC_4_23_1  (
            .in0(_gnd_net_),
            .in1(N__22706),
            .in2(_gnd_net_),
            .in3(N__20376),
            .lcout(n9148),
            .ltout(n9148_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_3_lut_4_lut_LC_4_23_2.C_ON=1'b0;
    defparam i2_3_lut_4_lut_LC_4_23_2.SEQ_MODE=4'b0000;
    defparam i2_3_lut_4_lut_LC_4_23_2.LUT_INIT=16'b0110100110010110;
    LogicCell40 i2_3_lut_4_lut_LC_4_23_2 (
            .in0(N__25021),
            .in1(N__21929),
            .in2(N__20573),
            .in3(N__25582),
            .lcout(n17585),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i45_LC_4_23_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i45_LC_4_23_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i45_LC_4_23_3 .LUT_INIT=16'b0000000011011000;
    LogicCell40 \c0.data_in_frame_0___i45_LC_4_23_3  (
            .in0(N__24255),
            .in1(N__25263),
            .in2(N__27407),
            .in3(N__31892),
            .lcout(data_in_frame_5_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50293),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1111_LC_4_23_4 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1111_LC_4_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1111_LC_4_23_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1111_LC_4_23_4  (
            .in0(N__20566),
            .in1(N__20513),
            .in2(N__25271),
            .in3(N__20537),
            .lcout(\c0.n17605 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i19_LC_4_23_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i19_LC_4_23_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i19_LC_4_23_5 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \c0.data_in_frame_0___i19_LC_4_23_5  (
            .in0(N__24254),
            .in1(N__24383),
            .in2(N__20523),
            .in3(N__31893),
            .lcout(\c0.data_in_frame_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50293),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1036_LC_4_23_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1036_LC_4_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1036_LC_4_23_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1036_LC_4_23_6  (
            .in0(N__20492),
            .in1(N__20462),
            .in2(_gnd_net_),
            .in3(N__20441),
            .lcout(\c0.n8751 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i77_LC_4_23_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i77_LC_4_23_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i77_LC_4_23_7 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \c0.data_out_frame2_0___i77_LC_4_23_7  (
            .in0(N__31219),
            .in1(_gnd_net_),
            .in2(N__36470),
            .in3(N__32678),
            .lcout(data_out_frame2_9_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50293),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1127_LC_4_24_0 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1127_LC_4_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1127_LC_4_24_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_1127_LC_4_24_0  (
            .in0(N__23024),
            .in1(N__20401),
            .in2(N__20381),
            .in3(N__20735),
            .lcout(\c0.n17647 ),
            .ltout(\c0.n17647_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_854_LC_4_24_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_854_LC_4_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_854_LC_4_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i2_3_lut_adj_854_LC_4_24_1  (
            .in0(_gnd_net_),
            .in1(N__28530),
            .in2(N__20738),
            .in3(N__24416),
            .lcout(\c0.n17648 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_1125_LC_4_24_2 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_1125_LC_4_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_1125_LC_4_24_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_1125_LC_4_24_2  (
            .in0(N__24693),
            .in1(N__20648),
            .in2(N__22405),
            .in3(N__24499),
            .lcout(\c0.n12_adj_2549 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i70_LC_4_24_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i70_LC_4_24_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i70_LC_4_24_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i70_LC_4_24_3  (
            .in0(N__45385),
            .in1(N__20712),
            .in2(_gnd_net_),
            .in3(N__32909),
            .lcout(data_in_8_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50301),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1035_LC_4_24_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1035_LC_4_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1035_LC_4_24_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1035_LC_4_24_4  (
            .in0(N__21976),
            .in1(N__22511),
            .in2(N__20696),
            .in3(N__20669),
            .lcout(\c0.n9345 ),
            .ltout(\c0.n9345_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_906_LC_4_24_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_906_LC_4_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_906_LC_4_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_906_LC_4_24_5  (
            .in0(_gnd_net_),
            .in1(N__28342),
            .in2(N__20642),
            .in3(N__24694),
            .lcout(\c0.n17532 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_LC_4_25_0 .C_ON=1'b0;
    defparam \c0.i4_4_lut_LC_4_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_LC_4_25_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_LC_4_25_0  (
            .in0(N__25193),
            .in1(N__32983),
            .in2(N__20905),
            .in3(N__32064),
            .lcout(),
            .ltout(\c0.n10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i160_LC_4_25_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i160_LC_4_25_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i160_LC_4_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_out_frame2_0___i160_LC_4_25_1  (
            .in0(_gnd_net_),
            .in1(N__23099),
            .in2(N__20639),
            .in3(N__21073),
            .lcout(\c0.data_out_frame2_19_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50309),
            .ce(N__32828),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i167_LC_4_25_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i167_LC_4_25_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i167_LC_4_25_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.data_out_frame2_0___i167_LC_4_25_2  (
            .in0(N__21074),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29506),
            .lcout(\c0.data_out_frame2_20_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50309),
            .ce(N__32828),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_837_LC_4_25_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_837_LC_4_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_837_LC_4_25_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_837_LC_4_25_3  (
            .in0(N__24319),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29389),
            .lcout(\c0.n8995 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i161_LC_4_25_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i161_LC_4_25_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i161_LC_4_25_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_frame2_0___i161_LC_4_25_4  (
            .in0(N__20912),
            .in1(N__32214),
            .in2(N__20906),
            .in3(N__20891),
            .lcout(\c0.data_out_frame2_20_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50309),
            .ce(N__32828),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_975_LC_4_25_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_975_LC_4_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_975_LC_4_25_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_975_LC_4_25_5  (
            .in0(N__24320),
            .in1(N__28693),
            .in2(_gnd_net_),
            .in3(N__29390),
            .lcout(),
            .ltout(\c0.n6_adj_2502_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i163_LC_4_25_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i163_LC_4_25_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i163_LC_4_25_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_frame2_0___i163_LC_4_25_6  (
            .in0(N__23528),
            .in1(N__29279),
            .in2(N__20864),
            .in3(N__28850),
            .lcout(\c0.data_out_frame2_20_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50309),
            .ce(N__32828),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i158_LC_4_25_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i158_LC_4_25_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i158_LC_4_25_7 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_frame2_0___i158_LC_4_25_7  (
            .in0(N__23527),
            .in1(N__29391),
            .in2(N__36806),
            .in3(N__23126),
            .lcout(\c0.data_out_frame2_19_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50309),
            .ce(N__32828),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i113_LC_4_26_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i113_LC_4_26_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i113_LC_4_26_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_out_frame2_0___i113_LC_4_26_0  (
            .in0(N__35406),
            .in1(N__32751),
            .in2(_gnd_net_),
            .in3(N__20830),
            .lcout(data_out_frame2_14_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50317),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i147_LC_4_26_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i147_LC_4_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i147_LC_4_26_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i147_LC_4_26_1  (
            .in0(N__32747),
            .in1(N__34100),
            .in2(_gnd_net_),
            .in3(N__20812),
            .lcout(data_out_frame2_18_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50317),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i47_LC_4_26_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i47_LC_4_26_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i47_LC_4_26_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_out_frame2_0___i47_LC_4_26_2  (
            .in0(N__36356),
            .in1(N__32752),
            .in2(_gnd_net_),
            .in3(N__20791),
            .lcout(data_out_frame2_5_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50317),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i52_LC_4_26_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i52_LC_4_26_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i52_LC_4_26_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i52_LC_4_26_3  (
            .in0(N__32748),
            .in1(N__35261),
            .in2(_gnd_net_),
            .in3(N__20773),
            .lcout(data_out_frame2_6_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50317),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i103_LC_4_26_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i103_LC_4_26_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i103_LC_4_26_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_out_frame2_0___i103_LC_4_26_4  (
            .in0(N__35041),
            .in1(N__32750),
            .in2(_gnd_net_),
            .in3(N__20752),
            .lcout(data_out_frame2_12_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50317),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i93_LC_4_26_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i93_LC_4_26_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i93_LC_4_26_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i93_LC_4_26_5  (
            .in0(N__32749),
            .in1(N__35658),
            .in2(_gnd_net_),
            .in3(N__25670),
            .lcout(data_out_frame2_11_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50317),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i82_LC_4_26_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i82_LC_4_26_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i82_LC_4_26_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_out_frame2_0___i82_LC_4_26_6  (
            .in0(N__35357),
            .in1(N__32753),
            .in2(_gnd_net_),
            .in3(N__23300),
            .lcout(data_out_frame2_10_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50317),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i111_LC_4_26_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i111_LC_4_26_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i111_LC_4_26_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i111_LC_4_26_7  (
            .in0(N__32746),
            .in1(N__36355),
            .in2(_gnd_net_),
            .in3(N__20959),
            .lcout(data_out_frame2_13_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50317),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i65_LC_4_27_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i65_LC_4_27_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i65_LC_4_27_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i65_LC_4_27_0  (
            .in0(N__32633),
            .in1(N__34212),
            .in2(_gnd_net_),
            .in3(N__20938),
            .lcout(data_out_frame2_8_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50326),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i148_LC_4_27_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i148_LC_4_27_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i148_LC_4_27_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i148_LC_4_27_1  (
            .in0(N__35209),
            .in1(N__26035),
            .in2(_gnd_net_),
            .in3(N__32638),
            .lcout(data_out_frame2_18_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50326),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i144_LC_4_27_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i144_LC_4_27_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i144_LC_4_27_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i144_LC_4_27_2  (
            .in0(N__32632),
            .in1(N__35459),
            .in2(_gnd_net_),
            .in3(N__21205),
            .lcout(data_out_frame2_17_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50326),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i124_LC_4_27_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i124_LC_4_27_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i124_LC_4_27_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i124_LC_4_27_3  (
            .in0(N__35716),
            .in1(N__23363),
            .in2(_gnd_net_),
            .in3(N__32636),
            .lcout(data_out_frame2_15_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50326),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i88_LC_4_27_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i88_LC_4_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i88_LC_4_27_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i88_LC_4_27_4  (
            .in0(N__32634),
            .in1(N__36005),
            .in2(_gnd_net_),
            .in3(N__20924),
            .lcout(data_out_frame2_10_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50326),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i72_LC_4_27_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i72_LC_4_27_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i72_LC_4_27_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i72_LC_4_27_5  (
            .in0(N__34963),
            .in1(N__23419),
            .in2(_gnd_net_),
            .in3(N__32639),
            .lcout(data_out_frame2_8_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50326),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i90_LC_4_27_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i90_LC_4_27_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i90_LC_4_27_6 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \c0.data_out_frame2_0___i90_LC_4_27_6  (
            .in0(N__32635),
            .in1(N__34817),
            .in2(N__23315),
            .in3(_gnd_net_),
            .lcout(data_out_frame2_11_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50326),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i140_LC_4_27_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i140_LC_4_27_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i140_LC_4_27_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i140_LC_4_27_7  (
            .in0(N__35717),
            .in1(N__25978),
            .in2(_gnd_net_),
            .in3(N__32637),
            .lcout(data_out_frame2_17_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50326),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i125_LC_4_28_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i125_LC_4_28_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i125_LC_4_28_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i125_LC_4_28_0  (
            .in0(N__35647),
            .in1(N__20995),
            .in2(_gnd_net_),
            .in3(N__32790),
            .lcout(data_out_frame2_15_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50335),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i39_LC_4_28_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i39_LC_4_28_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i39_LC_4_28_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i39_LC_4_28_1  (
            .in0(N__45292),
            .in1(N__28365),
            .in2(_gnd_net_),
            .in3(N__31270),
            .lcout(\c0.data_in_4_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50335),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i149_LC_4_28_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i149_LC_4_28_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i149_LC_4_28_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i149_LC_4_28_2  (
            .in0(N__35138),
            .in1(N__26260),
            .in2(_gnd_net_),
            .in3(N__32791),
            .lcout(data_out_frame2_18_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50335),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i85_LC_4_28_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i85_LC_4_28_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i85_LC_4_28_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i85_LC_4_28_3  (
            .in0(N__32788),
            .in1(N__36143),
            .in2(_gnd_net_),
            .in3(N__25687),
            .lcout(data_out_frame2_10_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50335),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i80_LC_4_28_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i80_LC_4_28_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i80_LC_4_28_5 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \c0.data_out_frame2_0___i80_LC_4_28_5  (
            .in0(N__32787),
            .in1(N__36306),
            .in2(N__23435),
            .in3(_gnd_net_),
            .lcout(data_out_frame2_9_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50335),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i101_LC_4_28_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i101_LC_4_28_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i101_LC_4_28_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i101_LC_4_28_6  (
            .in0(N__35137),
            .in1(N__20980),
            .in2(_gnd_net_),
            .in3(N__32789),
            .lcout(data_out_frame2_12_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50335),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1096_LC_4_28_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1096_LC_4_28_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1096_LC_4_28_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1096_LC_4_28_7  (
            .in0(N__29392),
            .in1(N__28645),
            .in2(_gnd_net_),
            .in3(N__24318),
            .lcout(\c0.n17504 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_838_LC_4_29_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_838_LC_4_29_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_838_LC_4_29_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_838_LC_4_29_0  (
            .in0(_gnd_net_),
            .in1(N__28974),
            .in2(_gnd_net_),
            .in3(N__28937),
            .lcout(),
            .ltout(\c0.n17535_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i159_LC_4_29_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i159_LC_4_29_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i159_LC_4_29_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_frame2_0___i159_LC_4_29_1  (
            .in0(N__29323),
            .in1(N__21086),
            .in2(N__21104),
            .in3(N__36743),
            .lcout(\c0.data_out_frame2_19_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50345),
            .ce(N__32792),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_852_LC_4_29_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_852_LC_4_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_852_LC_4_29_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_852_LC_4_29_2  (
            .in0(_gnd_net_),
            .in1(N__28694),
            .in2(_gnd_net_),
            .in3(N__32066),
            .lcout(\c0.n9240 ),
            .ltout(\c0.n9240_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1117_LC_4_29_3 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1117_LC_4_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1117_LC_4_29_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1117_LC_4_29_3  (
            .in0(N__21064),
            .in1(N__29393),
            .in2(N__21077),
            .in3(N__29479),
            .lcout(\c0.n10_adj_2470 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1110_LC_4_29_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1110_LC_4_29_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1110_LC_4_29_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1110_LC_4_29_4  (
            .in0(N__32114),
            .in1(N__29257),
            .in2(N__31520),
            .in3(N__25637),
            .lcout(\c0.n9131 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1121_LC_4_29_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1121_LC_4_29_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1121_LC_4_29_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1121_LC_4_29_5  (
            .in0(_gnd_net_),
            .in1(N__36742),
            .in2(_gnd_net_),
            .in3(N__36692),
            .lcout(),
            .ltout(\c0.n17409_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i162_LC_4_29_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i162_LC_4_29_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i162_LC_4_29_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_frame2_0___i162_LC_4_29_6  (
            .in0(N__36632),
            .in1(N__32216),
            .in2(N__21053),
            .in3(N__21050),
            .lcout(\c0.data_out_frame2_20_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50345),
            .ce(N__32792),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i154_LC_4_29_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i154_LC_4_29_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i154_LC_4_29_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_out_frame2_0___i154_LC_4_29_7  (
            .in0(N__32215),
            .in1(N__36631),
            .in2(_gnd_net_),
            .in3(N__28880),
            .lcout(\c0.data_out_frame2_19_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50345),
            .ce(N__32792),
            .sr(_gnd_net_));
    defparam \c0.n18420_bdd_4_lut_LC_4_30_0 .C_ON=1'b0;
    defparam \c0.n18420_bdd_4_lut_LC_4_30_0 .SEQ_MODE=4'b0000;
    defparam \c0.n18420_bdd_4_lut_LC_4_30_0 .LUT_INIT=16'b1110111001010000;
    LogicCell40 \c0.n18420_bdd_4_lut_LC_4_30_0  (
            .in0(N__26673),
            .in1(N__21020),
            .in2(N__23450),
            .in3(N__21173),
            .lcout(),
            .ltout(\c0.n18423_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i7_LC_4_30_1 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i7_LC_4_30_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i7_LC_4_30_1 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \c0.tx2.r_Tx_Data_i7_LC_4_30_1  (
            .in0(N__21188),
            .in1(N__26674),
            .in2(N__21008),
            .in3(N__26520),
            .lcout(\c0.tx2.r_Tx_Data_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50355),
            .ce(N__26417),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16091_LC_4_30_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16091_LC_4_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16091_LC_4_30_2 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_16091_LC_4_30_2  (
            .in0(N__21232),
            .in1(N__31094),
            .in2(N__21221),
            .in3(N__30791),
            .lcout(),
            .ltout(\c0.n18576_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18576_bdd_4_lut_LC_4_30_3 .C_ON=1'b0;
    defparam \c0.n18576_bdd_4_lut_LC_4_30_3 .SEQ_MODE=4'b0000;
    defparam \c0.n18576_bdd_4_lut_LC_4_30_3 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n18576_bdd_4_lut_LC_4_30_3  (
            .in0(N__31095),
            .in1(N__22427),
            .in2(N__21209),
            .in3(N__21206),
            .lcout(),
            .ltout(\c0.n18579_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_7_i22_4_lut_LC_4_30_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_7_i22_4_lut_LC_4_30_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_7_i22_4_lut_LC_4_30_4 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_7_i22_4_lut_LC_4_30_4  (
            .in0(N__26841),
            .in1(N__23171),
            .in2(N__21191),
            .in3(N__26941),
            .lcout(\c0.n22_adj_2520 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15970_LC_4_30_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15970_LC_4_30_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15970_LC_4_30_5 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_15970_LC_4_30_5  (
            .in0(N__23396),
            .in1(N__26672),
            .in2(N__21182),
            .in3(N__26840),
            .lcout(\c0.n18420 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i2_LC_4_31_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i2_LC_4_31_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i2_LC_4_31_0 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \c0.FRAME_MATCHER_state_i2_LC_4_31_0  (
            .in0(N__33491),
            .in1(N__33326),
            .in2(_gnd_net_),
            .in3(N__33265),
            .lcout(\c0.FRAME_MATCHER_state_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50366),
            .ce(),
            .sr(N__21167));
    defparam \c0.rx.i1_2_lut_LC_4_31_1 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_LC_4_31_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_LC_4_31_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.rx.i1_2_lut_LC_4_31_1  (
            .in0(_gnd_net_),
            .in1(N__39656),
            .in2(_gnd_net_),
            .in3(N__39565),
            .lcout(\c0.rx.n79 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i1_2_lut_adj_824_LC_4_31_2 .C_ON=1'b0;
    defparam \c0.tx2.i1_2_lut_adj_824_LC_4_31_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i1_2_lut_adj_824_LC_4_31_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \c0.tx2.i1_2_lut_adj_824_LC_4_31_2  (
            .in0(_gnd_net_),
            .in1(N__21326),
            .in2(_gnd_net_),
            .in3(N__21501),
            .lcout(\c0.tx2.n4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.o_Tx_Serial_I_0_1_lut_LC_4_31_3 .C_ON=1'b0;
    defparam \c0.tx.o_Tx_Serial_I_0_1_lut_LC_4_31_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx.o_Tx_Serial_I_0_1_lut_LC_4_31_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \c0.tx.o_Tx_Serial_I_0_1_lut_LC_4_31_3  (
            .in0(N__37162),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(tx_enable),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.o_Tx_Serial_I_0_1_lut_LC_4_31_4 .C_ON=1'b0;
    defparam \c0.tx2.o_Tx_Serial_I_0_1_lut_LC_4_31_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.o_Tx_Serial_I_0_1_lut_LC_4_31_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \c0.tx2.o_Tx_Serial_I_0_1_lut_LC_4_31_4  (
            .in0(N__21148),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(tx2_enable),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i1_4_lut_LC_4_32_0 .C_ON=1'b0;
    defparam \c0.tx2.i1_4_lut_LC_4_32_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i1_4_lut_LC_4_32_0 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \c0.tx2.i1_4_lut_LC_4_32_0  (
            .in0(N__21288),
            .in1(N__21533),
            .in2(N__21434),
            .in3(N__21512),
            .lcout(),
            .ltout(\c0.tx2.n9568_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Active_47_LC_4_32_1 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Active_47_LC_4_32_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Active_47_LC_4_32_1 .LUT_INIT=16'b0011111100110000;
    LogicCell40 \c0.tx2.r_Tx_Active_47_LC_4_32_1  (
            .in0(_gnd_net_),
            .in1(N__21292),
            .in2(N__21527),
            .in3(N__21524),
            .lcout(\c0.tx2.tx2_active ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50374),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i2_4_lut_adj_823_LC_4_32_2 .C_ON=1'b0;
    defparam \c0.tx2.i2_4_lut_adj_823_LC_4_32_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i2_4_lut_adj_823_LC_4_32_2 .LUT_INIT=16'b0001000100000001;
    LogicCell40 \c0.tx2.i2_4_lut_adj_823_LC_4_32_2  (
            .in0(N__21323),
            .in1(N__21426),
            .in2(N__21295),
            .in3(N__21467),
            .lcout(n9652),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i1_2_lut_LC_4_32_3 .C_ON=1'b0;
    defparam \c0.tx2.i1_2_lut_LC_4_32_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i1_2_lut_LC_4_32_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.tx2.i1_2_lut_LC_4_32_3  (
            .in0(N__21468),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21324),
            .lcout(\c0.tx2.n23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i29_4_lut_LC_4_32_4 .C_ON=1'b0;
    defparam \c0.tx2.i29_4_lut_LC_4_32_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i29_4_lut_LC_4_32_4 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \c0.tx2.i29_4_lut_LC_4_32_4  (
            .in0(N__26131),
            .in1(N__21506),
            .in2(N__21296),
            .in3(N__21479),
            .lcout(),
            .ltout(\c0.tx2.n12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_i0_LC_4_32_5 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_i0_LC_4_32_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_SM_Main_i0_LC_4_32_5 .LUT_INIT=16'b0000000001110100;
    LogicCell40 \c0.tx2.r_SM_Main_i0_LC_4_32_5  (
            .in0(N__21469),
            .in1(N__21325),
            .in2(N__21437),
            .in3(N__21430),
            .lcout(\c0.tx2.r_SM_Main_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50374),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i4452_2_lut_LC_4_32_6 .C_ON=1'b0;
    defparam \c0.tx2.i4452_2_lut_LC_4_32_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i4452_2_lut_LC_4_32_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.tx2.i4452_2_lut_LC_4_32_6  (
            .in0(N__25888),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26185),
            .lcout(),
            .ltout(\c0.tx2.n6812_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i7506_4_lut_LC_4_32_7 .C_ON=1'b0;
    defparam \c0.tx2.i7506_4_lut_LC_4_32_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i7506_4_lut_LC_4_32_7 .LUT_INIT=16'b1101010100000000;
    LogicCell40 \c0.tx2.i7506_4_lut_LC_4_32_7  (
            .in0(N__21293),
            .in1(N__26130),
            .in2(N__21236),
            .in3(N__25926),
            .lcout(n9922),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i44_LC_5_16_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i44_LC_5_16_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i44_LC_5_16_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i44_LC_5_16_1  (
            .in0(N__45496),
            .in1(N__23678),
            .in2(_gnd_net_),
            .in3(N__22297),
            .lcout(data_in_5_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50270),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i52_LC_5_16_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i52_LC_5_16_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i52_LC_5_16_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i52_LC_5_16_7  (
            .in0(N__45497),
            .in1(N__25727),
            .in2(_gnd_net_),
            .in3(N__22296),
            .lcout(data_in_6_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50270),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i8_LC_5_17_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i8_LC_5_17_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i8_LC_5_17_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i8_LC_5_17_0  (
            .in0(N__21646),
            .in1(N__45488),
            .in2(_gnd_net_),
            .in3(N__27037),
            .lcout(data_in_0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50260),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15249_2_lut_LC_5_17_1 .C_ON=1'b0;
    defparam \c0.i15249_2_lut_LC_5_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.i15249_2_lut_LC_5_17_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i15249_2_lut_LC_5_17_1  (
            .in0(_gnd_net_),
            .in1(N__21645),
            .in2(_gnd_net_),
            .in3(N__27629),
            .lcout(),
            .ltout(\c0.n17697_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15315_4_lut_LC_5_17_2 .C_ON=1'b0;
    defparam \c0.i15315_4_lut_LC_5_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.i15315_4_lut_LC_5_17_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i15315_4_lut_LC_5_17_2  (
            .in0(N__24002),
            .in1(N__21624),
            .in2(N__21632),
            .in3(N__36242),
            .lcout(\c0.n17765 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i12_LC_5_17_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i12_LC_5_17_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i12_LC_5_17_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i12_LC_5_17_3  (
            .in0(N__45487),
            .in1(N__37566),
            .in2(_gnd_net_),
            .in3(N__27630),
            .lcout(\c0.data_in_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50260),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i5_LC_5_17_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i5_LC_5_17_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i5_LC_5_17_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_0___i5_LC_5_17_4  (
            .in0(N__21628),
            .in1(N__37660),
            .in2(_gnd_net_),
            .in3(N__45493),
            .lcout(data_in_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50260),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i14_LC_5_17_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i14_LC_5_17_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i14_LC_5_17_5 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \c0.data_in_0___i14_LC_5_17_5  (
            .in0(N__36243),
            .in1(_gnd_net_),
            .in2(N__45505),
            .in3(N__26989),
            .lcout(data_in_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50260),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i9_LC_5_17_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i9_LC_5_17_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i9_LC_5_17_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i9_LC_5_17_6  (
            .in0(N__24003),
            .in1(N__45489),
            .in2(_gnd_net_),
            .in3(N__27115),
            .lcout(\c0.data_in_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50260),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1057_LC_5_18_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1057_LC_5_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1057_LC_5_18_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1057_LC_5_18_0  (
            .in0(N__24970),
            .in1(N__21607),
            .in2(N__21554),
            .in3(N__22034),
            .lcout(n9054),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i11_LC_5_18_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i11_LC_5_18_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i11_LC_5_18_1 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \c0.data_in_0___i11_LC_5_18_1  (
            .in0(N__24378),
            .in1(N__28142),
            .in2(N__45503),
            .in3(_gnd_net_),
            .lcout(data_in_1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50271),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i3_LC_5_18_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i3_LC_5_18_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i3_LC_5_18_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i3_LC_5_18_2  (
            .in0(N__28143),
            .in1(N__45474),
            .in2(_gnd_net_),
            .in3(N__23737),
            .lcout(data_in_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50271),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i11_LC_5_18_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i11_LC_5_18_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i11_LC_5_18_3 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \c0.data_in_frame_0___i11_LC_5_18_3  (
            .in0(N__24125),
            .in1(N__28144),
            .in2(N__22042),
            .in3(N__31974),
            .lcout(\c0.data_in_frame_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50271),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_951_LC_5_18_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_951_LC_5_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_951_LC_5_18_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_951_LC_5_18_4  (
            .in0(N__22010),
            .in1(N__27509),
            .in2(_gnd_net_),
            .in3(N__28773),
            .lcout(\c0.n9208 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1113_LC_5_18_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1113_LC_5_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1113_LC_5_18_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1113_LC_5_18_5  (
            .in0(N__24759),
            .in1(N__21977),
            .in2(N__21953),
            .in3(N__22544),
            .lcout(n9100),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_969_LC_5_18_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_969_LC_5_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_969_LC_5_18_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_969_LC_5_18_6  (
            .in0(N__22451),
            .in1(N__21908),
            .in2(N__28979),
            .in3(N__21833),
            .lcout(n6_adj_2583),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i19_LC_5_18_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i19_LC_5_18_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i19_LC_5_18_7 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \c0.data_in_0___i19_LC_5_18_7  (
            .in0(N__37518),
            .in1(N__24377),
            .in2(N__45504),
            .in3(_gnd_net_),
            .lcout(data_in_2_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50271),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_861_LC_5_19_0 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_861_LC_5_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_861_LC_5_19_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_861_LC_5_19_0  (
            .in0(N__22155),
            .in1(N__21869),
            .in2(N__21838),
            .in3(N__21785),
            .lcout(),
            .ltout(\c0.n10_adj_2430_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_adj_959_LC_5_19_1 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_adj_959_LC_5_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_adj_959_LC_5_19_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_adj_959_LC_5_19_1  (
            .in0(N__21768),
            .in1(N__21727),
            .in2(N__21689),
            .in3(N__21686),
            .lcout(\c0.n8695 ),
            .ltout(\c0.n8695_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_886_LC_5_19_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_886_LC_5_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_886_LC_5_19_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_886_LC_5_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22193),
            .in3(N__28335),
            .lcout(\c0.n8064 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1049_LC_5_19_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1049_LC_5_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1049_LC_5_19_3 .LUT_INIT=16'b0110011000111100;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1049_LC_5_19_3  (
            .in0(N__25112),
            .in1(N__23065),
            .in2(N__36961),
            .in3(N__24069),
            .lcout(\c0.n8867 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i7_LC_5_19_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i7_LC_5_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i7_LC_5_19_4 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \c0.data_in_frame_0___i7_LC_5_19_4  (
            .in0(N__24071),
            .in1(N__22161),
            .in2(N__31996),
            .in3(N__27749),
            .lcout(\c0.data_in_frame_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50277),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i29_LC_5_19_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i29_LC_5_19_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i29_LC_5_19_5 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \c0.data_in_frame_0___i29_LC_5_19_5  (
            .in0(N__27908),
            .in1(N__24072),
            .in2(N__22133),
            .in3(N__31988),
            .lcout(\c0.data_in_frame_3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50277),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i3_LC_5_19_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i3_LC_5_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i3_LC_5_19_6 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \c0.data_in_frame_0___i3_LC_5_19_6  (
            .in0(N__24070),
            .in1(N__29001),
            .in2(N__31995),
            .in3(N__23741),
            .lcout(\c0.data_in_frame_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50277),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i41_LC_5_19_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i41_LC_5_19_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i41_LC_5_19_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i41_LC_5_19_7  (
            .in0(N__45460),
            .in1(N__22086),
            .in2(_gnd_net_),
            .in3(N__23830),
            .lcout(data_in_5_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50277),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3919_3_lut_4_lut_LC_5_20_0 .C_ON=1'b0;
    defparam \c0.i3919_3_lut_4_lut_LC_5_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3919_3_lut_4_lut_LC_5_20_0 .LUT_INIT=16'b1010101011100010;
    LogicCell40 \c0.i3919_3_lut_4_lut_LC_5_20_0  (
            .in0(N__22856),
            .in1(N__34553),
            .in2(N__22063),
            .in3(N__28008),
            .lcout(n2585),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i63_LC_5_20_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i63_LC_5_20_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i63_LC_5_20_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i63_LC_5_20_1  (
            .in0(N__45455),
            .in1(N__38761),
            .in2(_gnd_net_),
            .in3(N__22059),
            .lcout(data_in_7_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50283),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i55_LC_5_20_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i55_LC_5_20_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i55_LC_5_20_2 .LUT_INIT=16'b1110001011100010;
    LogicCell40 \c0.data_in_0___i55_LC_5_20_2  (
            .in0(N__31287),
            .in1(N__45456),
            .in2(N__22064),
            .in3(_gnd_net_),
            .lcout(data_in_6_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50283),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i57_LC_5_20_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i57_LC_5_20_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i57_LC_5_20_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i57_LC_5_20_3  (
            .in0(N__45454),
            .in1(N__23905),
            .in2(_gnd_net_),
            .in3(N__24598),
            .lcout(data_in_7_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50283),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3935_3_lut_4_lut_LC_5_20_4 .C_ON=1'b0;
    defparam \c0.i3935_3_lut_4_lut_LC_5_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3935_3_lut_4_lut_LC_5_20_4 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \c0.i3935_3_lut_4_lut_LC_5_20_4  (
            .in0(N__23043),
            .in1(N__34552),
            .in2(N__31291),
            .in3(N__28007),
            .lcout(n2593),
            .ltout(n2593_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_LC_5_20_5 .C_ON=1'b0;
    defparam \c0.i6_4_lut_LC_5_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_LC_5_20_5 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \c0.i6_4_lut_LC_5_20_5  (
            .in0(N__28920),
            .in1(N__22261),
            .in2(N__22361),
            .in3(N__24901),
            .lcout(\c0.n22_adj_2461 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3921_3_lut_4_lut_LC_5_20_6 .C_ON=1'b0;
    defparam \c0.i3921_3_lut_4_lut_LC_5_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3921_3_lut_4_lut_LC_5_20_6 .LUT_INIT=16'b1010101011100010;
    LogicCell40 \c0.i3921_3_lut_4_lut_LC_5_20_6  (
            .in0(N__28492),
            .in1(N__34554),
            .in2(N__36223),
            .in3(N__28009),
            .lcout(n2586),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1103_LC_5_20_7 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1103_LC_5_20_7 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1103_LC_5_20_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1103_LC_5_20_7  (
            .in0(N__27516),
            .in1(N__22334),
            .in2(N__22705),
            .in3(N__24781),
            .lcout(\c0.n17412 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3929_3_lut_4_lut_LC_5_21_1 .C_ON=1'b0;
    defparam \c0.i3929_3_lut_4_lut_LC_5_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3929_3_lut_4_lut_LC_5_21_1 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \c0.i3929_3_lut_4_lut_LC_5_21_1  (
            .in0(N__37016),
            .in1(N__34569),
            .in2(N__22695),
            .in3(N__28004),
            .lcout(n2590),
            .ltout(n2590_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_885_LC_5_21_2 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_885_LC_5_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_885_LC_5_21_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_885_LC_5_21_2  (
            .in0(N__22768),
            .in1(N__22496),
            .in2(N__22313),
            .in3(N__24758),
            .lcout(\c0.n10_adj_2450 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3941_3_lut_4_lut_LC_5_21_3 .C_ON=1'b0;
    defparam \c0.i3941_3_lut_4_lut_LC_5_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3941_3_lut_4_lut_LC_5_21_3 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \c0.i3941_3_lut_4_lut_LC_5_21_3  (
            .in0(N__22902),
            .in1(N__34570),
            .in2(N__22304),
            .in3(N__28005),
            .lcout(n2596),
            .ltout(n2596_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_971_LC_5_21_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_971_LC_5_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_971_LC_5_21_4 .LUT_INIT=16'b1011111001111101;
    LogicCell40 \c0.i3_4_lut_adj_971_LC_5_21_4  (
            .in0(N__22262),
            .in1(N__25346),
            .in2(N__22244),
            .in3(N__24476),
            .lcout(\c0.n10_adj_2498 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3925_3_lut_4_lut_LC_5_21_5 .C_ON=1'b0;
    defparam \c0.i3925_3_lut_4_lut_LC_5_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3925_3_lut_4_lut_LC_5_21_5 .LUT_INIT=16'b1010101011100010;
    LogicCell40 \c0.i3925_3_lut_4_lut_LC_5_21_5  (
            .in0(N__22224),
            .in1(N__34571),
            .in2(N__25723),
            .in3(N__28006),
            .lcout(n2588),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_adj_1053_LC_5_21_6 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_adj_1053_LC_5_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_adj_1053_LC_5_21_6 .LUT_INIT=16'b1111111101101001;
    LogicCell40 \c0.i1_3_lut_4_lut_adj_1053_LC_5_21_6  (
            .in0(N__22769),
            .in1(N__22729),
            .in2(N__24698),
            .in3(N__24482),
            .lcout(\c0.n17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i58_LC_5_21_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i58_LC_5_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i58_LC_5_21_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.data_in_frame_0___i58_LC_5_21_7  (
            .in0(_gnd_net_),
            .in1(N__22712),
            .in2(_gnd_net_),
            .in3(N__31906),
            .lcout(\c0.data_in_frame_7_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50288),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1106_LC_5_22_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1106_LC_5_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1106_LC_5_22_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1106_LC_5_22_0  (
            .in0(N__22653),
            .in1(N__22636),
            .in2(N__22590),
            .in3(N__22552),
            .lcout(\c0.n17403 ),
            .ltout(\c0.n17403_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_985_LC_5_22_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_985_LC_5_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_985_LC_5_22_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_985_LC_5_22_1  (
            .in0(N__24438),
            .in1(N__22926),
            .in2(N__22499),
            .in3(N__22492),
            .lcout(n9283),
            .ltout(n9283_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_2_lut_3_lut_4_lut_LC_5_22_2.C_ON=1'b0;
    defparam i3_2_lut_3_lut_4_lut_LC_5_22_2.SEQ_MODE=4'b0000;
    defparam i3_2_lut_3_lut_4_lut_LC_5_22_2.LUT_INIT=16'b0110100110010110;
    LogicCell40 i3_2_lut_3_lut_4_lut_LC_5_22_2 (
            .in0(N__25587),
            .in1(N__25064),
            .in2(N__22430),
            .in3(N__28094),
            .lcout(n16_adj_2656),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i136_LC_5_22_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i136_LC_5_22_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i136_LC_5_22_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i136_LC_5_22_3  (
            .in0(N__34964),
            .in1(N__22420),
            .in2(_gnd_net_),
            .in3(N__32833),
            .lcout(data_out_frame2_16_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50294),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13614_3_lut_4_lut_LC_5_22_4 .C_ON=1'b0;
    defparam \c0.i13614_3_lut_4_lut_LC_5_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i13614_3_lut_4_lut_LC_5_22_4 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \c0.i13614_3_lut_4_lut_LC_5_22_4  (
            .in0(N__38801),
            .in1(N__34605),
            .in2(N__29245),
            .in3(N__34446),
            .lcout(\c0.n15927 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_974_LC_5_22_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_974_LC_5_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_974_LC_5_22_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_974_LC_5_22_6  (
            .in0(N__22927),
            .in1(N__24439),
            .in2(_gnd_net_),
            .in3(N__28481),
            .lcout(\c0.n9219 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_829_LC_5_23_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_829_LC_5_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_829_LC_5_23_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_829_LC_5_23_0  (
            .in0(_gnd_net_),
            .in1(N__28339),
            .in2(_gnd_net_),
            .in3(N__25331),
            .lcout(\c0.n17519 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_LC_5_23_1 .C_ON=1'b0;
    defparam \c0.i9_4_lut_LC_5_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_LC_5_23_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_LC_5_23_1  (
            .in0(N__28254),
            .in1(N__28563),
            .in2(N__24614),
            .in3(N__23066),
            .lcout(),
            .ltout(\c0.n22_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_LC_5_23_2 .C_ON=1'b0;
    defparam \c0.i11_4_lut_LC_5_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_LC_5_23_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_LC_5_23_2  (
            .in0(N__23051),
            .in1(N__23023),
            .in2(N__22991),
            .in3(N__22988),
            .lcout(),
            .ltout(\c0.n24_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_LC_5_23_3 .C_ON=1'b0;
    defparam \c0.i12_4_lut_LC_5_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_LC_5_23_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_4_lut_LC_5_23_3  (
            .in0(N__28397),
            .in1(N__22982),
            .in2(N__22976),
            .in3(N__22862),
            .lcout(\c0.n9355 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i86_LC_5_23_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i86_LC_5_23_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i86_LC_5_23_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.data_in_frame_0___i86_LC_5_23_4  (
            .in0(_gnd_net_),
            .in1(N__32936),
            .in2(_gnd_net_),
            .in3(N__31973),
            .lcout(\c0.data_in_frame_10_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50302),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_3_lut_4_lut_adj_907_LC_5_23_5 .C_ON=1'b0;
    defparam \c0.i4_3_lut_4_lut_adj_907_LC_5_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_3_lut_4_lut_adj_907_LC_5_23_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_3_lut_4_lut_adj_907_LC_5_23_5  (
            .in0(N__25332),
            .in1(N__28341),
            .in2(N__24691),
            .in3(N__22871),
            .lcout(\c0.n11_adj_2453 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_LC_5_23_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_LC_5_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_LC_5_23_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_LC_5_23_6  (
            .in0(N__22961),
            .in1(N__22903),
            .in2(_gnd_net_),
            .in3(N__22928),
            .lcout(\c0.n9144 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_3_lut_LC_5_23_7 .C_ON=1'b0;
    defparam \c0.i7_3_lut_LC_5_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.i7_3_lut_LC_5_23_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i7_3_lut_LC_5_23_7  (
            .in0(N__22904),
            .in1(N__25525),
            .in2(_gnd_net_),
            .in3(N__22870),
            .lcout(\c0.n20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_980_LC_5_24_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_980_LC_5_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_980_LC_5_24_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_980_LC_5_24_0  (
            .in0(N__22846),
            .in1(N__28491),
            .in2(N__22801),
            .in3(N__22784),
            .lcout(\c0.n17582 ),
            .ltout(\c0.n17582_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i168_LC_5_24_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i168_LC_5_24_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i168_LC_5_24_1 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.data_out_frame2_0___i168_LC_5_24_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23174),
            .in3(N__23098),
            .lcout(\c0.data_out_frame2_20_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50310),
            .ce(N__32814),
            .sr(_gnd_net_));
    defparam \c0.i3869_3_lut_4_lut_LC_5_24_2 .C_ON=1'b0;
    defparam \c0.i3869_3_lut_4_lut_LC_5_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3869_3_lut_4_lut_LC_5_24_2 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \c0.i3869_3_lut_4_lut_LC_5_24_2  (
            .in0(N__34628),
            .in1(N__30473),
            .in2(N__36685),
            .in3(N__34445),
            .lcout(n2560),
            .ltout(n2560_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_860_LC_5_24_3 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_860_LC_5_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_860_LC_5_24_3 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \c0.i2_4_lut_adj_860_LC_5_24_3  (
            .in0(N__23144),
            .in1(N__23135),
            .in2(N__23129),
            .in3(N__23083),
            .lcout(),
            .ltout(\c0.n18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_867_LC_5_24_4 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_867_LC_5_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_867_LC_5_24_4 .LUT_INIT=16'b1111011111111011;
    LogicCell40 \c0.i9_4_lut_adj_867_LC_5_24_4  (
            .in0(N__23125),
            .in1(N__23108),
            .in2(N__23102),
            .in3(N__24470),
            .lcout(\c0.n25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_928_LC_5_24_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_928_LC_5_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_928_LC_5_24_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_928_LC_5_24_5  (
            .in0(N__36872),
            .in1(N__32264),
            .in2(N__36625),
            .in3(N__36579),
            .lcout(\c0.n17418 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3893_3_lut_4_lut_LC_5_24_6 .C_ON=1'b0;
    defparam \c0.i3893_3_lut_4_lut_LC_5_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3893_3_lut_4_lut_LC_5_24_6 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \c0.i3893_3_lut_4_lut_LC_5_24_6  (
            .in0(N__34627),
            .in1(N__29681),
            .in2(N__36581),
            .in3(N__34444),
            .lcout(n2572),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_2_lut_LC_5_25_0 .C_ON=1'b1;
    defparam \c0.tx.add_59_2_lut_LC_5_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_2_lut_LC_5_25_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx.add_59_2_lut_LC_5_25_0  (
            .in0(N__29700),
            .in1(N__29659),
            .in2(_gnd_net_),
            .in3(N__23072),
            .lcout(n18104),
            .ltout(),
            .carryin(bfn_5_25_0_),
            .carryout(\c0.tx.n16357 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_3_lut_LC_5_25_1 .C_ON=1'b1;
    defparam \c0.tx.add_59_3_lut_LC_5_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_3_lut_LC_5_25_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx.add_59_3_lut_LC_5_25_1  (
            .in0(N__29712),
            .in1(N__29582),
            .in2(_gnd_net_),
            .in3(N__23069),
            .lcout(n18101),
            .ltout(),
            .carryin(\c0.tx.n16357 ),
            .carryout(\c0.tx.n16358 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_4_lut_LC_5_25_2 .C_ON=1'b1;
    defparam \c0.tx.add_59_4_lut_LC_5_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_4_lut_LC_5_25_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx.add_59_4_lut_LC_5_25_2  (
            .in0(N__29699),
            .in1(N__33794),
            .in2(_gnd_net_),
            .in3(N__23228),
            .lcout(n18102),
            .ltout(),
            .carryin(\c0.tx.n16358 ),
            .carryout(\c0.tx.n16359 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_5_lut_LC_5_25_3 .C_ON=1'b1;
    defparam \c0.tx.add_59_5_lut_LC_5_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_5_lut_LC_5_25_3 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx.add_59_5_lut_LC_5_25_3  (
            .in0(N__29713),
            .in1(N__29620),
            .in2(_gnd_net_),
            .in3(N__23225),
            .lcout(n18103),
            .ltout(),
            .carryin(\c0.tx.n16359 ),
            .carryout(\c0.tx.n16360 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_6_lut_LC_5_25_4 .C_ON=1'b1;
    defparam \c0.tx.add_59_6_lut_LC_5_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_6_lut_LC_5_25_4 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx.add_59_6_lut_LC_5_25_4  (
            .in0(N__29701),
            .in1(N__29602),
            .in2(_gnd_net_),
            .in3(N__23222),
            .lcout(n18097),
            .ltout(),
            .carryin(\c0.tx.n16360 ),
            .carryout(\c0.tx.n16361 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_7_lut_LC_5_25_5 .C_ON=1'b1;
    defparam \c0.tx.add_59_7_lut_LC_5_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_7_lut_LC_5_25_5 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx.add_59_7_lut_LC_5_25_5  (
            .in0(N__29714),
            .in1(N__29640),
            .in2(_gnd_net_),
            .in3(N__23219),
            .lcout(n18054),
            .ltout(),
            .carryin(\c0.tx.n16361 ),
            .carryout(\c0.tx.n16362 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_8_lut_LC_5_25_6 .C_ON=1'b1;
    defparam \c0.tx.add_59_8_lut_LC_5_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_8_lut_LC_5_25_6 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx.add_59_8_lut_LC_5_25_6  (
            .in0(N__33832),
            .in1(N__37265),
            .in2(_gnd_net_),
            .in3(N__23216),
            .lcout(n18010),
            .ltout(),
            .carryin(\c0.tx.n16362 ),
            .carryout(\c0.tx.n16363 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_9_lut_LC_5_25_7 .C_ON=1'b1;
    defparam \c0.tx.add_59_9_lut_LC_5_25_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_9_lut_LC_5_25_7 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.tx.add_59_9_lut_LC_5_25_7  (
            .in0(N__33831),
            .in1(N__37229),
            .in2(_gnd_net_),
            .in3(N__23213),
            .lcout(n17952),
            .ltout(),
            .carryin(\c0.tx.n16363 ),
            .carryout(\c0.tx.n16364 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_10_lut_LC_5_26_0 .C_ON=1'b0;
    defparam \c0.tx.add_59_10_lut_LC_5_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_10_lut_LC_5_26_0 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \c0.tx.add_59_10_lut_LC_5_26_0  (
            .in0(N__37325),
            .in1(N__33833),
            .in2(_gnd_net_),
            .in3(N__23210),
            .lcout(n17950),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i133_LC_5_26_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i133_LC_5_26_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i133_LC_5_26_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \c0.data_out_frame2_0___i133_LC_5_26_2  (
            .in0(N__32743),
            .in1(_gnd_net_),
            .in2(N__35149),
            .in3(N__26221),
            .lcout(data_out_frame2_16_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50327),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1081_LC_5_26_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1081_LC_5_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1081_LC_5_26_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1081_LC_5_26_3  (
            .in0(N__25636),
            .in1(N__28692),
            .in2(_gnd_net_),
            .in3(N__32045),
            .lcout(n9051),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_870_LC_5_26_5 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_870_LC_5_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_870_LC_5_26_5 .LUT_INIT=16'b1111110111111000;
    LogicCell40 \c0.i1_4_lut_adj_870_LC_5_26_5  (
            .in0(N__33272),
            .in1(N__25132),
            .in2(N__33367),
            .in3(N__23207),
            .lcout(\c0.n136 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i79_LC_5_26_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i79_LC_5_26_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i79_LC_5_26_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i79_LC_5_26_6  (
            .in0(N__32744),
            .in1(N__36354),
            .in2(_gnd_net_),
            .in3(N__23377),
            .lcout(data_out_frame2_9_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50327),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i116_LC_5_26_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i116_LC_5_26_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i116_LC_5_26_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i116_LC_5_26_7  (
            .in0(N__35250),
            .in1(N__23350),
            .in2(_gnd_net_),
            .in3(N__32745),
            .lcout(data_out_frame2_14_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50327),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16041_LC_5_27_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16041_LC_5_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16041_LC_5_27_0 .LUT_INIT=16'b1101100010101010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_16041_LC_5_27_0  (
            .in0(N__30695),
            .in1(N__23362),
            .in2(N__23351),
            .in3(N__31052),
            .lcout(),
            .ltout(\c0.n18516_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18516_bdd_4_lut_LC_5_27_1 .C_ON=1'b0;
    defparam \c0.n18516_bdd_4_lut_LC_5_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.n18516_bdd_4_lut_LC_5_27_1 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n18516_bdd_4_lut_LC_5_27_1  (
            .in0(N__31053),
            .in1(N__25777),
            .in2(N__23336),
            .in3(N__23333),
            .lcout(\c0.n17818 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16011_LC_5_27_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16011_LC_5_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16011_LC_5_27_3 .LUT_INIT=16'b1010111111000000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_16011_LC_5_27_3  (
            .in0(N__23311),
            .in1(N__23299),
            .in2(N__31096),
            .in3(N__30694),
            .lcout(\c0.n18480 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12304_4_lut_LC_5_27_4 .C_ON=1'b0;
    defparam \c0.i12304_4_lut_LC_5_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.i12304_4_lut_LC_5_27_4 .LUT_INIT=16'b0010001001110010;
    LogicCell40 \c0.i12304_4_lut_LC_5_27_4  (
            .in0(N__33514),
            .in1(N__23276),
            .in2(N__33148),
            .in3(N__23270),
            .lcout(\c0.n14631 ),
            .ltout(\c0.n14631_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i5_LC_5_27_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i5_LC_5_27_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i5_LC_5_27_5 .LUT_INIT=16'b1111010111110000;
    LogicCell40 \c0.data_out_frame2_0___i5_LC_5_27_5  (
            .in0(N__33666),
            .in1(_gnd_net_),
            .in2(N__23252),
            .in3(N__26710),
            .lcout(\c0.data_out_frame2_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50336),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i3_LC_5_27_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i3_LC_5_27_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i3_LC_5_27_6 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \c0.data_out_frame2_0___i3_LC_5_27_6  (
            .in0(N__23242),
            .in1(N__33667),
            .in2(_gnd_net_),
            .in3(N__25789),
            .lcout(\c0.data_out_frame2_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50336),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i45_LC_5_28_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i45_LC_5_28_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i45_LC_5_28_0 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \c0.data_out_frame2_0___i45_LC_5_28_0  (
            .in0(N__36459),
            .in1(N__26863),
            .in2(N__32842),
            .in3(_gnd_net_),
            .lcout(data_out_frame2_5_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50346),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i68_LC_5_28_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i68_LC_5_28_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i68_LC_5_28_1 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \c0.data_out_frame2_0___i68_LC_5_28_1  (
            .in0(_gnd_net_),
            .in1(N__32834),
            .in2(N__23492),
            .in3(N__35194),
            .lcout(data_out_frame2_8_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50346),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_843_LC_5_28_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_843_LC_5_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_843_LC_5_28_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_843_LC_5_28_2  (
            .in0(_gnd_net_),
            .in1(N__32987),
            .in2(_gnd_net_),
            .in3(N__36686),
            .lcout(\c0.n17482 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18522_bdd_4_lut_LC_5_28_3 .C_ON=1'b0;
    defparam \c0.n18522_bdd_4_lut_LC_5_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.n18522_bdd_4_lut_LC_5_28_3 .LUT_INIT=16'b1110111001010000;
    LogicCell40 \c0.n18522_bdd_4_lut_LC_5_28_3  (
            .in0(N__31075),
            .in1(N__23509),
            .in2(N__23491),
            .in3(N__23477),
            .lcout(\c0.n17815 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15819_3_lut_LC_5_28_4 .C_ON=1'b0;
    defparam \c0.i15819_3_lut_LC_5_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.i15819_3_lut_LC_5_28_4 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \c0.i15819_3_lut_LC_5_28_4  (
            .in0(N__30722),
            .in1(N__23468),
            .in2(_gnd_net_),
            .in3(N__31074),
            .lcout(\c0.n18076 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18588_bdd_4_lut_LC_5_28_7 .C_ON=1'b0;
    defparam \c0.n18588_bdd_4_lut_LC_5_28_7 .SEQ_MODE=4'b0000;
    defparam \c0.n18588_bdd_4_lut_LC_5_28_7 .LUT_INIT=16'b1110111001010000;
    LogicCell40 \c0.n18588_bdd_4_lut_LC_5_28_7  (
            .in0(N__31073),
            .in1(N__23431),
            .in2(N__23420),
            .in3(N__23405),
            .lcout(\c0.n17785 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2269__i0_LC_5_29_0.C_ON=1'b1;
    defparam rand_data_2269__i0_LC_5_29_0.SEQ_MODE=4'b1000;
    defparam rand_data_2269__i0_LC_5_29_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2269__i0_LC_5_29_0 (
            .in0(_gnd_net_),
            .in1(N__34201),
            .in2(_gnd_net_),
            .in3(N__23387),
            .lcout(rand_data_0),
            .ltout(),
            .carryin(bfn_5_29_0_),
            .carryout(n16319),
            .clk(N__50356),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2269__i1_LC_5_29_1.C_ON=1'b1;
    defparam rand_data_2269__i1_LC_5_29_1.SEQ_MODE=4'b1000;
    defparam rand_data_2269__i1_LC_5_29_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2269__i1_LC_5_29_1 (
            .in0(_gnd_net_),
            .in1(N__34139),
            .in2(_gnd_net_),
            .in3(N__23384),
            .lcout(rand_data_1),
            .ltout(),
            .carryin(n16319),
            .carryout(n16320),
            .clk(N__50356),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2269__i2_LC_5_29_2.C_ON=1'b1;
    defparam rand_data_2269__i2_LC_5_29_2.SEQ_MODE=4'b1000;
    defparam rand_data_2269__i2_LC_5_29_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2269__i2_LC_5_29_2 (
            .in0(_gnd_net_),
            .in1(N__34078),
            .in2(_gnd_net_),
            .in3(N__23381),
            .lcout(rand_data_2),
            .ltout(),
            .carryin(n16320),
            .carryout(n16321),
            .clk(N__50356),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2269__i3_LC_5_29_3.C_ON=1'b1;
    defparam rand_data_2269__i3_LC_5_29_3.SEQ_MODE=4'b1000;
    defparam rand_data_2269__i3_LC_5_29_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2269__i3_LC_5_29_3 (
            .in0(_gnd_net_),
            .in1(N__35190),
            .in2(_gnd_net_),
            .in3(N__23555),
            .lcout(rand_data_3),
            .ltout(),
            .carryin(n16321),
            .carryout(n16322),
            .clk(N__50356),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2269__i4_LC_5_29_4.C_ON=1'b1;
    defparam rand_data_2269__i4_LC_5_29_4.SEQ_MODE=4'b1000;
    defparam rand_data_2269__i4_LC_5_29_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2269__i4_LC_5_29_4 (
            .in0(_gnd_net_),
            .in1(N__35133),
            .in2(_gnd_net_),
            .in3(N__23552),
            .lcout(rand_data_4),
            .ltout(),
            .carryin(n16322),
            .carryout(n16323),
            .clk(N__50356),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2269__i5_LC_5_29_5.C_ON=1'b1;
    defparam rand_data_2269__i5_LC_5_29_5.SEQ_MODE=4'b1000;
    defparam rand_data_2269__i5_LC_5_29_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2269__i5_LC_5_29_5 (
            .in0(_gnd_net_),
            .in1(N__35071),
            .in2(_gnd_net_),
            .in3(N__23549),
            .lcout(rand_data_5),
            .ltout(),
            .carryin(n16323),
            .carryout(n16324),
            .clk(N__50356),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2269__i6_LC_5_29_6.C_ON=1'b1;
    defparam rand_data_2269__i6_LC_5_29_6.SEQ_MODE=4'b1000;
    defparam rand_data_2269__i6_LC_5_29_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2269__i6_LC_5_29_6 (
            .in0(_gnd_net_),
            .in1(N__35013),
            .in2(_gnd_net_),
            .in3(N__23546),
            .lcout(rand_data_6),
            .ltout(),
            .carryin(n16324),
            .carryout(n16325),
            .clk(N__50356),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2269__i7_LC_5_29_7.C_ON=1'b1;
    defparam rand_data_2269__i7_LC_5_29_7.SEQ_MODE=4'b1000;
    defparam rand_data_2269__i7_LC_5_29_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2269__i7_LC_5_29_7 (
            .in0(_gnd_net_),
            .in1(N__34938),
            .in2(_gnd_net_),
            .in3(N__23543),
            .lcout(rand_data_7),
            .ltout(),
            .carryin(n16325),
            .carryout(n16326),
            .clk(N__50356),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2269__i8_LC_5_30_0.C_ON=1'b1;
    defparam rand_data_2269__i8_LC_5_30_0.SEQ_MODE=4'b1000;
    defparam rand_data_2269__i8_LC_5_30_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2269__i8_LC_5_30_0 (
            .in0(_gnd_net_),
            .in1(N__34856),
            .in2(_gnd_net_),
            .in3(N__23540),
            .lcout(rand_data_8),
            .ltout(),
            .carryin(bfn_5_30_0_),
            .carryout(n16327),
            .clk(N__50367),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2269__i9_LC_5_30_1.C_ON=1'b1;
    defparam rand_data_2269__i9_LC_5_30_1.SEQ_MODE=4'b1000;
    defparam rand_data_2269__i9_LC_5_30_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2269__i9_LC_5_30_1 (
            .in0(_gnd_net_),
            .in1(N__34801),
            .in2(_gnd_net_),
            .in3(N__23537),
            .lcout(rand_data_9),
            .ltout(),
            .carryin(n16327),
            .carryout(n16328),
            .clk(N__50367),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2269__i10_LC_5_30_2.C_ON=1'b1;
    defparam rand_data_2269__i10_LC_5_30_2.SEQ_MODE=4'b1000;
    defparam rand_data_2269__i10_LC_5_30_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2269__i10_LC_5_30_2 (
            .in0(_gnd_net_),
            .in1(N__34736),
            .in2(_gnd_net_),
            .in3(N__23534),
            .lcout(rand_data_10),
            .ltout(),
            .carryin(n16328),
            .carryout(n16329),
            .clk(N__50367),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2269__i11_LC_5_30_3.C_ON=1'b1;
    defparam rand_data_2269__i11_LC_5_30_3.SEQ_MODE=4'b1000;
    defparam rand_data_2269__i11_LC_5_30_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2269__i11_LC_5_30_3 (
            .in0(_gnd_net_),
            .in1(N__35685),
            .in2(_gnd_net_),
            .in3(N__23531),
            .lcout(rand_data_11),
            .ltout(),
            .carryin(n16329),
            .carryout(n16330),
            .clk(N__50367),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2269__i12_LC_5_30_4.C_ON=1'b1;
    defparam rand_data_2269__i12_LC_5_30_4.SEQ_MODE=4'b1000;
    defparam rand_data_2269__i12_LC_5_30_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2269__i12_LC_5_30_4 (
            .in0(_gnd_net_),
            .in1(N__35632),
            .in2(_gnd_net_),
            .in3(N__23585),
            .lcout(rand_data_12),
            .ltout(),
            .carryin(n16330),
            .carryout(n16331),
            .clk(N__50367),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2269__i13_LC_5_30_5.C_ON=1'b1;
    defparam rand_data_2269__i13_LC_5_30_5.SEQ_MODE=4'b1000;
    defparam rand_data_2269__i13_LC_5_30_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2269__i13_LC_5_30_5 (
            .in0(_gnd_net_),
            .in1(N__35563),
            .in2(_gnd_net_),
            .in3(N__23582),
            .lcout(rand_data_13),
            .ltout(),
            .carryin(n16331),
            .carryout(n16332),
            .clk(N__50367),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2269__i14_LC_5_30_6.C_ON=1'b1;
    defparam rand_data_2269__i14_LC_5_30_6.SEQ_MODE=4'b1000;
    defparam rand_data_2269__i14_LC_5_30_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2269__i14_LC_5_30_6 (
            .in0(_gnd_net_),
            .in1(N__35503),
            .in2(_gnd_net_),
            .in3(N__23579),
            .lcout(rand_data_14),
            .ltout(),
            .carryin(n16332),
            .carryout(n16333),
            .clk(N__50367),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2269__i15_LC_5_30_7.C_ON=1'b1;
    defparam rand_data_2269__i15_LC_5_30_7.SEQ_MODE=4'b1000;
    defparam rand_data_2269__i15_LC_5_30_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2269__i15_LC_5_30_7 (
            .in0(_gnd_net_),
            .in1(N__35437),
            .in2(_gnd_net_),
            .in3(N__23576),
            .lcout(rand_data_15),
            .ltout(),
            .carryin(n16333),
            .carryout(n16334),
            .clk(N__50367),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2269__i16_LC_5_31_0.C_ON=1'b1;
    defparam rand_data_2269__i16_LC_5_31_0.SEQ_MODE=4'b1000;
    defparam rand_data_2269__i16_LC_5_31_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2269__i16_LC_5_31_0 (
            .in0(_gnd_net_),
            .in1(N__35386),
            .in2(_gnd_net_),
            .in3(N__23573),
            .lcout(rand_data_16),
            .ltout(),
            .carryin(bfn_5_31_0_),
            .carryout(n16335),
            .clk(N__50375),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2269__i17_LC_5_31_1.C_ON=1'b1;
    defparam rand_data_2269__i17_LC_5_31_1.SEQ_MODE=4'b1000;
    defparam rand_data_2269__i17_LC_5_31_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2269__i17_LC_5_31_1 (
            .in0(_gnd_net_),
            .in1(N__35335),
            .in2(_gnd_net_),
            .in3(N__23570),
            .lcout(rand_data_17),
            .ltout(),
            .carryin(n16335),
            .carryout(n16336),
            .clk(N__50375),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2269__i18_LC_5_31_2.C_ON=1'b1;
    defparam rand_data_2269__i18_LC_5_31_2.SEQ_MODE=4'b1000;
    defparam rand_data_2269__i18_LC_5_31_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2269__i18_LC_5_31_2 (
            .in0(_gnd_net_),
            .in1(N__35283),
            .in2(_gnd_net_),
            .in3(N__23567),
            .lcout(rand_data_18),
            .ltout(),
            .carryin(n16336),
            .carryout(n16337),
            .clk(N__50375),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2269__i19_LC_5_31_3.C_ON=1'b1;
    defparam rand_data_2269__i19_LC_5_31_3.SEQ_MODE=4'b1000;
    defparam rand_data_2269__i19_LC_5_31_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2269__i19_LC_5_31_3 (
            .in0(_gnd_net_),
            .in1(N__35239),
            .in2(_gnd_net_),
            .in3(N__23564),
            .lcout(rand_data_19),
            .ltout(),
            .carryin(n16337),
            .carryout(n16338),
            .clk(N__50375),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2269__i20_LC_5_31_4.C_ON=1'b1;
    defparam rand_data_2269__i20_LC_5_31_4.SEQ_MODE=4'b1000;
    defparam rand_data_2269__i20_LC_5_31_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2269__i20_LC_5_31_4 (
            .in0(_gnd_net_),
            .in1(N__36131),
            .in2(_gnd_net_),
            .in3(N__23561),
            .lcout(rand_data_20),
            .ltout(),
            .carryin(n16338),
            .carryout(n16339),
            .clk(N__50375),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2269__i21_LC_5_31_5.C_ON=1'b1;
    defparam rand_data_2269__i21_LC_5_31_5.SEQ_MODE=4'b1000;
    defparam rand_data_2269__i21_LC_5_31_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2269__i21_LC_5_31_5 (
            .in0(_gnd_net_),
            .in1(N__36076),
            .in2(_gnd_net_),
            .in3(N__23558),
            .lcout(rand_data_21),
            .ltout(),
            .carryin(n16339),
            .carryout(n16340),
            .clk(N__50375),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2269__i22_LC_5_31_6.C_ON=1'b1;
    defparam rand_data_2269__i22_LC_5_31_6.SEQ_MODE=4'b1000;
    defparam rand_data_2269__i22_LC_5_31_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2269__i22_LC_5_31_6 (
            .in0(_gnd_net_),
            .in1(N__36027),
            .in2(_gnd_net_),
            .in3(N__23612),
            .lcout(rand_data_22),
            .ltout(),
            .carryin(n16340),
            .carryout(n16341),
            .clk(N__50375),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2269__i23_LC_5_31_7.C_ON=1'b1;
    defparam rand_data_2269__i23_LC_5_31_7.SEQ_MODE=4'b1000;
    defparam rand_data_2269__i23_LC_5_31_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2269__i23_LC_5_31_7 (
            .in0(_gnd_net_),
            .in1(N__35978),
            .in2(_gnd_net_),
            .in3(N__23609),
            .lcout(rand_data_23),
            .ltout(),
            .carryin(n16341),
            .carryout(n16342),
            .clk(N__50375),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2269__i24_LC_5_32_0.C_ON=1'b1;
    defparam rand_data_2269__i24_LC_5_32_0.SEQ_MODE=4'b1000;
    defparam rand_data_2269__i24_LC_5_32_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2269__i24_LC_5_32_0 (
            .in0(_gnd_net_),
            .in1(N__35920),
            .in2(_gnd_net_),
            .in3(N__23606),
            .lcout(rand_data_24),
            .ltout(),
            .carryin(bfn_5_32_0_),
            .carryout(n16343),
            .clk(N__50383),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2269__i25_LC_5_32_1.C_ON=1'b1;
    defparam rand_data_2269__i25_LC_5_32_1.SEQ_MODE=4'b1000;
    defparam rand_data_2269__i25_LC_5_32_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2269__i25_LC_5_32_1 (
            .in0(_gnd_net_),
            .in1(N__35860),
            .in2(_gnd_net_),
            .in3(N__23603),
            .lcout(rand_data_25),
            .ltout(),
            .carryin(n16343),
            .carryout(n16344),
            .clk(N__50383),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2269__i26_LC_5_32_2.C_ON=1'b1;
    defparam rand_data_2269__i26_LC_5_32_2.SEQ_MODE=4'b1000;
    defparam rand_data_2269__i26_LC_5_32_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2269__i26_LC_5_32_2 (
            .in0(_gnd_net_),
            .in1(N__35796),
            .in2(_gnd_net_),
            .in3(N__23600),
            .lcout(rand_data_26),
            .ltout(),
            .carryin(n16344),
            .carryout(n16345),
            .clk(N__50383),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2269__i27_LC_5_32_3.C_ON=1'b1;
    defparam rand_data_2269__i27_LC_5_32_3.SEQ_MODE=4'b1000;
    defparam rand_data_2269__i27_LC_5_32_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2269__i27_LC_5_32_3 (
            .in0(_gnd_net_),
            .in1(N__35749),
            .in2(_gnd_net_),
            .in3(N__23597),
            .lcout(rand_data_27),
            .ltout(),
            .carryin(n16345),
            .carryout(n16346),
            .clk(N__50383),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2269__i28_LC_5_32_4.C_ON=1'b1;
    defparam rand_data_2269__i28_LC_5_32_4.SEQ_MODE=4'b1000;
    defparam rand_data_2269__i28_LC_5_32_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2269__i28_LC_5_32_4 (
            .in0(_gnd_net_),
            .in1(N__36437),
            .in2(_gnd_net_),
            .in3(N__23594),
            .lcout(rand_data_28),
            .ltout(),
            .carryin(n16346),
            .carryout(n16347),
            .clk(N__50383),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2269__i29_LC_5_32_5.C_ON=1'b1;
    defparam rand_data_2269__i29_LC_5_32_5.SEQ_MODE=4'b1000;
    defparam rand_data_2269__i29_LC_5_32_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2269__i29_LC_5_32_5 (
            .in0(_gnd_net_),
            .in1(N__36383),
            .in2(_gnd_net_),
            .in3(N__23591),
            .lcout(rand_data_29),
            .ltout(),
            .carryin(n16347),
            .carryout(n16348),
            .clk(N__50383),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2269__i30_LC_5_32_6.C_ON=1'b1;
    defparam rand_data_2269__i30_LC_5_32_6.SEQ_MODE=4'b1000;
    defparam rand_data_2269__i30_LC_5_32_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2269__i30_LC_5_32_6 (
            .in0(_gnd_net_),
            .in1(N__36335),
            .in2(_gnd_net_),
            .in3(N__23588),
            .lcout(rand_data_30),
            .ltout(),
            .carryin(n16348),
            .carryout(n16349),
            .clk(N__50383),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2269__i31_LC_5_32_7.C_ON=1'b0;
    defparam rand_data_2269__i31_LC_5_32_7.SEQ_MODE=4'b1000;
    defparam rand_data_2269__i31_LC_5_32_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2269__i31_LC_5_32_7 (
            .in0(_gnd_net_),
            .in1(N__36287),
            .in2(_gnd_net_),
            .in3(N__23705),
            .lcout(rand_data_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50383),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i24_LC_6_16_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i24_LC_6_16_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i24_LC_6_16_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i24_LC_6_16_1  (
            .in0(N__45501),
            .in1(N__27275),
            .in2(_gnd_net_),
            .in3(N__23947),
            .lcout(data_in_2_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50278),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i36_LC_6_16_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i36_LC_6_16_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i36_LC_6_16_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i36_LC_6_16_7  (
            .in0(N__45502),
            .in1(N__27564),
            .in2(_gnd_net_),
            .in3(N__23679),
            .lcout(data_in_4_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50278),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15296_4_lut_LC_6_17_0 .C_ON=1'b0;
    defparam \c0.i15296_4_lut_LC_6_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.i15296_4_lut_LC_6_17_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i15296_4_lut_LC_6_17_0  (
            .in0(N__23945),
            .in1(N__27173),
            .in2(N__23977),
            .in3(N__27782),
            .lcout(\c0.n17745 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i30_LC_6_17_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i30_LC_6_17_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i30_LC_6_17_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i30_LC_6_17_1  (
            .in0(N__27174),
            .in1(N__45418),
            .in2(_gnd_net_),
            .in3(N__27199),
            .lcout(data_in_3_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50265),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15266_3_lut_LC_6_17_2 .C_ON=1'b0;
    defparam \c0.i15266_3_lut_LC_6_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.i15266_3_lut_LC_6_17_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.i15266_3_lut_LC_6_17_2  (
            .in0(N__27271),
            .in1(N__26977),
            .in2(_gnd_net_),
            .in3(N__27062),
            .lcout(),
            .ltout(\c0.n17715_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_941_LC_6_17_3 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_941_LC_6_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_941_LC_6_17_3 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \c0.i3_4_lut_adj_941_LC_6_17_3  (
            .in0(N__24370),
            .in1(N__27103),
            .in2(N__23654),
            .in3(N__23924),
            .lcout(\c0.n8_adj_2474 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16061_LC_6_17_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16061_LC_6_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16061_LC_6_17_4 .LUT_INIT=16'b1110010010101010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_16061_LC_6_17_4  (
            .in0(N__30770),
            .in1(N__25655),
            .in2(N__23651),
            .in3(N__31124),
            .lcout(\c0.n18540 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i32_LC_6_17_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i32_LC_6_17_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i32_LC_6_17_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i32_LC_6_17_5  (
            .in0(N__27232),
            .in1(N__45419),
            .in2(_gnd_net_),
            .in3(N__23946),
            .lcout(data_in_3_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50265),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i1_LC_6_17_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i1_LC_6_17_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i1_LC_6_17_6 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \c0.data_in_0___i1_LC_6_17_6  (
            .in0(N__23973),
            .in1(_gnd_net_),
            .in2(N__45484),
            .in3(N__24007),
            .lcout(\c0.data_in_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50265),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_940_LC_6_17_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_940_LC_6_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_940_LC_6_17_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i1_2_lut_adj_940_LC_6_17_7  (
            .in0(_gnd_net_),
            .in1(N__23969),
            .in2(_gnd_net_),
            .in3(N__23944),
            .lcout(\c0.n6_adj_2473 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i53_LC_6_18_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i53_LC_6_18_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i53_LC_6_18_1 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i53_LC_6_18_1  (
            .in0(N__27454),
            .in1(_gnd_net_),
            .in2(N__45485),
            .in3(N__27426),
            .lcout(\c0.data_in_6_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50279),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i65_LC_6_18_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i65_LC_6_18_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i65_LC_6_18_3 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i65_LC_6_18_3  (
            .in0(N__29419),
            .in1(_gnd_net_),
            .in2(N__45486),
            .in3(N__23893),
            .lcout(data_in_8_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50279),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i2_LC_6_18_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i2_LC_6_18_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i2_LC_6_18_5 .LUT_INIT=16'b0000110010101110;
    LogicCell40 \c0.data_out_frame2_0___i2_LC_6_18_5  (
            .in0(N__33158),
            .in1(N__31171),
            .in2(N__33693),
            .in3(N__23882),
            .lcout(\c0.data_out_frame2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50279),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3947_3_lut_LC_6_18_6 .C_ON=1'b0;
    defparam \c0.i3947_3_lut_LC_6_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3947_3_lut_LC_6_18_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.i3947_3_lut_LC_6_18_6  (
            .in0(N__23831),
            .in1(N__23804),
            .in2(_gnd_net_),
            .in3(N__24118),
            .lcout(n2599),
            .ltout(n2599_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_893_LC_6_18_7 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_893_LC_6_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_893_LC_6_18_7 .LUT_INIT=16'b1101111001111011;
    LogicCell40 \c0.i4_4_lut_adj_893_LC_6_18_7  (
            .in0(N__24560),
            .in1(N__28591),
            .in2(N__23756),
            .in3(N__27466),
            .lcout(\c0.n20_adj_2452 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_934_LC_6_19_0 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_934_LC_6_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_934_LC_6_19_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i5_4_lut_adj_934_LC_6_19_0  (
            .in0(N__27315),
            .in1(N__27536),
            .in2(N__31410),
            .in3(N__27707),
            .lcout(),
            .ltout(\c0.n12_adj_2472_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_937_LC_6_19_1 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_937_LC_6_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_937_LC_6_19_1 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \c0.i6_4_lut_adj_937_LC_6_19_1  (
            .in0(N__27680),
            .in1(N__23736),
            .in2(N__23720),
            .in3(N__23717),
            .lcout(\c0.n8556 ),
            .ltout(\c0.n8556_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_944_LC_6_19_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_944_LC_6_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_944_LC_6_19_2 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \c0.i1_2_lut_adj_944_LC_6_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24395),
            .in3(N__27740),
            .lcout(\c0.n6_adj_2478 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_LC_6_19_3 .C_ON=1'b0;
    defparam \c0.i2_2_lut_LC_6_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_LC_6_19_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i2_2_lut_LC_6_19_3  (
            .in0(_gnd_net_),
            .in1(N__27133),
            .in2(_gnd_net_),
            .in3(N__24343),
            .lcout(),
            .ltout(\c0.n7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_947_LC_6_19_4 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_947_LC_6_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_947_LC_6_19_4 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \c0.i4_4_lut_adj_947_LC_6_19_4  (
            .in0(N__28141),
            .in1(N__28183),
            .in2(N__24392),
            .in3(N__31378),
            .lcout(n63),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_946_LC_6_19_5 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_946_LC_6_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_946_LC_6_19_5 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \c0.i4_4_lut_adj_946_LC_6_19_5  (
            .in0(N__37652),
            .in1(N__27872),
            .in2(N__37553),
            .in3(N__24389),
            .lcout(\c0.n8460 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_956_LC_6_20_0 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_956_LC_6_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_956_LC_6_20_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i6_4_lut_adj_956_LC_6_20_0  (
            .in0(N__24379),
            .in1(N__27280),
            .in2(N__28117),
            .in3(N__24344),
            .lcout(),
            .ltout(\c0.n16_adj_2485_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_1010_LC_6_20_1 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_1010_LC_6_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_1010_LC_6_20_1 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \c0.i9_4_lut_adj_1010_LC_6_20_1  (
            .in0(N__27604),
            .in1(N__24332),
            .in2(N__24323),
            .in3(N__26951),
            .lcout(n63_adj_2642),
            .ltout(n63_adj_2642_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10279_3_lut_4_lut_LC_6_20_2 .C_ON=1'b0;
    defparam \c0.i10279_3_lut_4_lut_LC_6_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i10279_3_lut_4_lut_LC_6_20_2 .LUT_INIT=16'b1100111011000100;
    LogicCell40 \c0.i10279_3_lut_4_lut_LC_6_20_2  (
            .in0(N__34550),
            .in1(N__24317),
            .in2(N__24281),
            .in3(N__39845),
            .lcout(n2561),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_adj_1009_LC_6_20_3 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_adj_1009_LC_6_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_adj_1009_LC_6_20_3 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \c0.i2_2_lut_3_lut_adj_1009_LC_6_20_3  (
            .in0(N__34307),
            .in1(_gnd_net_),
            .in2(N__34408),
            .in3(N__34548),
            .lcout(n16468),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1011_LC_6_20_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1011_LC_6_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1011_LC_6_20_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_1011_LC_6_20_4  (
            .in0(_gnd_net_),
            .in1(N__34308),
            .in2(_gnd_net_),
            .in3(N__34367),
            .lcout(\c0.n4_adj_2512 ),
            .ltout(\c0.n4_adj_2512_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10772_3_lut_4_lut_LC_6_20_5 .C_ON=1'b0;
    defparam \c0.i10772_3_lut_4_lut_LC_6_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i10772_3_lut_4_lut_LC_6_20_5 .LUT_INIT=16'b1100101011001100;
    LogicCell40 \c0.i10772_3_lut_4_lut_LC_6_20_5  (
            .in0(N__24594),
            .in1(N__25472),
            .in2(N__24578),
            .in3(N__34549),
            .lcout(n2591),
            .ltout(n2591_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_902_LC_6_20_6 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_902_LC_6_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_902_LC_6_20_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_902_LC_6_20_6  (
            .in0(N__24555),
            .in1(N__24524),
            .in2(N__24506),
            .in3(N__24503),
            .lcout(\c0.n17533 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3959_3_lut_4_lut_LC_6_20_7 .C_ON=1'b0;
    defparam \c0.i3959_3_lut_4_lut_LC_6_20_7 .SEQ_MODE=4'b0000;
    defparam \c0.i3959_3_lut_4_lut_LC_6_20_7 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \c0.i3959_3_lut_4_lut_LC_6_20_7  (
            .in0(N__24763),
            .in1(N__34551),
            .in2(N__33037),
            .in3(N__28035),
            .lcout(\c0.n2605 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3889_3_lut_4_lut_LC_6_21_0 .C_ON=1'b0;
    defparam \c0.i3889_3_lut_4_lut_LC_6_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3889_3_lut_4_lut_LC_6_21_0 .LUT_INIT=16'b1101110010001100;
    LogicCell40 \c0.i3889_3_lut_4_lut_LC_6_21_0  (
            .in0(N__34394),
            .in1(N__36597),
            .in2(N__34642),
            .in3(N__32908),
            .lcout(n2570),
            .ltout(n2570_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i78_LC_6_21_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i78_LC_6_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i78_LC_6_21_1 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \c0.data_in_frame_0___i78_LC_6_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__24458),
            .in3(N__31907),
            .lcout(\c0.data_in_frame_9_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50295),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1013_LC_6_21_2 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1013_LC_6_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1013_LC_6_21_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i7_4_lut_adj_1013_LC_6_21_2  (
            .in0(N__24455),
            .in1(N__27904),
            .in2(N__28118),
            .in3(N__27140),
            .lcout(),
            .ltout(\c0.n17_adj_2514_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_1014_LC_6_21_3 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_1014_LC_6_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_1014_LC_6_21_3 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \c0.i9_4_lut_adj_1014_LC_6_21_3  (
            .in0(N__27741),
            .in1(N__27824),
            .in2(N__24446),
            .in3(N__37472),
            .lcout(FRAME_MATCHER_next_state_31_N_2026_1),
            .ltout(FRAME_MATCHER_next_state_31_N_2026_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3943_3_lut_4_lut_LC_6_21_4 .C_ON=1'b0;
    defparam \c0.i3943_3_lut_4_lut_LC_6_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3943_3_lut_4_lut_LC_6_21_4 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \c0.i3943_3_lut_4_lut_LC_6_21_4  (
            .in0(N__33061),
            .in1(N__24443),
            .in2(N__24419),
            .in3(N__28033),
            .lcout(n2597),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3883_3_lut_4_lut_LC_6_21_5 .C_ON=1'b0;
    defparam \c0.i3883_3_lut_4_lut_LC_6_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3883_3_lut_4_lut_LC_6_21_5 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \c0.i3883_3_lut_4_lut_LC_6_21_5  (
            .in0(N__29926),
            .in1(N__34594),
            .in2(N__25631),
            .in3(N__34393),
            .lcout(n2567),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_898_LC_6_21_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_898_LC_6_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_898_LC_6_21_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_898_LC_6_21_6  (
            .in0(N__25389),
            .in1(N__24879),
            .in2(_gnd_net_),
            .in3(N__24994),
            .lcout(\c0.n17575 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3961_3_lut_4_lut_LC_6_22_0 .C_ON=1'b0;
    defparam \c0.i3961_3_lut_4_lut_LC_6_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3961_3_lut_4_lut_LC_6_22_0 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \c0.i3961_3_lut_4_lut_LC_6_22_0  (
            .in0(N__28043),
            .in1(N__24971),
            .in2(N__39892),
            .in3(N__34575),
            .lcout(\c0.n2606 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3951_3_lut_4_lut_LC_6_22_1 .C_ON=1'b0;
    defparam \c0.i3951_3_lut_4_lut_LC_6_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3951_3_lut_4_lut_LC_6_22_1 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \c0.i3951_3_lut_4_lut_LC_6_22_1  (
            .in0(N__34574),
            .in1(N__28042),
            .in2(N__24692),
            .in3(N__31263),
            .lcout(),
            .ltout(\c0.n2601_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_968_LC_6_22_2 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_968_LC_6_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_968_LC_6_22_2 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \c0.i3_4_lut_adj_968_LC_6_22_2  (
            .in0(N__24791),
            .in1(N__24935),
            .in2(N__24911),
            .in3(N__24900),
            .lcout(\c0.n11_adj_2494 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_adj_1043_LC_6_22_3 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_adj_1043_LC_6_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_adj_1043_LC_6_22_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_adj_1043_LC_6_22_3  (
            .in0(N__25444),
            .in1(N__24883),
            .in2(N__25403),
            .in3(N__28196),
            .lcout(),
            .ltout(\c0.n17428_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_981_LC_6_22_4 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_981_LC_6_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_981_LC_6_22_4 .LUT_INIT=16'b1111111111110110;
    LogicCell40 \c0.i6_4_lut_adj_981_LC_6_22_4  (
            .in0(N__24848),
            .in1(N__24821),
            .in2(N__24815),
            .in3(N__24812),
            .lcout(\c0.n14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1058_LC_6_22_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1058_LC_6_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1058_LC_6_22_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1058_LC_6_22_5  (
            .in0(N__24678),
            .in1(N__24753),
            .in2(_gnd_net_),
            .in3(N__24790),
            .lcout(\c0.n9103 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_900_LC_6_22_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_900_LC_6_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_900_LC_6_22_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_900_LC_6_22_6  (
            .in0(N__24754),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24682),
            .lcout(\c0.n17430 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3955_3_lut_4_lut_LC_6_22_7 .C_ON=1'b0;
    defparam \c0.i3955_3_lut_4_lut_LC_6_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.i3955_3_lut_4_lut_LC_6_22_7 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \c0.i3955_3_lut_4_lut_LC_6_22_7  (
            .in0(N__34576),
            .in1(N__28044),
            .in2(N__27403),
            .in3(N__25277),
            .lcout(\c0.n2603 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3885_3_lut_4_lut_LC_6_23_0 .C_ON=1'b0;
    defparam \c0.i3885_3_lut_4_lut_LC_6_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3885_3_lut_4_lut_LC_6_23_0 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \c0.i3885_3_lut_4_lut_LC_6_23_0  (
            .in0(N__29828),
            .in1(N__34640),
            .in2(N__32263),
            .in3(N__34434),
            .lcout(n2568),
            .ltout(n2568_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_LC_6_23_1 .C_ON=1'b0;
    defparam \c0.i5_4_lut_LC_6_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_LC_6_23_1 .LUT_INIT=16'b1011111001111101;
    LogicCell40 \c0.i5_4_lut_LC_6_23_1  (
            .in0(N__25208),
            .in1(N__25189),
            .in2(N__25178),
            .in3(N__31450),
            .lcout(),
            .ltout(\c0.n21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_866_LC_6_23_2 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_866_LC_6_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_866_LC_6_23_2 .LUT_INIT=16'b1111110111111110;
    LogicCell40 \c0.i11_4_lut_adj_866_LC_6_23_2  (
            .in0(N__25174),
            .in1(N__27914),
            .in2(N__25145),
            .in3(N__32935),
            .lcout(),
            .ltout(\c0.n27_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_LC_6_23_3 .C_ON=1'b0;
    defparam \c0.i15_4_lut_LC_6_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_LC_6_23_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i15_4_lut_LC_6_23_3  (
            .in0(N__28781),
            .in1(N__25142),
            .in2(N__25136),
            .in3(N__28499),
            .lcout(\c0.n5_adj_2438 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3897_3_lut_4_lut_LC_6_23_4 .C_ON=1'b0;
    defparam \c0.i3897_3_lut_4_lut_LC_6_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3897_3_lut_4_lut_LC_6_23_4 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \c0.i3897_3_lut_4_lut_LC_6_23_4  (
            .in0(N__27657),
            .in1(N__34641),
            .in2(N__36741),
            .in3(N__34433),
            .lcout(n2574),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i74_LC_6_23_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i74_LC_6_23_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i74_LC_6_23_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i74_LC_6_23_5  (
            .in0(N__45344),
            .in1(N__29531),
            .in2(_gnd_net_),
            .in3(N__27658),
            .lcout(data_in_9_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50311),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1119_LC_6_24_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1119_LC_6_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1119_LC_6_24_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1119_LC_6_24_1  (
            .in0(_gnd_net_),
            .in1(N__28098),
            .in2(_gnd_net_),
            .in3(N__25108),
            .lcout(\c0.n4_adj_2548 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_1131_LC_6_24_2.C_ON=1'b0;
    defparam i1_2_lut_adj_1131_LC_6_24_2.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_1131_LC_6_24_2.LUT_INIT=16'b0101010110101010;
    LogicCell40 i1_2_lut_adj_1131_LC_6_24_2 (
            .in0(N__28099),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25063),
            .lcout(n19_adj_2651),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i35_LC_6_24_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i35_LC_6_24_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i35_LC_6_24_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i35_LC_6_24_3  (
            .in0(N__45280),
            .in1(N__29844),
            .in2(_gnd_net_),
            .in3(N__33027),
            .lcout(data_in_4_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50318),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_LC_6_24_4.C_ON=1'b0;
    defparam i1_2_lut_LC_6_24_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_LC_6_24_4.LUT_INIT=16'b0011001111001100;
    LogicCell40 i1_2_lut_LC_6_24_4 (
            .in0(_gnd_net_),
            .in1(N__25588),
            .in2(_gnd_net_),
            .in3(N__28439),
            .lcout(),
            .ltout(n6_adj_2604_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i4_4_lut_LC_6_24_5.C_ON=1'b0;
    defparam i4_4_lut_LC_6_24_5.SEQ_MODE=4'b0000;
    defparam i4_4_lut_LC_6_24_5.LUT_INIT=16'b0110100110010110;
    LogicCell40 i4_4_lut_LC_6_24_5 (
            .in0(N__25529),
            .in1(N__25501),
            .in2(N__25475),
            .in3(N__25471),
            .lcout(n17547),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_adj_1046_LC_6_24_6 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_adj_1046_LC_6_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_adj_1046_LC_6_24_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_adj_1046_LC_6_24_6  (
            .in0(N__25443),
            .in1(N__29762),
            .in2(N__25399),
            .in3(N__25361),
            .lcout(\c0.n8666 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i114_LC_6_24_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i114_LC_6_24_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i114_LC_6_24_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i114_LC_6_24_7  (
            .in0(N__35356),
            .in1(N__25309),
            .in2(_gnd_net_),
            .in3(N__32815),
            .lcout(data_out_frame2_14_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50318),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i0_LC_6_25_1 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i0_LC_6_25_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i0_LC_6_25_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.tx.r_Clock_Count__i0_LC_6_25_1  (
            .in0(N__40371),
            .in1(N__25295),
            .in2(_gnd_net_),
            .in3(N__29660),
            .lcout(r_Clock_Count_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50328),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i13_LC_6_25_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i13_LC_6_25_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i13_LC_6_25_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_0___i13_LC_6_25_2  (
            .in0(N__27326),
            .in1(N__37648),
            .in2(_gnd_net_),
            .in3(N__45245),
            .lcout(data_in_1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50328),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i4_LC_6_25_3 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i4_LC_6_25_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i4_LC_6_25_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.tx.r_Clock_Count__i4_LC_6_25_3  (
            .in0(N__40372),
            .in1(N__29603),
            .in2(_gnd_net_),
            .in3(N__25289),
            .lcout(r_Clock_Count_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50328),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i3_LC_6_25_4 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i3_LC_6_25_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i3_LC_6_25_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.tx.r_Clock_Count__i3_LC_6_25_4  (
            .in0(N__29621),
            .in1(N__25283),
            .in2(_gnd_net_),
            .in3(N__40374),
            .lcout(r_Clock_Count_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50328),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i60_LC_6_25_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i60_LC_6_25_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i60_LC_6_25_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_0___i60_LC_6_25_6  (
            .in0(N__25710),
            .in1(N__29734),
            .in2(_gnd_net_),
            .in3(N__45246),
            .lcout(data_in_7_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50328),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i5_LC_6_25_7 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i5_LC_6_25_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i5_LC_6_25_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.tx.r_Clock_Count__i5_LC_6_25_7  (
            .in0(N__40373),
            .in1(N__25694),
            .in2(_gnd_net_),
            .in3(N__29641),
            .lcout(r_Clock_Count_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50328),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i9_3_lut_LC_6_26_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i9_3_lut_LC_6_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i9_3_lut_LC_6_26_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_4_i9_3_lut_LC_6_26_0  (
            .in0(N__25688),
            .in1(N__25669),
            .in2(_gnd_net_),
            .in3(N__30753),
            .lcout(\c0.n9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i123_LC_6_26_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i123_LC_6_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i123_LC_6_26_1 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i123_LC_6_26_1  (
            .in0(N__34049),
            .in1(_gnd_net_),
            .in2(N__45347),
            .in3(N__29881),
            .lcout(data_in_15_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50337),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i61_LC_6_26_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i61_LC_6_26_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i61_LC_6_26_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_out_frame2_0___i61_LC_6_26_2  (
            .in0(N__30235),
            .in1(N__35662),
            .in2(_gnd_net_),
            .in3(N__32823),
            .lcout(data_out_frame2_7_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50337),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i80_LC_6_26_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i80_LC_6_26_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i80_LC_6_26_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i80_LC_6_26_3  (
            .in0(N__45238),
            .in1(N__29826),
            .in2(_gnd_net_),
            .in3(N__30472),
            .lcout(data_in_9_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50337),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i118_LC_6_26_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i118_LC_6_26_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i118_LC_6_26_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i118_LC_6_26_4  (
            .in0(N__36099),
            .in1(N__25651),
            .in2(_gnd_net_),
            .in3(N__32822),
            .lcout(data_out_frame2_14_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50337),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i165_LC_6_26_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i165_LC_6_26_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i165_LC_6_26_5 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \c0.data_in_0___i165_LC_6_26_5  (
            .in0(N__38443),
            .in1(_gnd_net_),
            .in2(N__45348),
            .in3(N__29896),
            .lcout(data_in_20_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50337),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_953_LC_6_26_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_953_LC_6_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_953_LC_6_26_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_953_LC_6_26_6  (
            .in0(_gnd_net_),
            .in1(N__29258),
            .in2(_gnd_net_),
            .in3(N__25635),
            .lcout(\c0.n17559 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i11212_2_lut_LC_6_26_7 .C_ON=1'b0;
    defparam \c0.rx.i11212_2_lut_LC_6_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i11212_2_lut_LC_6_26_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.rx.i11212_2_lut_LC_6_26_7  (
            .in0(_gnd_net_),
            .in1(N__39245),
            .in2(_gnd_net_),
            .in3(N__39307),
            .lcout(n13597),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i107_LC_6_27_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i107_LC_6_27_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i107_LC_6_27_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i107_LC_6_27_0  (
            .in0(N__45226),
            .in1(N__34705),
            .in2(_gnd_net_),
            .in3(N__29870),
            .lcout(data_in_13_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50347),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i4_LC_6_27_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i4_LC_6_27_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i4_LC_6_27_2 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \c0.data_out_frame2_0___i4_LC_6_27_2  (
            .in0(N__33645),
            .in1(N__25810),
            .in2(_gnd_net_),
            .in3(N__25790),
            .lcout(\c0.data_out_frame2_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50347),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i100_LC_6_27_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i100_LC_6_27_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i100_LC_6_27_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_out_frame2_0___i100_LC_6_27_3  (
            .in0(N__25778),
            .in1(N__35204),
            .in2(_gnd_net_),
            .in3(N__32832),
            .lcout(data_out_frame2_12_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50347),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i51_LC_6_27_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i51_LC_6_27_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i51_LC_6_27_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_0___i51_LC_6_27_5  (
            .in0(N__33060),
            .in1(N__33763),
            .in2(_gnd_net_),
            .in3(N__45231),
            .lcout(data_in_6_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50347),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i155_LC_6_27_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i155_LC_6_27_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i155_LC_6_27_6 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i155_LC_6_27_6  (
            .in0(N__25766),
            .in1(_gnd_net_),
            .in2(N__45345),
            .in3(N__38464),
            .lcout(data_in_19_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50347),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i163_LC_6_27_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i163_LC_6_27_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i163_LC_6_27_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i163_LC_6_27_7  (
            .in0(N__30014),
            .in1(N__45227),
            .in2(_gnd_net_),
            .in3(N__25765),
            .lcout(data_in_20_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50347),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15930_LC_6_28_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15930_LC_6_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15930_LC_6_28_1 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_15930_LC_6_28_1  (
            .in0(N__26663),
            .in1(N__25757),
            .in2(N__25751),
            .in3(N__26846),
            .lcout(),
            .ltout(\c0.n18372_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18372_bdd_4_lut_LC_6_28_2 .C_ON=1'b0;
    defparam \c0.n18372_bdd_4_lut_LC_6_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.n18372_bdd_4_lut_LC_6_28_2 .LUT_INIT=16'b1111000011001010;
    LogicCell40 \c0.n18372_bdd_4_lut_LC_6_28_2  (
            .in0(N__25796),
            .in1(N__25742),
            .in2(N__25730),
            .in3(N__26664),
            .lcout(),
            .ltout(\c0.n18375_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i3_LC_6_28_3 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i3_LC_6_28_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i3_LC_6_28_3 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \c0.tx2.r_Tx_Data_i3_LC_6_28_3  (
            .in0(N__26665),
            .in1(N__25949),
            .in2(N__26054),
            .in3(N__26521),
            .lcout(\c0.tx2.r_Tx_Data_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50357),
            .ce(N__26416),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16036_LC_6_28_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16036_LC_6_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16036_LC_6_28_4 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_16036_LC_6_28_4  (
            .in0(N__26039),
            .in1(N__31076),
            .in2(N__26021),
            .in3(N__30789),
            .lcout(),
            .ltout(\c0.n18510_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18510_bdd_4_lut_LC_6_28_5 .C_ON=1'b0;
    defparam \c0.n18510_bdd_4_lut_LC_6_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.n18510_bdd_4_lut_LC_6_28_5 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n18510_bdd_4_lut_LC_6_28_5  (
            .in0(N__31077),
            .in1(N__26003),
            .in2(N__25985),
            .in3(N__25982),
            .lcout(),
            .ltout(\c0.n18513_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_3_i22_4_lut_LC_6_28_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_3_i22_4_lut_LC_6_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_3_i22_4_lut_LC_6_28_6 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_3_i22_4_lut_LC_6_28_6  (
            .in0(N__26845),
            .in1(N__25964),
            .in2(N__25952),
            .in3(N__26925),
            .lcout(\c0.n22_adj_2527 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Bit_Index_i2_LC_6_29_0 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_i2_LC_6_29_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Bit_Index_i2_LC_6_29_0 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \c0.tx2.r_Bit_Index_i2_LC_6_29_0  (
            .in0(N__25871),
            .in1(N__25943),
            .in2(N__26093),
            .in3(N__25910),
            .lcout(r_Bit_Index_2_adj_2635),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50368),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i153_LC_6_29_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i153_LC_6_29_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i153_LC_6_29_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i153_LC_6_29_1  (
            .in0(N__45232),
            .in1(N__37823),
            .in2(_gnd_net_),
            .in3(N__29938),
            .lcout(data_in_19_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50368),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i1_LC_6_29_3 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i1_LC_6_29_3 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i1_LC_6_29_3 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \c0.rx.r_Clock_Count__i1_LC_6_29_3  (
            .in0(N__26081),
            .in1(N__30375),
            .in2(N__29969),
            .in3(N__30316),
            .lcout(r_Clock_Count_1_adj_2623),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50368),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_955_LC_6_29_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_955_LC_6_29_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_955_LC_6_29_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_955_LC_6_29_4  (
            .in0(N__31516),
            .in1(N__32065),
            .in2(N__25847),
            .in3(N__28534),
            .lcout(n9135),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15817_3_lut_LC_6_29_5 .C_ON=1'b0;
    defparam \c0.i15817_3_lut_LC_6_29_5 .SEQ_MODE=4'b0000;
    defparam \c0.i15817_3_lut_LC_6_29_5 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \c0.i15817_3_lut_LC_6_29_5  (
            .in0(N__30790),
            .in1(N__25811),
            .in2(_gnd_net_),
            .in3(N__31123),
            .lcout(\c0.n18082 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i2450_2_lut_LC_6_29_7 .C_ON=1'b0;
    defparam \c0.tx2.i2450_2_lut_LC_6_29_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i2450_2_lut_LC_6_29_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.tx2.i2450_2_lut_LC_6_29_7  (
            .in0(N__26186),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26135),
            .lcout(n4980),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_2_lut_LC_6_30_0 .C_ON=1'b1;
    defparam \c0.rx.add_62_2_lut_LC_6_30_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_2_lut_LC_6_30_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.add_62_2_lut_LC_6_30_0  (
            .in0(_gnd_net_),
            .in1(N__29988),
            .in2(_gnd_net_),
            .in3(N__26084),
            .lcout(n226),
            .ltout(),
            .carryin(bfn_6_30_0_),
            .carryout(\c0.rx.n16365 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_3_lut_LC_6_30_1 .C_ON=1'b1;
    defparam \c0.rx.add_62_3_lut_LC_6_30_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_3_lut_LC_6_30_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.add_62_3_lut_LC_6_30_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29965),
            .in3(N__26075),
            .lcout(n225),
            .ltout(),
            .carryin(\c0.rx.n16365 ),
            .carryout(\c0.rx.n16366 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_4_lut_LC_6_30_2 .C_ON=1'b1;
    defparam \c0.rx.add_62_4_lut_LC_6_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_4_lut_LC_6_30_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.add_62_4_lut_LC_6_30_2  (
            .in0(_gnd_net_),
            .in1(N__30110),
            .in2(_gnd_net_),
            .in3(N__26072),
            .lcout(n224),
            .ltout(),
            .carryin(\c0.rx.n16366 ),
            .carryout(\c0.rx.n16367 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_5_lut_LC_6_30_3 .C_ON=1'b1;
    defparam \c0.rx.add_62_5_lut_LC_6_30_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_5_lut_LC_6_30_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.add_62_5_lut_LC_6_30_3  (
            .in0(_gnd_net_),
            .in1(N__30070),
            .in2(_gnd_net_),
            .in3(N__26069),
            .lcout(n223),
            .ltout(),
            .carryin(\c0.rx.n16367 ),
            .carryout(\c0.rx.n16368 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_6_lut_LC_6_30_4 .C_ON=1'b1;
    defparam \c0.rx.add_62_6_lut_LC_6_30_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_6_lut_LC_6_30_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.add_62_6_lut_LC_6_30_4  (
            .in0(_gnd_net_),
            .in1(N__30334),
            .in2(_gnd_net_),
            .in3(N__26066),
            .lcout(n222),
            .ltout(),
            .carryin(\c0.rx.n16368 ),
            .carryout(\c0.rx.n16369 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_7_lut_LC_6_30_5 .C_ON=1'b1;
    defparam \c0.rx.add_62_7_lut_LC_6_30_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_7_lut_LC_6_30_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.add_62_7_lut_LC_6_30_5  (
            .in0(_gnd_net_),
            .in1(N__38101),
            .in2(_gnd_net_),
            .in3(N__26063),
            .lcout(n221),
            .ltout(),
            .carryin(\c0.rx.n16369 ),
            .carryout(\c0.rx.n16370 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_8_lut_LC_6_30_6 .C_ON=1'b1;
    defparam \c0.rx.add_62_8_lut_LC_6_30_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_8_lut_LC_6_30_6 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.rx.add_62_8_lut_LC_6_30_6  (
            .in0(N__30119),
            .in1(N__37998),
            .in2(_gnd_net_),
            .in3(N__26060),
            .lcout(\c0.rx.n18001 ),
            .ltout(),
            .carryin(\c0.rx.n16370 ),
            .carryout(\c0.rx.n16371 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.add_62_9_lut_LC_6_30_7 .C_ON=1'b0;
    defparam \c0.rx.add_62_9_lut_LC_6_30_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.add_62_9_lut_LC_6_30_7 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \c0.rx.add_62_9_lut_LC_6_30_7  (
            .in0(N__38055),
            .in1(N__30118),
            .in2(_gnd_net_),
            .in3(N__26057),
            .lcout(\c0.rx.n17999 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i2_LC_6_31_0 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i2_LC_6_31_0 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i2_LC_6_31_0 .LUT_INIT=16'b0000000010101100;
    LogicCell40 \c0.rx.r_Clock_Count__i2_LC_6_31_0  (
            .in0(N__30108),
            .in1(N__26318),
            .in2(N__30317),
            .in3(N__30376),
            .lcout(r_Clock_Count_2_adj_2622),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50384),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i0_LC_6_31_1 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i0_LC_6_31_1 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i0_LC_6_31_1 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \c0.rx.r_Clock_Count__i0_LC_6_31_1  (
            .in0(N__26306),
            .in1(N__30373),
            .in2(N__29993),
            .in3(N__30310),
            .lcout(r_Clock_Count_0_adj_2624),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50384),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i5_LC_6_31_2 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i5_LC_6_31_2 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i5_LC_6_31_2 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \c0.rx.r_Clock_Count__i5_LC_6_31_2  (
            .in0(N__30315),
            .in1(N__30377),
            .in2(N__38110),
            .in3(N__26300),
            .lcout(r_Clock_Count_5_adj_2619),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50384),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i3_LC_6_31_3 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i3_LC_6_31_3 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i3_LC_6_31_3 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \c0.rx.r_Clock_Count__i3_LC_6_31_3  (
            .in0(N__26294),
            .in1(N__30374),
            .in2(N__30074),
            .in3(N__30314),
            .lcout(r_Clock_Count_3_adj_2621),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50384),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i11152_2_lut_LC_6_31_5 .C_ON=1'b0;
    defparam \c0.rx.i11152_2_lut_LC_6_31_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i11152_2_lut_LC_6_31_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.rx.i11152_2_lut_LC_6_31_5  (
            .in0(_gnd_net_),
            .in1(N__30107),
            .in2(_gnd_net_),
            .in3(N__30068),
            .lcout(\c0.rx.n13537 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i7_LC_6_31_6 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i7_LC_6_31_6 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i7_LC_6_31_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.rx.r_Clock_Count__i7_LC_6_31_6  (
            .in0(N__30309),
            .in1(N__38056),
            .in2(_gnd_net_),
            .in3(N__26288),
            .lcout(\c0.rx.r_Clock_Count_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50384),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18444_bdd_4_lut_LC_6_31_7 .C_ON=1'b0;
    defparam \c0.n18444_bdd_4_lut_LC_6_31_7 .SEQ_MODE=4'b0000;
    defparam \c0.n18444_bdd_4_lut_LC_6_31_7 .LUT_INIT=16'b1010101011011000;
    LogicCell40 \c0.n18444_bdd_4_lut_LC_6_31_7  (
            .in0(N__26282),
            .in1(N__26273),
            .in2(N__31190),
            .in3(N__26842),
            .lcout(\c0.n18447 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16051_LC_6_32_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16051_LC_6_32_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_16051_LC_6_32_0 .LUT_INIT=16'b1110010010101010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_16051_LC_6_32_0  (
            .in0(N__30795),
            .in1(N__26264),
            .in2(N__26243),
            .in3(N__31155),
            .lcout(),
            .ltout(\c0.n18528_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18528_bdd_4_lut_LC_6_32_1 .C_ON=1'b0;
    defparam \c0.n18528_bdd_4_lut_LC_6_32_1 .SEQ_MODE=4'b0000;
    defparam \c0.n18528_bdd_4_lut_LC_6_32_1 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n18528_bdd_4_lut_LC_6_32_1  (
            .in0(N__31156),
            .in1(N__26225),
            .in2(N__26207),
            .in3(N__26204),
            .lcout(),
            .ltout(\c0.n18531_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i22_4_lut_LC_6_32_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i22_4_lut_LC_6_32_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i22_4_lut_LC_6_32_2 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_4_i22_4_lut_LC_6_32_2  (
            .in0(N__29294),
            .in1(N__26934),
            .in2(N__26870),
            .in3(N__26798),
            .lcout(\c0.n22_adj_2525 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15709_2_lut_LC_6_32_3 .C_ON=1'b0;
    defparam \c0.i15709_2_lut_LC_6_32_3 .SEQ_MODE=4'b0000;
    defparam \c0.i15709_2_lut_LC_6_32_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i15709_2_lut_LC_6_32_3  (
            .in0(_gnd_net_),
            .in1(N__26867),
            .in2(_gnd_net_),
            .in3(N__30796),
            .lcout(),
            .ltout(\c0.n17955_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_1__bdd_4_lut_LC_6_32_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_1__bdd_4_lut_LC_6_32_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_1__bdd_4_lut_LC_6_32_4 .LUT_INIT=16'b1011100011001100;
    LogicCell40 \c0.byte_transmit_counter2_1__bdd_4_lut_LC_6_32_4  (
            .in0(N__30200),
            .in1(N__31157),
            .in2(N__26849),
            .in3(N__26799),
            .lcout(),
            .ltout(\c0.n18456_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18456_bdd_4_lut_4_lut_LC_6_32_5 .C_ON=1'b0;
    defparam \c0.n18456_bdd_4_lut_4_lut_LC_6_32_5 .SEQ_MODE=4'b0000;
    defparam \c0.n18456_bdd_4_lut_4_lut_LC_6_32_5 .LUT_INIT=16'b1111000010100100;
    LogicCell40 \c0.n18456_bdd_4_lut_4_lut_LC_6_32_5  (
            .in0(N__26800),
            .in1(N__26714),
            .in2(N__26696),
            .in3(N__30797),
            .lcout(),
            .ltout(\c0.n18459_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11600217_i1_3_lut_LC_6_32_6 .C_ON=1'b0;
    defparam \c0.i11600217_i1_3_lut_LC_6_32_6 .SEQ_MODE=4'b0000;
    defparam \c0.i11600217_i1_3_lut_LC_6_32_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \c0.i11600217_i1_3_lut_LC_6_32_6  (
            .in0(_gnd_net_),
            .in1(N__26693),
            .in2(N__26687),
            .in3(N__26666),
            .lcout(),
            .ltout(\c0.n15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i4_LC_6_32_7 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i4_LC_6_32_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i4_LC_6_32_7 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \c0.tx2.r_Tx_Data_i4_LC_6_32_7  (
            .in0(N__26684),
            .in1(N__26678),
            .in2(N__26528),
            .in3(N__26525),
            .lcout(\c0.tx2.r_Tx_Data_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50391),
            .ce(N__26404),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i29_LC_7_17_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i29_LC_7_17_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i29_LC_7_17_0 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i29_LC_7_17_0  (
            .in0(N__27364),
            .in1(_gnd_net_),
            .in2(N__45483),
            .in3(N__27895),
            .lcout(\c0.data_in_3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50272),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i2_LC_7_17_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i2_LC_7_17_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i2_LC_7_17_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_0___i2_LC_7_17_1  (
            .in0(N__27073),
            .in1(N__31377),
            .in2(_gnd_net_),
            .in3(N__45416),
            .lcout(data_in_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50272),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i22_LC_7_17_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i22_LC_7_17_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i22_LC_7_17_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i22_LC_7_17_2  (
            .in0(N__45410),
            .in1(N__27175),
            .in2(_gnd_net_),
            .in3(N__26985),
            .lcout(data_in_2_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50272),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i17_LC_7_17_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i17_LC_7_17_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i17_LC_7_17_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_0___i17_LC_7_17_3  (
            .in0(N__27111),
            .in1(N__27835),
            .in2(_gnd_net_),
            .in3(N__45415),
            .lcout(\c0.data_in_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50272),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i16_LC_7_17_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i16_LC_7_17_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i16_LC_7_17_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i16_LC_7_17_4  (
            .in0(N__45409),
            .in1(N__27032),
            .in2(_gnd_net_),
            .in3(N__27276),
            .lcout(data_in_1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50272),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i40_LC_7_17_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i40_LC_7_17_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i40_LC_7_17_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_0___i40_LC_7_17_5  (
            .in0(N__36916),
            .in1(N__27231),
            .in2(_gnd_net_),
            .in3(N__45417),
            .lcout(data_in_4_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50272),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i38_LC_7_17_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i38_LC_7_17_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i38_LC_7_17_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i38_LC_7_17_7  (
            .in0(N__29557),
            .in1(N__45411),
            .in2(_gnd_net_),
            .in3(N__27198),
            .lcout(data_in_4_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50272),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i46_2_lut_LC_7_18_0 .C_ON=1'b0;
    defparam \c0.i46_2_lut_LC_7_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.i46_2_lut_LC_7_18_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i46_2_lut_LC_7_18_0  (
            .in0(_gnd_net_),
            .in1(N__27596),
            .in2(_gnd_net_),
            .in3(N__27022),
            .lcout(),
            .ltout(\c0.n28_adj_2475_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_943_LC_7_18_1 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_943_LC_7_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_943_LC_7_18_1 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \c0.i1_4_lut_adj_943_LC_7_18_1  (
            .in0(N__27789),
            .in1(N__27172),
            .in2(N__27149),
            .in3(N__27146),
            .lcout(\c0.n8559 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_957_LC_7_18_2 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_957_LC_7_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_957_LC_7_18_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i7_4_lut_adj_957_LC_7_18_2  (
            .in0(N__27104),
            .in1(N__27063),
            .in2(N__27033),
            .in3(N__26978),
            .lcout(\c0.n17_adj_2486 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i20_LC_7_18_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i20_LC_7_18_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i20_LC_7_18_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i20_LC_7_18_3  (
            .in0(N__37552),
            .in1(N__45430),
            .in2(_gnd_net_),
            .in3(N__27538),
            .lcout(data_in_2_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50284),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i82_LC_7_18_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i82_LC_7_18_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i82_LC_7_18_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i82_LC_7_18_4  (
            .in0(N__45429),
            .in1(N__31316),
            .in2(_gnd_net_),
            .in3(N__29523),
            .lcout(data_in_10_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50284),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i4_LC_7_18_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i4_LC_7_18_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i4_LC_7_18_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i4_LC_7_18_5  (
            .in0(N__27597),
            .in1(N__45432),
            .in2(_gnd_net_),
            .in3(N__27644),
            .lcout(\c0.data_in_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50284),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i28_LC_7_18_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i28_LC_7_18_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i28_LC_7_18_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i28_LC_7_18_7  (
            .in0(N__27571),
            .in1(N__45431),
            .in2(_gnd_net_),
            .in3(N__27537),
            .lcout(data_in_3_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50284),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3923_3_lut_4_lut_LC_7_19_0 .C_ON=1'b0;
    defparam \c0.i3923_3_lut_4_lut_LC_7_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3923_3_lut_4_lut_LC_7_19_0 .LUT_INIT=16'b1010101011100010;
    LogicCell40 \c0.i3923_3_lut_4_lut_LC_7_19_0  (
            .in0(N__27517),
            .in1(N__34643),
            .in2(N__27455),
            .in3(N__28034),
            .lcout(n2587),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i61_LC_7_19_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i61_LC_7_19_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i61_LC_7_19_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i61_LC_7_19_1  (
            .in0(N__45329),
            .in1(N__38377),
            .in2(_gnd_net_),
            .in3(N__27453),
            .lcout(\c0.data_in_7_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50289),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i45_LC_7_19_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i45_LC_7_19_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i45_LC_7_19_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i45_LC_7_19_3  (
            .in0(N__27427),
            .in1(N__45295),
            .in2(_gnd_net_),
            .in3(N__27390),
            .lcout(data_in_5_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50289),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i37_LC_7_19_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i37_LC_7_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i37_LC_7_19_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i37_LC_7_19_4  (
            .in0(N__27389),
            .in1(N__45330),
            .in2(_gnd_net_),
            .in3(N__27357),
            .lcout(\c0.data_in_4_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50289),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i7_LC_7_19_5 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i7_LC_7_19_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i7_LC_7_19_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.tx.r_Clock_Count__i7_LC_7_19_5  (
            .in0(N__40375),
            .in1(N__27341),
            .in2(_gnd_net_),
            .in3(N__37199),
            .lcout(r_Clock_Count_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50289),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i21_LC_7_19_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i21_LC_7_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i21_LC_7_19_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i21_LC_7_19_6  (
            .in0(N__45294),
            .in1(N__27897),
            .in2(_gnd_net_),
            .in3(N__27314),
            .lcout(data_in_2_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50289),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15294_4_lut_LC_7_19_7 .C_ON=1'b0;
    defparam \c0.i15294_4_lut_LC_7_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.i15294_4_lut_LC_7_19_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i15294_4_lut_LC_7_19_7  (
            .in0(N__27896),
            .in1(N__27823),
            .in2(N__37612),
            .in3(N__37508),
            .lcout(\c0.n17743 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i25_LC_7_20_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i25_LC_7_20_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i25_LC_7_20_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_0___i25_LC_7_20_0  (
            .in0(N__27831),
            .in1(N__27866),
            .in2(_gnd_net_),
            .in3(N__45452),
            .lcout(\c0.data_in_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50296),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i7_LC_7_20_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i7_LC_7_20_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i7_LC_7_20_1 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i7_LC_7_20_1  (
            .in0(N__27796),
            .in1(_gnd_net_),
            .in2(N__45494),
            .in3(N__27742),
            .lcout(data_in_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50296),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i23_LC_7_20_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i23_LC_7_20_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i23_LC_7_20_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_0___i23_LC_7_20_2  (
            .in0(N__27714),
            .in1(N__28182),
            .in2(_gnd_net_),
            .in3(N__45451),
            .lcout(data_in_2_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50296),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13622_3_lut_4_lut_LC_7_20_3 .C_ON=1'b0;
    defparam \c0.i13622_3_lut_4_lut_LC_7_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i13622_3_lut_4_lut_LC_7_20_3 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \c0.i13622_3_lut_4_lut_LC_7_20_3  (
            .in0(N__38348),
            .in1(N__34606),
            .in2(N__31505),
            .in3(N__34426),
            .lcout(n2571),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i73_LC_7_20_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i73_LC_7_20_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i73_LC_7_20_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_0___i73_LC_7_20_4  (
            .in0(N__29927),
            .in1(N__29412),
            .in2(_gnd_net_),
            .in3(N__45453),
            .lcout(data_in_9_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50296),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i26_LC_7_20_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i26_LC_7_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i26_LC_7_20_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i26_LC_7_20_5  (
            .in0(N__45445),
            .in1(N__38506),
            .in2(_gnd_net_),
            .in3(N__27681),
            .lcout(data_in_3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50296),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i18_LC_7_20_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i18_LC_7_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i18_LC_7_20_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i18_LC_7_20_6  (
            .in0(N__27682),
            .in1(N__45447),
            .in2(_gnd_net_),
            .in3(N__31409),
            .lcout(data_in_2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50296),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i66_LC_7_20_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i66_LC_7_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i66_LC_7_20_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i66_LC_7_20_7  (
            .in0(N__45446),
            .in1(N__37032),
            .in2(_gnd_net_),
            .in3(N__27662),
            .lcout(data_in_8_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50296),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_828_LC_7_21_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_828_LC_7_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_828_LC_7_21_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_828_LC_7_21_0  (
            .in0(_gnd_net_),
            .in1(N__28493),
            .in2(_gnd_net_),
            .in3(N__28434),
            .lcout(\c0.n17473 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i31_LC_7_21_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i31_LC_7_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i31_LC_7_21_1 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \c0.data_in_0___i31_LC_7_21_1  (
            .in0(_gnd_net_),
            .in1(N__45346),
            .in2(N__28385),
            .in3(N__28181),
            .lcout(data_in_3_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50303),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3949_3_lut_4_lut_LC_7_21_2 .C_ON=1'b0;
    defparam \c0.i3949_3_lut_4_lut_LC_7_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3949_3_lut_4_lut_LC_7_21_2 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \c0.i3949_3_lut_4_lut_LC_7_21_2  (
            .in0(N__28343),
            .in1(N__34572),
            .in2(N__36912),
            .in3(N__28023),
            .lcout(),
            .ltout(\c0.n2600_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_966_LC_7_21_3 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_966_LC_7_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_966_LC_7_21_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_966_LC_7_21_3  (
            .in0(N__28274),
            .in1(N__28262),
            .in2(N__28220),
            .in3(N__28216),
            .lcout(\c0.n10_adj_2493 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_932_LC_7_21_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_932_LC_7_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_932_LC_7_21_5 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \c0.i2_3_lut_adj_932_LC_7_21_5  (
            .in0(N__28174),
            .in1(N__31376),
            .in2(_gnd_net_),
            .in3(N__28148),
            .lcout(\c0.n8572 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3937_3_lut_4_lut_LC_7_21_6 .C_ON=1'b0;
    defparam \c0.i3937_3_lut_4_lut_LC_7_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3937_3_lut_4_lut_LC_7_21_6 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \c0.i3937_3_lut_4_lut_LC_7_21_6  (
            .in0(N__28100),
            .in1(N__34573),
            .in2(N__36190),
            .in3(N__28024),
            .lcout(n2594),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i84_LC_7_21_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i84_LC_7_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i84_LC_7_21_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.data_in_frame_0___i84_LC_7_21_7  (
            .in0(_gnd_net_),
            .in1(N__31451),
            .in2(_gnd_net_),
            .in3(N__31972),
            .lcout(\c0.data_in_frame_10_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50303),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10244_3_lut_4_lut_LC_7_22_0 .C_ON=1'b0;
    defparam \c0.i10244_3_lut_4_lut_LC_7_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10244_3_lut_4_lut_LC_7_22_0 .LUT_INIT=16'b1110111101000000;
    LogicCell40 \c0.i10244_3_lut_4_lut_LC_7_22_0  (
            .in0(N__34436),
            .in1(N__36493),
            .in2(N__34644),
            .in3(N__32106),
            .lcout(n2573),
            .ltout(n2573_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_3_lut_4_lut_adj_1156_LC_7_22_1.C_ON=1'b0;
    defparam i2_3_lut_4_lut_adj_1156_LC_7_22_1.SEQ_MODE=4'b0000;
    defparam i2_3_lut_4_lut_adj_1156_LC_7_22_1.LUT_INIT=16'b0110100110010110;
    LogicCell40 i2_3_lut_4_lut_adj_1156_LC_7_22_1 (
            .in0(N__29173),
            .in1(N__28774),
            .in2(N__27917),
            .in3(N__28732),
            .lcout(n17481),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1122_LC_7_22_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1122_LC_7_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1122_LC_7_22_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1122_LC_7_22_2  (
            .in0(N__28978),
            .in1(N__28933),
            .in2(N__28646),
            .in3(N__28895),
            .lcout(\c0.n17536 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3879_3_lut_4_lut_LC_7_22_3 .C_ON=1'b0;
    defparam \c0.i3879_3_lut_4_lut_LC_7_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3879_3_lut_4_lut_LC_7_22_3 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \c0.i3879_3_lut_4_lut_LC_7_22_3  (
            .in0(N__36524),
            .in1(N__34601),
            .in2(N__32057),
            .in3(N__34435),
            .lcout(n2565),
            .ltout(n2565_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_LC_7_22_4 .C_ON=1'b0;
    defparam \c0.i7_4_lut_LC_7_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_LC_7_22_4 .LUT_INIT=16'b1101011111101011;
    LogicCell40 \c0.i7_4_lut_LC_7_22_4  (
            .in0(N__28873),
            .in1(N__28849),
            .in2(N__28829),
            .in3(N__28819),
            .lcout(),
            .ltout(\c0.n23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_862_LC_7_22_5 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_862_LC_7_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_862_LC_7_22_5 .LUT_INIT=16'b1111100111111111;
    LogicCell40 \c0.i12_4_lut_adj_862_LC_7_22_5  (
            .in0(N__28807),
            .in1(N__31537),
            .in2(N__28790),
            .in3(N__28787),
            .lcout(\c0.n28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_1130_LC_7_22_7.C_ON=1'b0;
    defparam i1_2_lut_adj_1130_LC_7_22_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_1130_LC_7_22_7.LUT_INIT=16'b0011001111001100;
    LogicCell40 i1_2_lut_adj_1130_LC_7_22_7 (
            .in0(_gnd_net_),
            .in1(N__28775),
            .in2(_gnd_net_),
            .in3(N__28733),
            .lcout(n17479),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3875_3_lut_4_lut_LC_7_23_0 .C_ON=1'b0;
    defparam \c0.i3875_3_lut_4_lut_LC_7_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3875_3_lut_4_lut_LC_7_23_0 .LUT_INIT=16'b1101110010001100;
    LogicCell40 \c0.i3875_3_lut_4_lut_LC_7_23_0  (
            .in0(N__34455),
            .in1(N__28679),
            .in2(N__34661),
            .in3(N__38330),
            .lcout(n2563),
            .ltout(n2563_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1118_LC_7_23_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1118_LC_7_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1118_LC_7_23_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1118_LC_7_23_1  (
            .in0(N__28641),
            .in1(N__28595),
            .in2(N__28568),
            .in3(N__28564),
            .lcout(),
            .ltout(\c0.n17592_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_LC_7_23_2 .C_ON=1'b0;
    defparam \c0.i10_4_lut_LC_7_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_LC_7_23_2 .LUT_INIT=16'b1111111111110110;
    LogicCell40 \c0.i10_4_lut_LC_7_23_2  (
            .in0(N__28535),
            .in1(N__29344),
            .in2(N__28502),
            .in3(N__29429),
            .lcout(\c0.n26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3881_3_lut_4_lut_LC_7_23_3 .C_ON=1'b0;
    defparam \c0.i3881_3_lut_4_lut_LC_7_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3881_3_lut_4_lut_LC_7_23_3 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \c0.i3881_3_lut_4_lut_LC_7_23_3  (
            .in0(N__29530),
            .in1(N__34622),
            .in2(N__36871),
            .in3(N__34454),
            .lcout(n2566),
            .ltout(n2566_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_841_LC_7_23_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_841_LC_7_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_841_LC_7_23_4 .LUT_INIT=16'b1101011111101011;
    LogicCell40 \c0.i3_4_lut_adj_841_LC_7_23_4  (
            .in0(N__29507),
            .in1(N__29480),
            .in2(N__29453),
            .in3(N__29446),
            .lcout(\c0.n19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3899_3_lut_4_lut_LC_7_23_5 .C_ON=1'b0;
    defparam \c0.i3899_3_lut_4_lut_LC_7_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3899_3_lut_4_lut_LC_7_23_5 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \c0.i3899_3_lut_4_lut_LC_7_23_5  (
            .in0(N__29423),
            .in1(N__34626),
            .in2(N__29388),
            .in3(N__34456),
            .lcout(n2575),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1091_LC_7_24_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1091_LC_7_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1091_LC_7_24_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1091_LC_7_24_0  (
            .in0(_gnd_net_),
            .in1(N__29246),
            .in2(_gnd_net_),
            .in3(N__36691),
            .lcout(),
            .ltout(\c0.n6_adj_2541_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i165_LC_7_24_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i165_LC_7_24_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i165_LC_7_24_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_frame2_0___i165_LC_7_24_1  (
            .in0(N__29333),
            .in1(N__29269),
            .in2(N__29312),
            .in3(N__29309),
            .lcout(\c0.data_out_frame2_20_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50329),
            .ce(N__32841),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_LC_7_24_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_LC_7_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_LC_7_24_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_LC_7_24_2  (
            .in0(N__32110),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31512),
            .lcout(\c0.n17488 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i155_LC_7_24_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i155_LC_7_24_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i155_LC_7_24_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_frame2_0___i155_LC_7_24_5  (
            .in0(N__29247),
            .in1(N__29210),
            .in2(N__29201),
            .in3(N__29177),
            .lcout(\c0.data_out_frame2_19_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50329),
            .ce(N__32841),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1059_LC_7_24_6 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1059_LC_7_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1059_LC_7_24_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1059_LC_7_24_6  (
            .in0(N__29138),
            .in1(N__29093),
            .in2(N__29060),
            .in3(N__29012),
            .lcout(\c0.n10_adj_2536 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i1_LC_7_25_0 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i1_LC_7_25_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i1_LC_7_25_0 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.tx.r_Clock_Count__i1_LC_7_25_0  (
            .in0(N__29578),
            .in1(_gnd_net_),
            .in2(N__40370),
            .in3(N__29756),
            .lcout(r_Clock_Count_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50338),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i68_LC_7_25_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i68_LC_7_25_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i68_LC_7_25_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i68_LC_7_25_1  (
            .in0(N__45250),
            .in1(N__29733),
            .in2(_gnd_net_),
            .in3(N__29677),
            .lcout(data_in_8_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50338),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_2_lut_LC_7_25_3 .C_ON=1'b0;
    defparam \c0.tx.i1_2_lut_LC_7_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_2_lut_LC_7_25_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.tx.i1_2_lut_LC_7_25_3  (
            .in0(_gnd_net_),
            .in1(N__40155),
            .in2(_gnd_net_),
            .in3(N__40350),
            .lcout(),
            .ltout(n8517_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_1138_LC_7_25_4.C_ON=1'b0;
    defparam i1_4_lut_adj_1138_LC_7_25_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_1138_LC_7_25_4.LUT_INIT=16'b0000000011011100;
    LogicCell40 i1_4_lut_adj_1138_LC_7_25_4 (
            .in0(N__33086),
            .in1(N__37346),
            .in2(N__29717),
            .in3(N__33852),
            .lcout(n17366),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i76_LC_7_25_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i76_LC_7_25_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i76_LC_7_25_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \c0.data_in_0___i76_LC_7_25_5  (
            .in0(N__45251),
            .in1(_gnd_net_),
            .in2(N__36989),
            .in3(N__29676),
            .lcout(data_in_9_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50338),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i4_4_lut_LC_7_25_6 .C_ON=1'b0;
    defparam \c0.tx.i4_4_lut_LC_7_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i4_4_lut_LC_7_25_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.tx.i4_4_lut_LC_7_25_6  (
            .in0(N__33789),
            .in1(N__29658),
            .in2(N__29642),
            .in3(N__29619),
            .lcout(),
            .ltout(\c0.tx.n10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i5_3_lut_LC_7_25_7 .C_ON=1'b0;
    defparam \c0.tx.i5_3_lut_LC_7_25_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i5_3_lut_LC_7_25_7 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \c0.tx.i5_3_lut_LC_7_25_7  (
            .in0(_gnd_net_),
            .in1(N__29601),
            .in2(N__29585),
            .in3(N__29577),
            .lcout(n16466),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i46_LC_7_26_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i46_LC_7_26_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i46_LC_7_26_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_0___i46_LC_7_26_0  (
            .in0(N__29553),
            .in1(N__36191),
            .in2(_gnd_net_),
            .in3(N__45248),
            .lcout(data_in_5_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50348),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i69_LC_7_26_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i69_LC_7_26_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i69_LC_7_26_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i69_LC_7_26_2  (
            .in0(N__35153),
            .in1(N__31204),
            .in2(_gnd_net_),
            .in3(N__32652),
            .lcout(data_out_frame2_8_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50348),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i6_LC_7_26_4 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i6_LC_7_26_4 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i6_LC_7_26_4 .LUT_INIT=16'b1111110100001000;
    LogicCell40 \c0.rx.r_Rx_Byte_i6_LC_7_26_4  (
            .in0(N__33724),
            .in1(N__37909),
            .in2(N__37946),
            .in3(N__33709),
            .lcout(rx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50348),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i145_LC_7_26_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i145_LC_7_26_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i145_LC_7_26_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i145_LC_7_26_5  (
            .in0(N__45247),
            .in1(N__37453),
            .in2(_gnd_net_),
            .in3(N__29942),
            .lcout(data_in_18_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50348),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i81_LC_7_26_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i81_LC_7_26_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i81_LC_7_26_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_0___i81_LC_7_26_6  (
            .in0(N__29919),
            .in1(N__36785),
            .in2(_gnd_net_),
            .in3(N__45249),
            .lcout(data_in_10_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50348),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i4_LC_7_26_7 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i4_LC_7_26_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i4_LC_7_26_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.rx.r_Rx_Byte_i4_LC_7_26_7  (
            .in0(N__33976),
            .in1(N__37941),
            .in2(N__29897),
            .in3(N__37910),
            .lcout(rx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50348),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i115_LC_7_27_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i115_LC_7_27_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i115_LC_7_27_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i115_LC_7_27_1  (
            .in0(N__45066),
            .in1(N__29869),
            .in2(_gnd_net_),
            .in3(N__29882),
            .lcout(data_in_14_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50358),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i136_LC_7_27_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i136_LC_7_27_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i136_LC_7_27_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i136_LC_7_27_2  (
            .in0(N__45077),
            .in1(N__30406),
            .in2(_gnd_net_),
            .in3(N__31472),
            .lcout(data_in_16_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50358),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i27_LC_7_27_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i27_LC_7_27_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i27_LC_7_27_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i27_LC_7_27_3  (
            .in0(N__45067),
            .in1(N__29851),
            .in2(_gnd_net_),
            .in3(N__37507),
            .lcout(data_in_3_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50358),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i72_LC_7_27_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i72_LC_7_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i72_LC_7_27_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_0___i72_LC_7_27_4  (
            .in0(N__29827),
            .in1(N__29784),
            .in2(_gnd_net_),
            .in3(N__45068),
            .lcout(data_in_8_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50358),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_4_lut_LC_7_28_0 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_4_lut_LC_7_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_4_lut_LC_7_28_0 .LUT_INIT=16'b1111111110111111;
    LogicCell40 \c0.rx.i1_2_lut_4_lut_LC_7_28_0  (
            .in0(N__30139),
            .in1(N__39654),
            .in2(N__40459),
            .in3(N__39584),
            .lcout(n8567),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i105_LC_7_28_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i105_LC_7_28_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i105_LC_7_28_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i105_LC_7_28_3  (
            .in0(N__35949),
            .in1(N__30040),
            .in2(_gnd_net_),
            .in3(N__32843),
            .lcout(data_out_frame2_13_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50369),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i150_LC_7_28_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i150_LC_7_28_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i150_LC_7_28_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i150_LC_7_28_4  (
            .in0(N__45233),
            .in1(N__30025),
            .in2(_gnd_net_),
            .in3(N__37721),
            .lcout(data_in_18_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50369),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i142_LC_7_28_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i142_LC_7_28_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i142_LC_7_28_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i142_LC_7_28_5  (
            .in0(N__30026),
            .in1(N__45234),
            .in2(_gnd_net_),
            .in3(N__34264),
            .lcout(data_in_17_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50369),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_4_lut_adj_820_LC_7_28_6 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_4_lut_adj_820_LC_7_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_4_lut_adj_820_LC_7_28_6 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \c0.rx.i1_2_lut_4_lut_adj_820_LC_7_28_6  (
            .in0(N__30140),
            .in1(N__39655),
            .in2(N__40460),
            .in3(N__39585),
            .lcout(n8562),
            .ltout(n8562_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i2_LC_7_28_7 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i2_LC_7_28_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i2_LC_7_28_7 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \c0.rx.r_Rx_Byte_i2_LC_7_28_7  (
            .in0(N__34033),
            .in1(N__30013),
            .in2(N__30017),
            .in3(N__37894),
            .lcout(rx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50369),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_3_lut_4_lut_LC_7_29_0 .C_ON=1'b0;
    defparam \c0.rx.i2_3_lut_4_lut_LC_7_29_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_3_lut_4_lut_LC_7_29_0 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \c0.rx.i2_3_lut_4_lut_LC_7_29_0  (
            .in0(N__39687),
            .in1(N__39556),
            .in2(N__37895),
            .in3(N__34245),
            .lcout(\c0.rx.n2 ),
            .ltout(\c0.rx.n2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_4_lut_adj_818_LC_7_29_1 .C_ON=1'b0;
    defparam \c0.rx.i1_4_lut_adj_818_LC_7_29_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_4_lut_adj_818_LC_7_29_1 .LUT_INIT=16'b0000001100000010;
    LogicCell40 \c0.rx.i1_4_lut_adj_818_LC_7_29_1  (
            .in0(N__39521),
            .in1(N__39752),
            .in2(N__30002),
            .in3(N__30383),
            .lcout(\c0.rx.n4_adj_2424 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_adj_819_LC_7_29_2 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_adj_819_LC_7_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_adj_819_LC_7_29_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \c0.rx.i1_2_lut_adj_819_LC_7_29_2  (
            .in0(N__39754),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29999),
            .lcout(n3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_3_lut_LC_7_29_3 .C_ON=1'b0;
    defparam \c0.rx.i2_3_lut_LC_7_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_3_lut_LC_7_29_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.rx.i2_3_lut_LC_7_29_3  (
            .in0(N__30333),
            .in1(N__29992),
            .in2(_gnd_net_),
            .in3(N__29958),
            .lcout(\c0.rx.n124 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_i1_LC_7_29_4 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_i1_LC_7_29_4 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_SM_Main_i1_LC_7_29_4 .LUT_INIT=16'b0000010000001110;
    LogicCell40 \c0.rx.r_SM_Main_i1_LC_7_29_4  (
            .in0(N__39690),
            .in1(N__34232),
            .in2(N__39771),
            .in3(N__30194),
            .lcout(\c0.rx.r_SM_Main_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50376),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.n18594_bdd_4_lut_4_lut_LC_7_29_5 .C_ON=1'b0;
    defparam \c0.rx.n18594_bdd_4_lut_4_lut_LC_7_29_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.n18594_bdd_4_lut_4_lut_LC_7_29_5 .LUT_INIT=16'b1111000010100011;
    LogicCell40 \c0.rx.n18594_bdd_4_lut_4_lut_LC_7_29_5  (
            .in0(N__34246),
            .in1(N__37876),
            .in2(N__38297),
            .in3(N__39689),
            .lcout(\c0.rx.n18597 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Data_50_LC_7_29_6 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Data_50_LC_7_29_6 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Data_50_LC_7_29_6 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \c0.rx.r_Rx_Data_50_LC_7_29_6  (
            .in0(_gnd_net_),
            .in1(N__30173),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(r_Rx_Data),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50376),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_adj_816_LC_7_29_7 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_adj_816_LC_7_29_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_adj_816_LC_7_29_7 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \c0.rx.i1_2_lut_adj_816_LC_7_29_7  (
            .in0(_gnd_net_),
            .in1(N__39753),
            .in2(_gnd_net_),
            .in3(N__39688),
            .lcout(\c0.rx.n17381 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_4_lut_LC_7_30_0 .C_ON=1'b0;
    defparam \c0.rx.i2_4_lut_LC_7_30_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_4_lut_LC_7_30_0 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \c0.rx.i2_4_lut_LC_7_30_0  (
            .in0(N__30250),
            .in1(N__30085),
            .in2(N__38106),
            .in3(N__30157),
            .lcout(\c0.rx.r_SM_Main_2_N_2386_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i15740_4_lut_LC_7_30_1 .C_ON=1'b0;
    defparam \c0.rx.i15740_4_lut_LC_7_30_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i15740_4_lut_LC_7_30_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.rx.i15740_4_lut_LC_7_30_1  (
            .in0(N__30158),
            .in1(N__38096),
            .in2(N__30089),
            .in3(N__30148),
            .lcout(),
            .ltout(\c0.rx.n18003_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i57_4_lut_LC_7_30_2 .C_ON=1'b0;
    defparam \c0.rx.i57_4_lut_LC_7_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i57_4_lut_LC_7_30_2 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.rx.i57_4_lut_LC_7_30_2  (
            .in0(N__30149),
            .in1(N__30138),
            .in2(N__30125),
            .in3(N__30251),
            .lcout(n13880),
            .ltout(n13880_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i7678_1_lut_LC_7_30_3 .C_ON=1'b0;
    defparam \c0.rx.i7678_1_lut_LC_7_30_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i7678_1_lut_LC_7_30_3 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \c0.rx.i7678_1_lut_LC_7_30_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30122),
            .in3(_gnd_net_),
            .lcout(\c0.rx.n10193 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_3_lut_adj_813_LC_7_30_4 .C_ON=1'b0;
    defparam \c0.rx.i2_3_lut_adj_813_LC_7_30_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_3_lut_adj_813_LC_7_30_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.rx.i2_3_lut_adj_813_LC_7_30_4  (
            .in0(N__30109),
            .in1(N__30084),
            .in2(_gnd_net_),
            .in3(N__30069),
            .lcout(\c0.rx.n97 ),
            .ltout(\c0.rx.n97_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_4_lut_adj_817_LC_7_30_5 .C_ON=1'b0;
    defparam \c0.rx.i1_4_lut_adj_817_LC_7_30_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_4_lut_adj_817_LC_7_30_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \c0.rx.i1_4_lut_adj_817_LC_7_30_5  (
            .in0(N__38100),
            .in1(N__38054),
            .in2(N__30386),
            .in3(N__37997),
            .lcout(\c0.rx.n17345 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i4_LC_7_30_6 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i4_LC_7_30_6 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i4_LC_7_30_6 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \c0.rx.r_Clock_Count__i4_LC_7_30_6  (
            .in0(N__30294),
            .in1(N__30372),
            .in2(N__30341),
            .in3(N__30347),
            .lcout(r_Clock_Count_4_adj_2620),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50385),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i6_LC_7_30_7 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i6_LC_7_30_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i6_LC_7_30_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.rx.r_Clock_Count__i6_LC_7_30_7  (
            .in0(N__37999),
            .in1(N__30293),
            .in2(_gnd_net_),
            .in3(N__30278),
            .lcout(\c0.rx.r_Clock_Count_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50385),
            .ce(),
            .sr(_gnd_net_));
    defparam i15405_4_lut_LC_7_31_0.C_ON=1'b0;
    defparam i15405_4_lut_LC_7_31_0.SEQ_MODE=4'b0000;
    defparam i15405_4_lut_LC_7_31_0.LUT_INIT=16'b1111001000110000;
    LogicCell40 i15405_4_lut_LC_7_31_0 (
            .in0(N__49063),
            .in1(N__49039),
            .in2(N__49112),
            .in3(N__49087),
            .lcout(n17855),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15406_4_lut_LC_7_31_1.C_ON=1'b0;
    defparam i15406_4_lut_LC_7_31_1.SEQ_MODE=4'b0000;
    defparam i15406_4_lut_LC_7_31_1.LUT_INIT=16'b1111110111001000;
    LogicCell40 i15406_4_lut_LC_7_31_1 (
            .in0(N__49088),
            .in1(N__49111),
            .in2(N__49043),
            .in3(N__49064),
            .lcout(),
            .ltout(n17856_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15407_3_lut_LC_7_31_2.C_ON=1'b0;
    defparam i15407_3_lut_LC_7_31_2.SEQ_MODE=4'b0000;
    defparam i15407_3_lut_LC_7_31_2.LUT_INIT=16'b0000101001011111;
    LogicCell40 i15407_3_lut_LC_7_31_2 (
            .in0(N__50459),
            .in1(_gnd_net_),
            .in2(N__30272),
            .in3(N__30269),
            .lcout(LED_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_i2_LC_7_31_3 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_i2_LC_7_31_3 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_SM_Main_i2_LC_7_31_3 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \c0.rx.r_SM_Main_i2_LC_7_31_3  (
            .in0(N__38102),
            .in1(N__38050),
            .in2(N__38020),
            .in3(N__37993),
            .lcout(\c0.rx.r_SM_Main_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50392),
            .ce(),
            .sr(N__39608));
    defparam \c0.rx.i1_2_lut_adj_814_LC_7_31_5 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_adj_814_LC_7_31_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_adj_814_LC_7_31_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.rx.i1_2_lut_adj_814_LC_7_31_5  (
            .in0(_gnd_net_),
            .in1(N__38049),
            .in2(_gnd_net_),
            .in3(N__37992),
            .lcout(\c0.rx.n112 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i5_3_lut_LC_7_31_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i5_3_lut_LC_7_31_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i5_3_lut_LC_7_31_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_4_i5_3_lut_LC_7_31_6  (
            .in0(N__30239),
            .in1(N__30221),
            .in2(_gnd_net_),
            .in3(N__30794),
            .lcout(\c0.n5_adj_2425 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i8_3_lut_LC_7_31_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i8_3_lut_LC_7_31_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i8_3_lut_LC_7_31_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_4_i8_3_lut_LC_7_31_7  (
            .in0(N__30793),
            .in1(N__31226),
            .in2(_gnd_net_),
            .in3(N__31205),
            .lcout(\c0.n8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15708_3_lut_LC_7_32_0 .C_ON=1'b0;
    defparam \c0.i15708_3_lut_LC_7_32_0 .SEQ_MODE=4'b0000;
    defparam \c0.i15708_3_lut_LC_7_32_0 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \c0.i15708_3_lut_LC_7_32_0  (
            .in0(N__31181),
            .in1(N__31154),
            .in2(_gnd_net_),
            .in3(N__30792),
            .lcout(\c0.n18086 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i88_LC_7_32_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i88_LC_7_32_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i88_LC_7_32_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i88_LC_7_32_1  (
            .in0(N__30446),
            .in1(N__44937),
            .in2(_gnd_net_),
            .in3(N__30462),
            .lcout(data_in_10_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50397),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i96_LC_7_32_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i96_LC_7_32_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i96_LC_7_32_2 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i96_LC_7_32_2  (
            .in0(N__30437),
            .in1(_gnd_net_),
            .in2(N__45153),
            .in3(N__30445),
            .lcout(data_in_11_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50397),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i104_LC_7_32_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i104_LC_7_32_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i104_LC_7_32_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i104_LC_7_32_3  (
            .in0(N__30428),
            .in1(N__44935),
            .in2(_gnd_net_),
            .in3(N__30436),
            .lcout(data_in_12_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50397),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i112_LC_7_32_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i112_LC_7_32_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i112_LC_7_32_4 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i112_LC_7_32_4  (
            .in0(N__30419),
            .in1(_gnd_net_),
            .in2(N__45152),
            .in3(N__30427),
            .lcout(data_in_13_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50397),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i120_LC_7_32_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i120_LC_7_32_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i120_LC_7_32_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i120_LC_7_32_5  (
            .in0(N__30395),
            .in1(N__44936),
            .in2(_gnd_net_),
            .in3(N__30418),
            .lcout(data_in_14_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50397),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i128_LC_7_32_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i128_LC_7_32_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i128_LC_7_32_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i128_LC_7_32_6  (
            .in0(N__44934),
            .in1(N__30394),
            .in2(_gnd_net_),
            .in3(N__30410),
            .lcout(data_in_15_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50397),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i114_LC_9_18_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i114_LC_9_18_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i114_LC_9_18_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i114_LC_9_18_0  (
            .in0(N__45433),
            .in1(N__31429),
            .in2(_gnd_net_),
            .in3(N__36761),
            .lcout(data_in_14_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50297),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_next_state_i1_LC_9_19_3 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_next_state_i1_LC_9_19_3 .SEQ_MODE=4'b1000;
    defparam \c0.FRAME_MATCHER_next_state_i1_LC_9_19_3 .LUT_INIT=16'b1010001010101010;
    LogicCell40 \c0.FRAME_MATCHER_next_state_i1_LC_9_19_3  (
            .in0(N__34683),
            .in1(N__34453),
            .in2(N__33548),
            .in3(N__34318),
            .lcout(FRAME_MATCHER_next_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50304),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3877_3_lut_4_lut_LC_9_20_0 .C_ON=1'b0;
    defparam \c0.i3877_3_lut_4_lut_LC_9_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3877_3_lut_4_lut_LC_9_20_0 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \c0.i3877_3_lut_4_lut_LC_9_20_0  (
            .in0(N__36978),
            .in1(N__34662),
            .in2(N__36836),
            .in3(N__34447),
            .lcout(n2564),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i106_LC_9_20_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i106_LC_9_20_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i106_LC_9_20_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_0___i106_LC_9_20_1  (
            .in0(N__31333),
            .in1(N__31433),
            .in2(_gnd_net_),
            .in3(N__45350),
            .lcout(data_in_13_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50312),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i10_LC_9_20_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i10_LC_9_20_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i10_LC_9_20_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_0___i10_LC_9_20_3  (
            .in0(N__31414),
            .in1(N__31363),
            .in2(_gnd_net_),
            .in3(N__45351),
            .lcout(data_in_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50312),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i102_LC_9_20_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i102_LC_9_20_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i102_LC_9_20_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i102_LC_9_20_4  (
            .in0(N__45349),
            .in1(N__38615),
            .in2(_gnd_net_),
            .in3(N__32869),
            .lcout(data_in_12_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50312),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i98_LC_9_20_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i98_LC_9_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i98_LC_9_20_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_0___i98_LC_9_20_5  (
            .in0(N__31334),
            .in1(N__31324),
            .in2(_gnd_net_),
            .in3(N__45352),
            .lcout(data_in_12_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50312),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i90_LC_9_20_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i90_LC_9_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i90_LC_9_20_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i90_LC_9_20_6  (
            .in0(N__31325),
            .in1(N__45353),
            .in2(_gnd_net_),
            .in3(N__31309),
            .lcout(data_in_11_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50312),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i47_LC_9_21_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i47_LC_9_21_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i47_LC_9_21_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i47_LC_9_21_0  (
            .in0(N__45253),
            .in1(N__31247),
            .in2(_gnd_net_),
            .in3(N__31298),
            .lcout(data_in_5_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50319),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i64_LC_9_21_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i64_LC_9_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i64_LC_9_21_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i64_LC_9_21_1  (
            .in0(N__35474),
            .in1(N__32278),
            .in2(_gnd_net_),
            .in3(N__32827),
            .lcout(data_out_frame2_7_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50319),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_935_LC_9_21_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_935_LC_9_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_935_LC_9_21_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_935_LC_9_21_2  (
            .in0(N__36857),
            .in1(N__32246),
            .in2(_gnd_net_),
            .in3(N__36831),
            .lcout(\c0.n17433 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i56_LC_9_21_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i56_LC_9_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i56_LC_9_21_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_0___i56_LC_9_21_3  (
            .in0(N__36948),
            .in1(N__32165),
            .in2(_gnd_net_),
            .in3(N__45254),
            .lcout(data_in_6_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50319),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i75_LC_9_21_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i75_LC_9_21_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i75_LC_9_21_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \c0.data_in_frame_0___i75_LC_9_21_4  (
            .in0(_gnd_net_),
            .in1(N__31969),
            .in2(_gnd_net_),
            .in3(N__32126),
            .lcout(\c0.data_in_frame_9_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50319),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i83_LC_9_21_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i83_LC_9_21_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i83_LC_9_21_5 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \c0.data_in_frame_0___i83_LC_9_21_5  (
            .in0(N__31971),
            .in1(N__32078),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.data_in_frame_10_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50319),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i82_LC_9_21_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i82_LC_9_21_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i82_LC_9_21_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \c0.data_in_frame_0___i82_LC_9_21_6  (
            .in0(_gnd_net_),
            .in1(N__31968),
            .in2(_gnd_net_),
            .in3(N__32009),
            .lcout(\c0.data_in_frame_10_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50319),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0___i77_LC_9_21_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0___i77_LC_9_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0___i77_LC_9_21_7 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \c0.data_in_frame_0___i77_LC_9_21_7  (
            .in0(N__31970),
            .in1(N__31541),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.data_in_frame_9_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50319),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i164_LC_9_22_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i164_LC_9_22_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i164_LC_9_22_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i164_LC_9_22_0  (
            .in0(N__45155),
            .in1(N__33998),
            .in2(_gnd_net_),
            .in3(N__38626),
            .lcout(data_in_20_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50330),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i144_LC_9_22_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i144_LC_9_22_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i144_LC_9_22_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i144_LC_9_22_4  (
            .in0(N__45154),
            .in1(N__31462),
            .in2(_gnd_net_),
            .in3(N__37133),
            .lcout(data_in_17_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50330),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Done_44_LC_9_22_5 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Done_44_LC_9_22_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Done_44_LC_9_22_5 .LUT_INIT=16'b1011111110111000;
    LogicCell40 \c0.tx.r_Tx_Done_44_LC_9_22_5  (
            .in0(N__33077),
            .in1(N__36767),
            .in2(N__40369),
            .in3(N__32849),
            .lcout(n7364),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50330),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i43_LC_9_22_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i43_LC_9_22_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i43_LC_9_22_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \c0.data_in_0___i43_LC_9_22_6  (
            .in0(N__45156),
            .in1(_gnd_net_),
            .in2(N__33071),
            .in3(N__33014),
            .lcout(data_in_5_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50330),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3873_3_lut_4_lut_LC_9_23_0 .C_ON=1'b0;
    defparam \c0.i3873_3_lut_4_lut_LC_9_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3873_3_lut_4_lut_LC_9_23_0 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \c0.i3873_3_lut_4_lut_LC_9_23_0  (
            .in0(N__34679),
            .in1(N__32919),
            .in2(N__32986),
            .in3(N__34448),
            .lcout(n2562),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i79_LC_9_23_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i79_LC_9_23_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i79_LC_9_23_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_0___i79_LC_9_23_1  (
            .in0(N__39844),
            .in1(N__38790),
            .in2(_gnd_net_),
            .in3(N__45163),
            .lcout(data_in_9_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50339),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i86_LC_9_23_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i86_LC_9_23_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i86_LC_9_23_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i86_LC_9_23_2  (
            .in0(N__45160),
            .in1(N__32858),
            .in2(_gnd_net_),
            .in3(N__32920),
            .lcout(data_in_10_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50339),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i78_LC_9_23_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i78_LC_9_23_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i78_LC_9_23_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i78_LC_9_23_3  (
            .in0(N__32921),
            .in1(N__45162),
            .in2(_gnd_net_),
            .in3(N__32892),
            .lcout(data_in_9_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50339),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i94_LC_9_23_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i94_LC_9_23_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i94_LC_9_23_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i94_LC_9_23_4  (
            .in0(N__45161),
            .in1(N__32857),
            .in2(_gnd_net_),
            .in3(N__32873),
            .lcout(data_in_11_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50339),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i15809_2_lut_3_lut_LC_9_23_5 .C_ON=1'b0;
    defparam \c0.tx.i15809_2_lut_3_lut_LC_9_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i15809_2_lut_3_lut_LC_9_23_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.tx.i15809_2_lut_3_lut_LC_9_23_5  (
            .in0(N__40159),
            .in1(N__40403),
            .in2(_gnd_net_),
            .in3(N__40215),
            .lcout(n18098),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i4717_4_lut_LC_9_23_7 .C_ON=1'b0;
    defparam \c0.tx.i4717_4_lut_LC_9_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i4717_4_lut_LC_9_23_7 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \c0.tx.i4717_4_lut_LC_9_23_7  (
            .in0(N__42979),
            .in1(N__37280),
            .in2(N__40163),
            .in3(N__40402),
            .lcout(n7080),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_220_Select_0_i1_2_lut_4_lut_LC_9_24_0 .C_ON=1'b0;
    defparam \c0.select_220_Select_0_i1_2_lut_4_lut_LC_9_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.select_220_Select_0_i1_2_lut_4_lut_LC_9_24_0 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \c0.select_220_Select_0_i1_2_lut_4_lut_LC_9_24_0  (
            .in0(N__33267),
            .in1(N__34289),
            .in2(N__33388),
            .in3(N__33460),
            .lcout(\c0.n1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i0_LC_9_24_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i0_LC_9_24_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i0_LC_9_24_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \c0.FRAME_MATCHER_state_i0_LC_9_24_1  (
            .in0(N__33461),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33682),
            .lcout(\c0.FRAME_MATCHER_state_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50349),
            .ce(),
            .sr(N__33560));
    defparam \c0.select_220_Select_1_i1_2_lut_4_lut_LC_9_24_2 .C_ON=1'b0;
    defparam \c0.select_220_Select_1_i1_2_lut_4_lut_LC_9_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.select_220_Select_1_i1_2_lut_4_lut_LC_9_24_2 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \c0.select_220_Select_1_i1_2_lut_4_lut_LC_9_24_2  (
            .in0(N__33268),
            .in1(N__33547),
            .in2(N__33389),
            .in3(N__33459),
            .lcout(\c0.n1_adj_2437 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_2_lut_4_lut_adj_826_LC_9_24_4 .C_ON=1'b0;
    defparam \c0.tx.i1_2_lut_4_lut_adj_826_LC_9_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_2_lut_4_lut_adj_826_LC_9_24_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.tx.i1_2_lut_4_lut_adj_826_LC_9_24_4  (
            .in0(N__37321),
            .in1(N__37215),
            .in2(N__37261),
            .in3(N__33860),
            .lcout(r_SM_Main_2_N_2323_1),
            .ltout(r_SM_Main_2_N_2323_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i15308_4_lut_LC_9_24_5 .C_ON=1'b0;
    defparam \c0.tx.i15308_4_lut_LC_9_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i15308_4_lut_LC_9_24_5 .LUT_INIT=16'b1111111111001110;
    LogicCell40 \c0.tx.i15308_4_lut_LC_9_24_5  (
            .in0(N__40145),
            .in1(N__40339),
            .in2(N__33395),
            .in3(N__40213),
            .lcout(n17757),
            .ltout(n17757_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9716_4_lut_LC_9_24_6.C_ON=1'b0;
    defparam i9716_4_lut_LC_9_24_6.SEQ_MODE=4'b0000;
    defparam i9716_4_lut_LC_9_24_6.LUT_INIT=16'b1111010000001000;
    LogicCell40 i9716_4_lut_LC_9_24_6 (
            .in0(N__39126),
            .in1(N__37442),
            .in2(N__33392),
            .in3(N__37395),
            .lcout(n12123),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1048_LC_9_24_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1048_LC_9_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1048_LC_9_24_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \c0.i1_2_lut_adj_1048_LC_9_24_7  (
            .in0(_gnd_net_),
            .in1(N__33380),
            .in2(_gnd_net_),
            .in3(N__33266),
            .lcout(\c0.n157 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i6_LC_9_25_0 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i6_LC_9_25_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i6_LC_9_25_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.tx.r_Clock_Count__i6_LC_9_25_0  (
            .in0(N__40325),
            .in1(N__33098),
            .in2(_gnd_net_),
            .in3(N__37254),
            .lcout(r_Clock_Count_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50359),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i2_2_lut_4_lut_LC_9_25_1 .C_ON=1'b0;
    defparam \c0.tx.i2_2_lut_4_lut_LC_9_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i2_2_lut_4_lut_LC_9_25_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.tx.i2_2_lut_4_lut_LC_9_25_1  (
            .in0(N__37253),
            .in1(N__37315),
            .in2(N__40237),
            .in3(N__37222),
            .lcout(n9390),
            .ltout(n9390_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15234_3_lut_4_lut_LC_9_25_2.C_ON=1'b0;
    defparam i15234_3_lut_4_lut_LC_9_25_2.SEQ_MODE=4'b0000;
    defparam i15234_3_lut_4_lut_LC_9_25_2.LUT_INIT=16'b1011101111111011;
    LogicCell40 i15234_3_lut_4_lut_LC_9_25_2 (
            .in0(N__40324),
            .in1(N__40102),
            .in2(N__33866),
            .in3(N__37362),
            .lcout(),
            .ltout(n17681_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15277_4_lut_LC_9_25_3.C_ON=1'b0;
    defparam i15277_4_lut_LC_9_25_3.SEQ_MODE=4'b0000;
    defparam i15277_4_lut_LC_9_25_3.LUT_INIT=16'b0000000000101111;
    LogicCell40 i15277_4_lut_LC_9_25_3 (
            .in0(N__37363),
            .in1(N__33770),
            .in2(N__33863),
            .in3(N__33859),
            .lcout(n17356),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i2_LC_9_25_4 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i2_LC_9_25_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i2_LC_9_25_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.tx.r_Clock_Count__i2_LC_9_25_4  (
            .in0(N__33803),
            .in1(N__40289),
            .in2(_gnd_net_),
            .in3(N__33793),
            .lcout(r_Clock_Count_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50359),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i83_LC_9_25_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i83_LC_9_25_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i83_LC_9_25_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i83_LC_9_25_5  (
            .in0(N__45117),
            .in1(N__33881),
            .in2(_gnd_net_),
            .in3(N__36516),
            .lcout(data_in_10_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50359),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i11216_2_lut_LC_9_25_6 .C_ON=1'b0;
    defparam \c0.tx.i11216_2_lut_LC_9_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i11216_2_lut_LC_9_25_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.tx.i11216_2_lut_LC_9_25_6  (
            .in0(_gnd_net_),
            .in1(N__40101),
            .in2(_gnd_net_),
            .in3(N__40288),
            .lcout(n13601),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i59_LC_9_25_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i59_LC_9_25_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i59_LC_9_25_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i59_LC_9_25_7  (
            .in0(N__45116),
            .in1(N__33931),
            .in2(_gnd_net_),
            .in3(N__33750),
            .lcout(data_in_7_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50359),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i7_LC_9_26_0 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i7_LC_9_26_0 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i7_LC_9_26_0 .LUT_INIT=16'b1100101011001100;
    LogicCell40 \c0.rx.r_Rx_Byte_i7_LC_9_26_0  (
            .in0(N__37917),
            .in1(N__37117),
            .in2(N__33911),
            .in3(N__33731),
            .lcout(rx_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50370),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i167_LC_9_26_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i167_LC_9_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i167_LC_9_26_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_0___i167_LC_9_26_1  (
            .in0(N__33953),
            .in1(N__33713),
            .in2(_gnd_net_),
            .in3(N__45141),
            .lcout(data_in_20_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50370),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_i1_LC_9_26_2 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_i1_LC_9_26_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Bit_Index_i1_LC_9_26_2 .LUT_INIT=16'b1100110000101000;
    LogicCell40 \c0.tx.r_Bit_Index_i1_LC_9_26_2  (
            .in0(N__37440),
            .in1(N__39122),
            .in2(N__38925),
            .in3(N__38950),
            .lcout(r_Bit_Index_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50370),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i131_LC_9_26_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i131_LC_9_26_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i131_LC_9_26_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_0___i131_LC_9_26_3  (
            .in0(N__38405),
            .in1(N__34045),
            .in2(_gnd_net_),
            .in3(N__45140),
            .lcout(data_in_16_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50370),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i3_LC_9_26_5 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i3_LC_9_26_5 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i3_LC_9_26_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.rx.r_Rx_Byte_i3_LC_9_26_5  (
            .in0(N__34034),
            .in1(N__33903),
            .in2(N__33997),
            .in3(N__37918),
            .lcout(rx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50370),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i5_LC_9_26_6 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i5_LC_9_26_6 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i5_LC_9_26_6 .LUT_INIT=16'b1100110011001010;
    LogicCell40 \c0.rx.r_Rx_Byte_i5_LC_9_26_6  (
            .in0(N__37916),
            .in1(N__37702),
            .in2(N__33910),
            .in3(N__33980),
            .lcout(rx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50370),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_8__7__3526_LC_9_27_0 .C_ON=1'b0;
    defparam \c0.data_out_8__7__3526_LC_9_27_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_8__7__3526_LC_9_27_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_8__7__3526_LC_9_27_0  (
            .in0(N__46049),
            .in1(N__34907),
            .in2(_gnd_net_),
            .in3(N__45899),
            .lcout(data_out_8_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50377),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i159_LC_9_27_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i159_LC_9_27_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i159_LC_9_27_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i159_LC_9_27_1  (
            .in0(N__33952),
            .in1(N__45105),
            .in2(_gnd_net_),
            .in3(N__37774),
            .lcout(data_in_19_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50377),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_8__6__3527_LC_9_27_2 .C_ON=1'b0;
    defparam \c0.data_out_8__6__3527_LC_9_27_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_8__6__3527_LC_9_27_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_8__6__3527_LC_9_27_2  (
            .in0(N__46048),
            .in1(N__34982),
            .in2(_gnd_net_),
            .in3(N__46134),
            .lcout(data_out_8_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50377),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i67_LC_9_27_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i67_LC_9_27_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i67_LC_9_27_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_0___i67_LC_9_27_3  (
            .in0(N__36497),
            .in1(N__33924),
            .in2(_gnd_net_),
            .in3(N__45110),
            .lcout(data_in_8_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50377),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i1_LC_9_27_5 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i1_LC_9_27_5 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i1_LC_9_27_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.rx.r_Rx_Byte_i1_LC_9_27_5  (
            .in0(N__37952),
            .in1(N__33902),
            .in2(N__37754),
            .in3(N__37919),
            .lcout(rx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50377),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i91_LC_9_27_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i91_LC_9_27_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i91_LC_9_27_6 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i91_LC_9_27_6  (
            .in0(N__34694),
            .in1(_gnd_net_),
            .in2(N__45252),
            .in3(N__33877),
            .lcout(data_in_11_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50377),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i99_LC_9_27_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i99_LC_9_27_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i99_LC_9_27_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i99_LC_9_27_7  (
            .in0(N__34709),
            .in1(N__45106),
            .in2(_gnd_net_),
            .in3(N__34693),
            .lcout(data_in_12_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50377),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15728_2_lut_LC_9_28_0 .C_ON=1'b0;
    defparam \c0.i15728_2_lut_LC_9_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.i15728_2_lut_LC_9_28_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i15728_2_lut_LC_9_28_0  (
            .in0(_gnd_net_),
            .in1(N__43650),
            .in2(_gnd_net_),
            .in3(N__48420),
            .lcout(\c0.n17911 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_next_state_i0_LC_9_28_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_next_state_i0_LC_9_28_1 .SEQ_MODE=4'b1000;
    defparam \c0.FRAME_MATCHER_next_state_i0_LC_9_28_1 .LUT_INIT=16'b1111011101110111;
    LogicCell40 \c0.FRAME_MATCHER_next_state_i0_LC_9_28_1  (
            .in0(N__34685),
            .in1(N__34457),
            .in2(N__34288),
            .in3(N__34325),
            .lcout(FRAME_MATCHER_next_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50386),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i5_3_lut_LC_9_28_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i5_3_lut_LC_9_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i5_3_lut_LC_9_28_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_0_i5_3_lut_LC_9_28_2  (
            .in0(N__41476),
            .in1(N__41825),
            .in2(_gnd_net_),
            .in3(N__48421),
            .lcout(\c0.n5_adj_2488 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i134_LC_9_28_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i134_LC_9_28_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i134_LC_9_28_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i134_LC_9_28_5  (
            .in0(N__45142),
            .in1(N__38725),
            .in2(_gnd_net_),
            .in3(N__34268),
            .lcout(data_in_16_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50386),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i15793_2_lut_3_lut_LC_9_28_7 .C_ON=1'b0;
    defparam \c0.rx.i15793_2_lut_3_lut_LC_9_28_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i15793_2_lut_3_lut_LC_9_28_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \c0.rx.i15793_2_lut_3_lut_LC_9_28_7  (
            .in0(N__37914),
            .in1(N__39571),
            .in2(_gnd_net_),
            .in3(N__34253),
            .lcout(\c0.rx.n18066 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2270__i0_LC_9_29_0.C_ON=1'b1;
    defparam rand_setpoint_2270__i0_LC_9_29_0.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2270__i0_LC_9_29_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2270__i0_LC_9_29_0 (
            .in0(_gnd_net_),
            .in1(N__34211),
            .in2(N__39436),
            .in3(_gnd_net_),
            .lcout(rand_setpoint_0),
            .ltout(),
            .carryin(bfn_9_29_0_),
            .carryout(n16412),
            .clk(N__50393),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2270__i1_LC_9_29_1.C_ON=1'b1;
    defparam rand_setpoint_2270__i1_LC_9_29_1.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2270__i1_LC_9_29_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2270__i1_LC_9_29_1 (
            .in0(_gnd_net_),
            .in1(N__34148),
            .in2(N__39160),
            .in3(N__34115),
            .lcout(rand_setpoint_1),
            .ltout(),
            .carryin(n16412),
            .carryout(n16413),
            .clk(N__50393),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2270__i2_LC_9_29_2.C_ON=1'b1;
    defparam rand_setpoint_2270__i2_LC_9_29_2.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2270__i2_LC_9_29_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2270__i2_LC_9_29_2 (
            .in0(_gnd_net_),
            .in1(N__34088),
            .in2(N__37738),
            .in3(N__34052),
            .lcout(rand_setpoint_2),
            .ltout(),
            .carryin(n16413),
            .carryout(n16414),
            .clk(N__50393),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2270__i3_LC_9_29_3.C_ON=1'b1;
    defparam rand_setpoint_2270__i3_LC_9_29_3.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2270__i3_LC_9_29_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2270__i3_LC_9_29_3 (
            .in0(_gnd_net_),
            .in1(N__35205),
            .in2(N__43351),
            .in3(N__35156),
            .lcout(rand_setpoint_3),
            .ltout(),
            .carryin(n16414),
            .carryout(n16415),
            .clk(N__50393),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2270__i4_LC_9_29_4.C_ON=1'b1;
    defparam rand_setpoint_2270__i4_LC_9_29_4.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2270__i4_LC_9_29_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2270__i4_LC_9_29_4 (
            .in0(_gnd_net_),
            .in1(N__35139),
            .in2(N__38216),
            .in3(N__35102),
            .lcout(rand_setpoint_4),
            .ltout(),
            .carryin(n16415),
            .carryout(n16416),
            .clk(N__50393),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2270__i5_LC_9_29_5.C_ON=1'b1;
    defparam rand_setpoint_2270__i5_LC_9_29_5.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2270__i5_LC_9_29_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2270__i5_LC_9_29_5 (
            .in0(_gnd_net_),
            .in1(N__35087),
            .in2(N__39412),
            .in3(N__35045),
            .lcout(rand_setpoint_5),
            .ltout(),
            .carryin(n16416),
            .carryout(n16417),
            .clk(N__50393),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2270__i6_LC_9_29_6.C_ON=1'b1;
    defparam rand_setpoint_2270__i6_LC_9_29_6.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2270__i6_LC_9_29_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2270__i6_LC_9_29_6 (
            .in0(_gnd_net_),
            .in1(N__34978),
            .in2(N__35039),
            .in3(N__34967),
            .lcout(rand_setpoint_6),
            .ltout(),
            .carryin(n16417),
            .carryout(n16418),
            .clk(N__50393),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2270__i7_LC_9_29_7.C_ON=1'b1;
    defparam rand_setpoint_2270__i7_LC_9_29_7.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2270__i7_LC_9_29_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2270__i7_LC_9_29_7 (
            .in0(_gnd_net_),
            .in1(N__34951),
            .in2(N__34906),
            .in3(N__34889),
            .lcout(rand_setpoint_7),
            .ltout(),
            .carryin(n16418),
            .carryout(n16419),
            .clk(N__50393),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2270__i8_LC_9_30_0.C_ON=1'b1;
    defparam rand_setpoint_2270__i8_LC_9_30_0.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2270__i8_LC_9_30_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2270__i8_LC_9_30_0 (
            .in0(_gnd_net_),
            .in1(N__34867),
            .in2(N__41500),
            .in3(N__34832),
            .lcout(rand_setpoint_8),
            .ltout(),
            .carryin(bfn_9_30_0_),
            .carryout(n16420),
            .clk(N__50398),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2270__i9_LC_9_30_1.C_ON=1'b1;
    defparam rand_setpoint_2270__i9_LC_9_30_1.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2270__i9_LC_9_30_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2270__i9_LC_9_30_1 (
            .in0(_gnd_net_),
            .in1(N__34813),
            .in2(N__44209),
            .in3(N__34772),
            .lcout(rand_setpoint_9),
            .ltout(),
            .carryin(n16420),
            .carryout(n16421),
            .clk(N__50398),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2270__i10_LC_9_30_2.C_ON=1'b1;
    defparam rand_setpoint_2270__i10_LC_9_30_2.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2270__i10_LC_9_30_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2270__i10_LC_9_30_2 (
            .in0(_gnd_net_),
            .in1(N__34745),
            .in2(N__38126),
            .in3(N__34712),
            .lcout(rand_setpoint_10),
            .ltout(),
            .carryin(n16421),
            .carryout(n16422),
            .clk(N__50398),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2270__i11_LC_9_30_3.C_ON=1'b1;
    defparam rand_setpoint_2270__i11_LC_9_30_3.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2270__i11_LC_9_30_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2270__i11_LC_9_30_3 (
            .in0(_gnd_net_),
            .in1(N__35689),
            .in2(N__38192),
            .in3(N__35666),
            .lcout(rand_setpoint_11),
            .ltout(),
            .carryin(n16422),
            .carryout(n16423),
            .clk(N__50398),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2270__i12_LC_9_30_4.C_ON=1'b1;
    defparam rand_setpoint_2270__i12_LC_9_30_4.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2270__i12_LC_9_30_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2270__i12_LC_9_30_4 (
            .in0(_gnd_net_),
            .in1(N__35657),
            .in2(N__41716),
            .in3(N__35606),
            .lcout(rand_setpoint_12),
            .ltout(),
            .carryin(n16423),
            .carryout(n16424),
            .clk(N__50398),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2270__i13_LC_9_30_5.C_ON=1'b1;
    defparam rand_setpoint_2270__i13_LC_9_30_5.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2270__i13_LC_9_30_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2270__i13_LC_9_30_5 (
            .in0(_gnd_net_),
            .in1(N__35585),
            .in2(N__41410),
            .in3(N__35537),
            .lcout(rand_setpoint_13),
            .ltout(),
            .carryin(n16424),
            .carryout(n16425),
            .clk(N__50398),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2270__i14_LC_9_30_6.C_ON=1'b1;
    defparam rand_setpoint_2270__i14_LC_9_30_6.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2270__i14_LC_9_30_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2270__i14_LC_9_30_6 (
            .in0(_gnd_net_),
            .in1(N__40561),
            .in2(N__35522),
            .in3(N__35477),
            .lcout(rand_setpoint_14),
            .ltout(),
            .carryin(n16425),
            .carryout(n16426),
            .clk(N__50398),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2270__i15_LC_9_30_7.C_ON=1'b1;
    defparam rand_setpoint_2270__i15_LC_9_30_7.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2270__i15_LC_9_30_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2270__i15_LC_9_30_7 (
            .in0(_gnd_net_),
            .in1(N__35458),
            .in2(N__40588),
            .in3(N__35411),
            .lcout(rand_setpoint_15),
            .ltout(),
            .carryin(n16426),
            .carryout(n16427),
            .clk(N__50398),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2270__i16_LC_9_31_0.C_ON=1'b1;
    defparam rand_setpoint_2270__i16_LC_9_31_0.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2270__i16_LC_9_31_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2270__i16_LC_9_31_0 (
            .in0(_gnd_net_),
            .in1(N__35396),
            .in2(N__41845),
            .in3(N__35360),
            .lcout(rand_setpoint_16),
            .ltout(),
            .carryin(bfn_9_31_0_),
            .carryout(n16428),
            .clk(N__50404),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2270__i17_LC_9_31_1.C_ON=1'b1;
    defparam rand_setpoint_2270__i17_LC_9_31_1.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2270__i17_LC_9_31_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2270__i17_LC_9_31_1 (
            .in0(_gnd_net_),
            .in1(N__35345),
            .in2(N__43858),
            .in3(N__35309),
            .lcout(rand_setpoint_17),
            .ltout(),
            .carryin(n16428),
            .carryout(n16429),
            .clk(N__50404),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2270__i18_LC_9_31_2.C_ON=1'b1;
    defparam rand_setpoint_2270__i18_LC_9_31_2.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2270__i18_LC_9_31_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2270__i18_LC_9_31_2 (
            .in0(_gnd_net_),
            .in1(N__35289),
            .in2(N__39505),
            .in3(N__35264),
            .lcout(rand_setpoint_18),
            .ltout(),
            .carryin(n16429),
            .carryout(n16430),
            .clk(N__50404),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2270__i19_LC_9_31_3.C_ON=1'b1;
    defparam rand_setpoint_2270__i19_LC_9_31_3.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2270__i19_LC_9_31_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2270__i19_LC_9_31_3 (
            .in0(_gnd_net_),
            .in1(N__35249),
            .in2(N__40765),
            .in3(N__35213),
            .lcout(rand_setpoint_19),
            .ltout(),
            .carryin(n16430),
            .carryout(n16431),
            .clk(N__50404),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2270__i20_LC_9_31_4.C_ON=1'b1;
    defparam rand_setpoint_2270__i20_LC_9_31_4.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2270__i20_LC_9_31_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2270__i20_LC_9_31_4 (
            .in0(_gnd_net_),
            .in1(N__36144),
            .in2(N__40615),
            .in3(N__36107),
            .lcout(rand_setpoint_20),
            .ltout(),
            .carryin(n16431),
            .carryout(n16432),
            .clk(N__50404),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2270__i21_LC_9_31_5.C_ON=1'b1;
    defparam rand_setpoint_2270__i21_LC_9_31_5.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2270__i21_LC_9_31_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2270__i21_LC_9_31_5 (
            .in0(_gnd_net_),
            .in1(N__43879),
            .in2(N__36098),
            .in3(N__36047),
            .lcout(rand_setpoint_21),
            .ltout(),
            .carryin(n16432),
            .carryout(n16433),
            .clk(N__50404),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2270__i22_LC_9_31_6.C_ON=1'b1;
    defparam rand_setpoint_2270__i22_LC_9_31_6.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2270__i22_LC_9_31_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2270__i22_LC_9_31_6 (
            .in0(_gnd_net_),
            .in1(N__38227),
            .in2(N__36034),
            .in3(N__36008),
            .lcout(rand_setpoint_22),
            .ltout(),
            .carryin(n16433),
            .carryout(n16434),
            .clk(N__50404),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2270__i23_LC_9_31_7.C_ON=1'b1;
    defparam rand_setpoint_2270__i23_LC_9_31_7.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2270__i23_LC_9_31_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2270__i23_LC_9_31_7 (
            .in0(_gnd_net_),
            .in1(N__35991),
            .in2(N__41881),
            .in3(N__35954),
            .lcout(rand_setpoint_23),
            .ltout(),
            .carryin(n16434),
            .carryout(n16435),
            .clk(N__50404),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2270__i24_LC_9_32_0.C_ON=1'b1;
    defparam rand_setpoint_2270__i24_LC_9_32_0.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2270__i24_LC_9_32_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2270__i24_LC_9_32_0 (
            .in0(_gnd_net_),
            .in1(N__35939),
            .in2(N__38249),
            .in3(N__35891),
            .lcout(rand_setpoint_24),
            .ltout(),
            .carryin(bfn_9_32_0_),
            .carryout(n16436),
            .clk(N__50410),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2270__i25_LC_9_32_1.C_ON=1'b1;
    defparam rand_setpoint_2270__i25_LC_9_32_1.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2270__i25_LC_9_32_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2270__i25_LC_9_32_1 (
            .in0(_gnd_net_),
            .in1(N__35867),
            .in2(N__38176),
            .in3(N__35831),
            .lcout(rand_setpoint_25),
            .ltout(),
            .carryin(n16436),
            .carryout(n16437),
            .clk(N__50410),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2270__i26_LC_9_32_2.C_ON=1'b1;
    defparam rand_setpoint_2270__i26_LC_9_32_2.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2270__i26_LC_9_32_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2270__i26_LC_9_32_2 (
            .in0(_gnd_net_),
            .in1(N__35802),
            .in2(N__39463),
            .in3(N__35777),
            .lcout(rand_setpoint_26),
            .ltout(),
            .carryin(n16437),
            .carryout(n16438),
            .clk(N__50410),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2270__i27_LC_9_32_3.C_ON=1'b1;
    defparam rand_setpoint_2270__i27_LC_9_32_3.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2270__i27_LC_9_32_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2270__i27_LC_9_32_3 (
            .in0(_gnd_net_),
            .in1(N__35759),
            .in2(N__38282),
            .in3(N__35720),
            .lcout(rand_setpoint_27),
            .ltout(),
            .carryin(n16438),
            .carryout(n16439),
            .clk(N__50410),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2270__i28_LC_9_32_4.C_ON=1'b1;
    defparam rand_setpoint_2270__i28_LC_9_32_4.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2270__i28_LC_9_32_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2270__i28_LC_9_32_4 (
            .in0(_gnd_net_),
            .in1(N__36458),
            .in2(N__41587),
            .in3(N__36413),
            .lcout(rand_setpoint_28),
            .ltout(),
            .carryin(n16439),
            .carryout(n16440),
            .clk(N__50410),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2270__i29_LC_9_32_5.C_ON=1'b1;
    defparam rand_setpoint_2270__i29_LC_9_32_5.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2270__i29_LC_9_32_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2270__i29_LC_9_32_5 (
            .in0(_gnd_net_),
            .in1(N__38264),
            .in2(N__36399),
            .in3(N__36359),
            .lcout(rand_setpoint_29),
            .ltout(),
            .carryin(n16440),
            .carryout(n16441),
            .clk(N__50410),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2270__i30_LC_9_32_6.C_ON=1'b1;
    defparam rand_setpoint_2270__i30_LC_9_32_6.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2270__i30_LC_9_32_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2270__i30_LC_9_32_6 (
            .in0(_gnd_net_),
            .in1(N__38155),
            .in2(N__36353),
            .in3(N__36311),
            .lcout(rand_setpoint_30),
            .ltout(),
            .carryin(n16441),
            .carryout(n16442),
            .clk(N__50410),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2270__i31_LC_9_32_7.C_ON=1'b0;
    defparam rand_setpoint_2270__i31_LC_9_32_7.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2270__i31_LC_9_32_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 rand_setpoint_2270__i31_LC_9_32_7 (
            .in0(N__36297),
            .in1(N__38140),
            .in2(_gnd_net_),
            .in3(N__36263),
            .lcout(rand_setpoint_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50410),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i6_LC_10_19_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i6_LC_10_19_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i6_LC_10_19_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i6_LC_10_19_1  (
            .in0(N__45340),
            .in1(N__37604),
            .in2(_gnd_net_),
            .in3(N__36260),
            .lcout(data_in_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50305),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i7_LC_10_20_0 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i7_LC_10_20_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i7_LC_10_20_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.tx.r_Tx_Data_i7_LC_10_20_0  (
            .in0(N__37417),
            .in1(N__48683),
            .in2(_gnd_net_),
            .in3(N__38690),
            .lcout(r_Tx_Data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50313),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i54_LC_10_20_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i54_LC_10_20_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i54_LC_10_20_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_0___i54_LC_10_20_2  (
            .in0(N__36177),
            .in1(N__36224),
            .in2(_gnd_net_),
            .in3(N__45202),
            .lcout(data_in_6_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50313),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i124_LC_10_20_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i124_LC_10_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i124_LC_10_20_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i124_LC_10_20_5  (
            .in0(N__45200),
            .in1(N__37106),
            .in2(_gnd_net_),
            .in3(N__37087),
            .lcout(data_in_15_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50313),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i50_LC_10_20_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i50_LC_10_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i50_LC_10_20_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_0___i50_LC_10_20_6  (
            .in0(N__37015),
            .in1(N__39918),
            .in2(_gnd_net_),
            .in3(N__45201),
            .lcout(\c0.data_in_6_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50313),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i58_LC_10_21_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i58_LC_10_21_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i58_LC_10_21_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i58_LC_10_21_0  (
            .in0(N__37043),
            .in1(N__45198),
            .in2(_gnd_net_),
            .in3(N__37008),
            .lcout(\c0.data_in_7_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50320),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i84_LC_10_21_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i84_LC_10_21_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i84_LC_10_21_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_0___i84_LC_10_21_2  (
            .in0(N__36982),
            .in1(N__38570),
            .in2(_gnd_net_),
            .in3(N__45199),
            .lcout(data_in_10_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50320),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i48_LC_10_21_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i48_LC_10_21_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i48_LC_10_21_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i48_LC_10_21_5  (
            .in0(N__45197),
            .in1(N__36947),
            .in2(_gnd_net_),
            .in3(N__36902),
            .lcout(data_in_5_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50320),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_844_LC_10_21_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_844_LC_10_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_844_LC_10_21_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_844_LC_10_21_6  (
            .in0(_gnd_net_),
            .in1(N__36858),
            .in2(_gnd_net_),
            .in3(N__36832),
            .lcout(\c0.n6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i89_LC_10_22_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i89_LC_10_22_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i89_LC_10_22_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i89_LC_10_22_1  (
            .in0(N__38843),
            .in1(N__45208),
            .in2(_gnd_net_),
            .in3(N__36778),
            .lcout(data_in_11_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50331),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i4723_2_lut_LC_10_22_2 .C_ON=1'b0;
    defparam \c0.tx.i4723_2_lut_LC_10_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i4723_2_lut_LC_10_22_2 .LUT_INIT=16'b1110111011101110;
    LogicCell40 \c0.tx.i4723_2_lut_LC_10_22_2  (
            .in0(N__40214),
            .in1(N__40160),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n7086),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i122_LC_10_22_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i122_LC_10_22_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i122_LC_10_22_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i122_LC_10_22_3  (
            .in0(N__36754),
            .in1(N__45206),
            .in2(_gnd_net_),
            .in3(N__38972),
            .lcout(data_in_15_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50331),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_976_LC_10_22_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_976_LC_10_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_976_LC_10_22_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_976_LC_10_22_4  (
            .in0(N__36729),
            .in1(N__36690),
            .in2(N__36624),
            .in3(N__36580),
            .lcout(\c0.n8989 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i75_LC_10_22_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i75_LC_10_22_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i75_LC_10_22_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i75_LC_10_22_6  (
            .in0(N__45205),
            .in1(N__36492),
            .in2(_gnd_net_),
            .in3(N__36523),
            .lcout(data_in_9_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50331),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i152_LC_10_22_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i152_LC_10_22_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i152_LC_10_22_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i152_LC_10_22_7  (
            .in0(N__37132),
            .in1(N__45207),
            .in2(_gnd_net_),
            .in3(N__37067),
            .lcout(data_in_18_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50331),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i168_LC_10_23_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i168_LC_10_23_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i168_LC_10_23_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i168_LC_10_23_0  (
            .in0(N__44948),
            .in1(N__37121),
            .in2(_gnd_net_),
            .in3(N__37075),
            .lcout(data_in_20_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50340),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i132_LC_10_23_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i132_LC_10_23_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i132_LC_10_23_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i132_LC_10_23_1  (
            .in0(N__45164),
            .in1(N__37102),
            .in2(_gnd_net_),
            .in3(N__38672),
            .lcout(data_in_16_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50340),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_3__7__3566_LC_10_23_2 .C_ON=1'b0;
    defparam \c0.data_out_3__7__3566_LC_10_23_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_3__7__3566_LC_10_23_2 .LUT_INIT=16'b1010110010101010;
    LogicCell40 \c0.data_out_3__7__3566_LC_10_23_2  (
            .in0(N__46412),
            .in1(N__46880),
            .in2(N__47143),
            .in3(N__47297),
            .lcout(data_out_5__7__N_931),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50340),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i116_LC_10_23_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i116_LC_10_23_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i116_LC_10_23_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i116_LC_10_23_4  (
            .in0(N__44947),
            .in1(N__38713),
            .in2(_gnd_net_),
            .in3(N__37091),
            .lcout(data_in_14_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50340),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i160_LC_10_23_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i160_LC_10_23_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i160_LC_10_23_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i160_LC_10_23_5  (
            .in0(N__37076),
            .in1(N__44949),
            .in2(_gnd_net_),
            .in3(N__37066),
            .lcout(data_in_19_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50340),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_i2_LC_10_23_6 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_i2_LC_10_23_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Bit_Index_i2_LC_10_23_6 .LUT_INIT=16'b1111100000001000;
    LogicCell40 \c0.tx.r_Bit_Index_i2_LC_10_23_6  (
            .in0(N__37396),
            .in1(N__37286),
            .in2(N__38927),
            .in3(N__37055),
            .lcout(r_Bit_Index_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50340),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_i0_LC_10_23_7 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_i0_LC_10_23_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_SM_Main_i0_LC_10_23_7 .LUT_INIT=16'b0000001100001010;
    LogicCell40 \c0.tx.r_SM_Main_i0_LC_10_23_7  (
            .in0(N__37049),
            .in1(N__40404),
            .in2(N__40376),
            .in3(N__40221),
            .lcout(r_SM_Main_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50340),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i2_LC_10_24_0 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i2_LC_10_24_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i2_LC_10_24_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.tx.r_Tx_Data_i2_LC_10_24_0  (
            .in0(N__37274),
            .in1(N__48674),
            .in2(_gnd_net_),
            .in3(N__38639),
            .lcout(r_Tx_Data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50350),
            .ce(),
            .sr(_gnd_net_));
    defparam i15317_2_lut_LC_10_24_1.C_ON=1'b0;
    defparam i15317_2_lut_LC_10_24_1.SEQ_MODE=4'b0000;
    defparam i15317_2_lut_LC_10_24_1.LUT_INIT=16'b1111111111001100;
    LogicCell40 i15317_2_lut_LC_10_24_1 (
            .in0(_gnd_net_),
            .in1(N__37441),
            .in2(_gnd_net_),
            .in3(N__38943),
            .lcout(n17767),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i2_3_lut_LC_10_24_2 .C_ON=1'b0;
    defparam \c0.tx.i2_3_lut_LC_10_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i2_3_lut_LC_10_24_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.tx.i2_3_lut_LC_10_24_2  (
            .in0(N__39125),
            .in1(N__37402),
            .in2(_gnd_net_),
            .in3(N__38918),
            .lcout(\c0.tx.n17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_Bit_Index_2__bdd_4_lut_LC_10_24_3.C_ON=1'b0;
    defparam r_Bit_Index_2__bdd_4_lut_LC_10_24_3.SEQ_MODE=4'b0000;
    defparam r_Bit_Index_2__bdd_4_lut_LC_10_24_3.LUT_INIT=16'b1010110011110000;
    LogicCell40 r_Bit_Index_2__bdd_4_lut_LC_10_24_3 (
            .in0(N__48614),
            .in1(N__37273),
            .in2(N__37403),
            .in3(N__39124),
            .lcout(n18462),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_2_lut_4_lut_LC_10_24_4 .C_ON=1'b0;
    defparam \c0.tx.i1_2_lut_4_lut_LC_10_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_2_lut_4_lut_LC_10_24_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \c0.tx.i1_2_lut_4_lut_LC_10_24_4  (
            .in0(N__37252),
            .in1(N__37320),
            .in2(N__40222),
            .in3(N__37209),
            .lcout(n12_adj_2618),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i11594214_i1_3_lut_LC_10_24_5.C_ON=1'b0;
    defparam i11594214_i1_3_lut_LC_10_24_5.SEQ_MODE=4'b0000;
    defparam i11594214_i1_3_lut_LC_10_24_5.LUT_INIT=16'b1010111110100000;
    LogicCell40 i11594214_i1_3_lut_LC_10_24_5 (
            .in0(N__39077),
            .in1(_gnd_net_),
            .in2(N__38926),
            .in3(N__38807),
            .lcout(),
            .ltout(n1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_2__I_0_56_i3_3_lut_LC_10_24_6 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_2__I_0_56_i3_3_lut_LC_10_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.r_SM_Main_2__I_0_56_i3_3_lut_LC_10_24_6 .LUT_INIT=16'b1111101001010101;
    LogicCell40 \c0.tx.r_SM_Main_2__I_0_56_i3_3_lut_LC_10_24_6  (
            .in0(N__40206),
            .in1(_gnd_net_),
            .in2(N__37181),
            .in3(N__40146),
            .lcout(),
            .ltout(n3_adj_2650_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.o_Tx_Serial_45_LC_10_24_7 .C_ON=1'b0;
    defparam \c0.tx.o_Tx_Serial_45_LC_10_24_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.o_Tx_Serial_45_LC_10_24_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \c0.tx.o_Tx_Serial_45_LC_10_24_7  (
            .in0(_gnd_net_),
            .in1(N__37144),
            .in2(N__37178),
            .in3(N__40346),
            .lcout(tx_o_adj_2584),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50350),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_831_LC_10_25_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_831_LC_10_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_831_LC_10_25_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_831_LC_10_25_0  (
            .in0(_gnd_net_),
            .in1(N__46148),
            .in2(_gnd_net_),
            .in3(N__41480),
            .lcout(\c0.n9087 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_881_LC_10_25_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_881_LC_10_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_881_LC_10_25_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_881_LC_10_25_2  (
            .in0(N__44489),
            .in1(N__43274),
            .in2(_gnd_net_),
            .in3(N__43332),
            .lcout(\c0.n17556 ),
            .ltout(\c0.n17556_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_9__3__3522_LC_10_25_3 .C_ON=1'b0;
    defparam \c0.data_out_9__3__3522_LC_10_25_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_9__3__3522_LC_10_25_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_9__3__3522_LC_10_25_3  (
            .in0(N__46149),
            .in1(N__37784),
            .in2(N__37664),
            .in3(N__43532),
            .lcout(\c0.data_out_9_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50360),
            .ce(N__46034),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1012_LC_10_25_4 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1012_LC_10_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1012_LC_10_25_4 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \c0.i6_4_lut_adj_1012_LC_10_25_4  (
            .in0(N__37656),
            .in1(N__37608),
            .in2(N__37574),
            .in3(N__37519),
            .lcout(\c0.n16_adj_2513 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i137_LC_10_26_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i137_LC_10_26_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i137_LC_10_26_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i137_LC_10_26_0  (
            .in0(N__37457),
            .in1(N__45111),
            .in2(_gnd_net_),
            .in3(N__39019),
            .lcout(data_in_17_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50371),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i7381_2_lut_4_lut_LC_10_26_1 .C_ON=1'b0;
    defparam \c0.tx.i7381_2_lut_4_lut_LC_10_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i7381_2_lut_4_lut_LC_10_26_1 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \c0.tx.i7381_2_lut_4_lut_LC_10_26_1  (
            .in0(N__37398),
            .in1(N__38906),
            .in2(N__40133),
            .in3(N__39107),
            .lcout(n9796),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_Bit_Index_2__bdd_4_lut_15992_LC_10_26_2.C_ON=1'b0;
    defparam r_Bit_Index_2__bdd_4_lut_15992_LC_10_26_2.SEQ_MODE=4'b0000;
    defparam r_Bit_Index_2__bdd_4_lut_15992_LC_10_26_2.LUT_INIT=16'b1011110010001100;
    LogicCell40 r_Bit_Index_2__bdd_4_lut_15992_LC_10_26_2 (
            .in0(N__37418),
            .in1(N__37397),
            .in2(N__39123),
            .in3(N__39052),
            .lcout(n18438),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_LC_10_26_3.C_ON=1'b0;
    defparam i1_3_lut_LC_10_26_3.SEQ_MODE=4'b0000;
    defparam i1_3_lut_LC_10_26_3.LUT_INIT=16'b0111011100000000;
    LogicCell40 i1_3_lut_LC_10_26_3 (
            .in0(N__40103),
            .in1(N__40290),
            .in2(_gnd_net_),
            .in3(N__37364),
            .lcout(n22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i8_LC_10_26_4 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i8_LC_10_26_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i8_LC_10_26_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.tx.r_Clock_Count__i8_LC_10_26_4  (
            .in0(N__40291),
            .in1(N__37334),
            .in2(_gnd_net_),
            .in3(N__37319),
            .lcout(r_Clock_Count_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50371),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_i1_LC_10_26_5 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_i1_LC_10_26_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_SM_Main_i1_LC_10_26_5 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \c0.tx.r_SM_Main_i1_LC_10_26_5  (
            .in0(N__40107),
            .in1(N__40414),
            .in2(N__40240),
            .in3(N__40292),
            .lcout(r_SM_Main_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50371),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_2_i5_3_lut_LC_10_26_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_2_i5_3_lut_LC_10_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_2_i5_3_lut_LC_10_26_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_2_i5_3_lut_LC_10_26_6  (
            .in0(N__46366),
            .in1(N__39485),
            .in2(_gnd_net_),
            .in3(N__48314),
            .lcout(\c0.n5_adj_2499 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_i2_LC_10_26_7 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_i2_LC_10_26_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_SM_Main_i2_LC_10_26_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \c0.tx.r_SM_Main_i2_LC_10_26_7  (
            .in0(N__40108),
            .in1(N__40415),
            .in2(N__40241),
            .in3(N__40293),
            .lcout(r_SM_Main_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50371),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1072_LC_10_27_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1072_LC_10_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1072_LC_10_27_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1072_LC_10_27_0  (
            .in0(N__40793),
            .in1(N__49706),
            .in2(_gnd_net_),
            .in3(N__43649),
            .lcout(\c0.n6_adj_2448 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i143_LC_10_27_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i143_LC_10_27_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i143_LC_10_27_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i143_LC_10_27_2  (
            .in0(N__37763),
            .in1(N__44792),
            .in2(_gnd_net_),
            .in3(N__37804),
            .lcout(data_in_17_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50378),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i151_LC_10_27_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i151_LC_10_27_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i151_LC_10_27_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i151_LC_10_27_3  (
            .in0(N__44791),
            .in1(N__37762),
            .in2(_gnd_net_),
            .in3(N__37775),
            .lcout(data_in_18_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50378),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i162_LC_10_27_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i162_LC_10_27_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i162_LC_10_27_5 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i162_LC_10_27_5  (
            .in0(N__37753),
            .in1(_gnd_net_),
            .in2(N__44968),
            .in3(N__39041),
            .lcout(data_in_20_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50378),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_8__2__3531_LC_10_27_7 .C_ON=1'b0;
    defparam \c0.data_out_8__2__3531_LC_10_27_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_8__2__3531_LC_10_27_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_8__2__3531_LC_10_27_7  (
            .in0(N__46041),
            .in1(N__37739),
            .in2(_gnd_net_),
            .in3(N__43328),
            .lcout(data_out_8_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50378),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i158_LC_10_28_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i158_LC_10_28_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i158_LC_10_28_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i158_LC_10_28_0  (
            .in0(N__37691),
            .in1(N__44866),
            .in2(_gnd_net_),
            .in3(N__37717),
            .lcout(data_in_19_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50387),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i166_LC_10_28_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i166_LC_10_28_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i166_LC_10_28_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i166_LC_10_28_1  (
            .in0(N__44865),
            .in1(N__37706),
            .in2(_gnd_net_),
            .in3(N__37690),
            .lcout(data_in_20_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50387),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_LC_10_28_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_LC_10_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_LC_10_28_2 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter_1__bdd_4_lut_LC_10_28_2  (
            .in0(N__37682),
            .in1(N__48110),
            .in2(N__37673),
            .in3(N__47984),
            .lcout(\c0.n18498 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i2_3_lut_LC_10_28_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i2_3_lut_LC_10_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i2_3_lut_LC_10_28_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_0_i2_3_lut_LC_10_28_3  (
            .in0(N__40701),
            .in1(N__44141),
            .in2(_gnd_net_),
            .in3(N__48425),
            .lcout(),
            .ltout(\c0.n2_adj_2487_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18498_bdd_4_lut_LC_10_28_4 .C_ON=1'b0;
    defparam \c0.n18498_bdd_4_lut_LC_10_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.n18498_bdd_4_lut_LC_10_28_4 .LUT_INIT=16'b1100110011100010;
    LogicCell40 \c0.n18498_bdd_4_lut_LC_10_28_4  (
            .in0(N__41336),
            .in1(N__37961),
            .in2(N__37955),
            .in3(N__48111),
            .lcout(\c0.n18501 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.equal_104_i4_2_lut_LC_10_28_5 .C_ON=1'b0;
    defparam \c0.rx.equal_104_i4_2_lut_LC_10_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.equal_104_i4_2_lut_LC_10_28_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.rx.equal_104_i4_2_lut_LC_10_28_5  (
            .in0(_gnd_net_),
            .in1(N__39230),
            .in2(_gnd_net_),
            .in3(N__39286),
            .lcout(n4_adj_2649),
            .ltout(n4_adj_2649_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i0_LC_10_28_6 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i0_LC_10_28_6 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i0_LC_10_28_6 .LUT_INIT=16'b1010101110101000;
    LogicCell40 \c0.rx.r_Rx_Byte_i0_LC_10_28_6  (
            .in0(N__37834),
            .in1(N__37945),
            .in2(N__37922),
            .in3(N__37915),
            .lcout(rx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50387),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__0__3597_LC_10_29_0 .C_ON=1'b0;
    defparam \c0.data_out_0__0__3597_LC_10_29_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__0__3597_LC_10_29_0 .LUT_INIT=16'b1010101011100010;
    LogicCell40 \c0.data_out_0__0__3597_LC_10_29_0  (
            .in0(N__47561),
            .in1(N__47400),
            .in2(N__46879),
            .in3(N__47079),
            .lcout(data_out_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50394),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i161_LC_10_29_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i161_LC_10_29_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i161_LC_10_29_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i161_LC_10_29_1  (
            .in0(N__37838),
            .in1(N__44890),
            .in2(_gnd_net_),
            .in3(N__37819),
            .lcout(data_in_20_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50394),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i135_LC_10_29_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i135_LC_10_29_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i135_LC_10_29_2 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i135_LC_10_29_2  (
            .in0(N__37808),
            .in1(_gnd_net_),
            .in2(N__45112),
            .in3(N__37792),
            .lcout(data_in_16_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50394),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i127_LC_10_29_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i127_LC_10_29_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i127_LC_10_29_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i127_LC_10_29_4  (
            .in0(N__44888),
            .in1(N__38200),
            .in2(_gnd_net_),
            .in3(N__37793),
            .lcout(data_in_15_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50394),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__3__3594_LC_10_29_5 .C_ON=1'b0;
    defparam \c0.data_out_0__3__3594_LC_10_29_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__3__3594_LC_10_29_5 .LUT_INIT=16'b1100010011001110;
    LogicCell40 \c0.data_out_0__3__3594_LC_10_29_5  (
            .in0(N__47399),
            .in1(N__47670),
            .in2(N__47111),
            .in3(N__46793),
            .lcout(data_out_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50394),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_8__4__3529_LC_10_29_6 .C_ON=1'b0;
    defparam \c0.data_out_8__4__3529_LC_10_29_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_8__4__3529_LC_10_29_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_8__4__3529_LC_10_29_6  (
            .in0(N__46033),
            .in1(N__38215),
            .in2(_gnd_net_),
            .in3(N__49603),
            .lcout(data_out_8_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50394),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i119_LC_10_29_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i119_LC_10_29_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i119_LC_10_29_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i119_LC_10_29_7  (
            .in0(N__38201),
            .in1(N__44889),
            .in2(_gnd_net_),
            .in3(N__44551),
            .lcout(data_in_14_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50394),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__3__3538_LC_10_30_0 .C_ON=1'b0;
    defparam \c0.data_out_7__3__3538_LC_10_30_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__3__3538_LC_10_30_0 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \c0.data_out_7__3__3538_LC_10_30_0  (
            .in0(N__47448),
            .in1(N__45677),
            .in2(N__46917),
            .in3(N__38191),
            .lcout(\c0.data_out_7_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50399),
            .ce(N__44192),
            .sr(_gnd_net_));
    defparam \c0.i15710_2_lut_LC_10_30_1 .C_ON=1'b0;
    defparam \c0.i15710_2_lut_LC_10_30_1 .SEQ_MODE=4'b0000;
    defparam \c0.i15710_2_lut_LC_10_30_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i15710_2_lut_LC_10_30_1  (
            .in0(N__38177),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47445),
            .lcout(\c0.n17962 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15722_2_lut_LC_10_30_2 .C_ON=1'b0;
    defparam \c0.i15722_2_lut_LC_10_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.i15722_2_lut_LC_10_30_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i15722_2_lut_LC_10_30_2  (
            .in0(N__47447),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38159),
            .lcout(\c0.n17972 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15723_2_lut_LC_10_30_3 .C_ON=1'b0;
    defparam \c0.i15723_2_lut_LC_10_30_3 .SEQ_MODE=4'b0000;
    defparam \c0.i15723_2_lut_LC_10_30_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i15723_2_lut_LC_10_30_3  (
            .in0(_gnd_net_),
            .in1(N__38141),
            .in2(_gnd_net_),
            .in3(N__47446),
            .lcout(\c0.n17974 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15760_2_lut_LC_10_30_4 .C_ON=1'b0;
    defparam \c0.i15760_2_lut_LC_10_30_4 .SEQ_MODE=4'b0000;
    defparam \c0.i15760_2_lut_LC_10_30_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i15760_2_lut_LC_10_30_4  (
            .in0(N__47444),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38125),
            .lcout(\c0.n17921 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i130_3_lut_4_lut_LC_10_30_5 .C_ON=1'b0;
    defparam \c0.rx.i130_3_lut_4_lut_LC_10_30_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i130_3_lut_4_lut_LC_10_30_5 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \c0.rx.i130_3_lut_4_lut_LC_10_30_5  (
            .in0(N__38111),
            .in1(N__38060),
            .in2(N__38021),
            .in3(N__38000),
            .lcout(\c0.rx.r_SM_Main_2_N_2380_2 ),
            .ltout(\c0.rx.r_SM_Main_2_N_2380_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i15739_2_lut_3_lut_4_lut_LC_10_30_6 .C_ON=1'b0;
    defparam \c0.rx.i15739_2_lut_3_lut_4_lut_LC_10_30_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i15739_2_lut_3_lut_4_lut_LC_10_30_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.rx.i15739_2_lut_3_lut_4_lut_LC_10_30_6  (
            .in0(N__40452),
            .in1(N__39236),
            .in2(N__37964),
            .in3(N__39300),
            .lcout(),
            .ltout(\c0.rx.n18000_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_0__bdd_4_lut_4_lut_LC_10_30_7 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_0__bdd_4_lut_4_lut_LC_10_30_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_SM_Main_0__bdd_4_lut_4_lut_LC_10_30_7 .LUT_INIT=16'b0111011111000000;
    LogicCell40 \c0.rx.r_SM_Main_0__bdd_4_lut_4_lut_LC_10_30_7  (
            .in0(N__39631),
            .in1(N__39711),
            .in2(N__38300),
            .in3(N__39590),
            .lcout(\c0.rx.n18594 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15874_4_lut_4_lut_4_lut_LC_10_31_0 .C_ON=1'b0;
    defparam \c0.i15874_4_lut_4_lut_4_lut_LC_10_31_0 .SEQ_MODE=4'b0000;
    defparam \c0.i15874_4_lut_4_lut_4_lut_LC_10_31_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \c0.i15874_4_lut_4_lut_4_lut_LC_10_31_0  (
            .in0(_gnd_net_),
            .in1(N__47106),
            .in2(_gnd_net_),
            .in3(N__47439),
            .lcout(n9519),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15714_2_lut_LC_10_31_1 .C_ON=1'b0;
    defparam \c0.i15714_2_lut_LC_10_31_1 .SEQ_MODE=4'b0000;
    defparam \c0.i15714_2_lut_LC_10_31_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i15714_2_lut_LC_10_31_1  (
            .in0(N__47441),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38281),
            .lcout(),
            .ltout(\c0.n17966_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_5__3__3554_LC_10_31_2 .C_ON=1'b0;
    defparam \c0.data_out_5__3__3554_LC_10_31_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_5__3__3554_LC_10_31_2 .LUT_INIT=16'b1111000011101110;
    LogicCell40 \c0.data_out_5__3__3554_LC_10_31_2  (
            .in0(N__40792),
            .in1(N__49443),
            .in2(N__38267),
            .in3(N__46891),
            .lcout(\c0.data_out_5_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50405),
            .ce(N__46516),
            .sr(_gnd_net_));
    defparam \c0.i15717_2_lut_LC_10_31_3 .C_ON=1'b0;
    defparam \c0.i15717_2_lut_LC_10_31_3 .SEQ_MODE=4'b0000;
    defparam \c0.i15717_2_lut_LC_10_31_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i15717_2_lut_LC_10_31_3  (
            .in0(N__47442),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38263),
            .lcout(),
            .ltout(\c0.n17970_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_5__5__3552_LC_10_31_4 .C_ON=1'b0;
    defparam \c0.data_out_5__5__3552_LC_10_31_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_5__5__3552_LC_10_31_4 .LUT_INIT=16'b1111010111100100;
    LogicCell40 \c0.data_out_5__5__3552_LC_10_31_4  (
            .in0(N__46892),
            .in1(N__49444),
            .in2(N__38252),
            .in3(N__49853),
            .lcout(\c0.data_out_7__5__N_543 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50405),
            .ce(N__46516),
            .sr(_gnd_net_));
    defparam \c0.i15705_2_lut_LC_10_31_5 .C_ON=1'b0;
    defparam \c0.i15705_2_lut_LC_10_31_5 .SEQ_MODE=4'b0000;
    defparam \c0.i15705_2_lut_LC_10_31_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i15705_2_lut_LC_10_31_5  (
            .in0(N__47440),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__38248),
            .lcout(),
            .ltout(\c0.n17957_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_5__0__3557_LC_10_31_6 .C_ON=1'b0;
    defparam \c0.data_out_5__0__3557_LC_10_31_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_5__0__3557_LC_10_31_6 .LUT_INIT=16'b1111000011011101;
    LogicCell40 \c0.data_out_5__0__3557_LC_10_31_6  (
            .in0(N__47771),
            .in1(N__49442),
            .in2(N__38234),
            .in3(N__46890),
            .lcout(\c0.data_out_6__3__N_788 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50405),
            .ce(N__46516),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__6__3543_LC_10_31_7 .C_ON=1'b0;
    defparam \c0.data_out_6__6__3543_LC_10_31_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__6__3543_LC_10_31_7 .LUT_INIT=16'b1010000000110011;
    LogicCell40 \c0.data_out_6__6__3543_LC_10_31_7  (
            .in0(N__47443),
            .in1(N__40631),
            .in2(N__38231),
            .in3(N__46893),
            .lcout(\c0.data_out_6_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50405),
            .ce(N__46516),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i147_LC_10_32_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i147_LC_10_32_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i147_LC_10_32_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i147_LC_10_32_2  (
            .in0(N__44649),
            .in1(N__38413),
            .in2(_gnd_net_),
            .in3(N__38474),
            .lcout(data_in_18_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50411),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i149_LC_10_32_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i149_LC_10_32_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i149_LC_10_32_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i149_LC_10_32_4  (
            .in0(N__38432),
            .in1(N__44652),
            .in2(_gnd_net_),
            .in3(N__38422),
            .lcout(data_in_18_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50411),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i157_LC_10_32_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i157_LC_10_32_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i157_LC_10_32_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i157_LC_10_32_5  (
            .in0(N__44651),
            .in1(N__38453),
            .in2(_gnd_net_),
            .in3(N__38431),
            .lcout(data_in_19_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50411),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i141_LC_10_32_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i141_LC_10_32_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i141_LC_10_32_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i141_LC_10_32_6  (
            .in0(N__44648),
            .in1(N__38536),
            .in2(_gnd_net_),
            .in3(N__38423),
            .lcout(data_in_17_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50411),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i139_LC_10_32_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i139_LC_10_32_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i139_LC_10_32_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i139_LC_10_32_7  (
            .in0(N__38414),
            .in1(N__44650),
            .in2(_gnd_net_),
            .in3(N__38398),
            .lcout(data_in_17_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50411),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i69_LC_11_20_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i69_LC_11_20_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i69_LC_11_20_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i69_LC_11_20_0  (
            .in0(N__38347),
            .in1(N__45212),
            .in2(_gnd_net_),
            .in3(N__38364),
            .lcout(data_in_8_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50321),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i77_LC_11_20_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i77_LC_11_20_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i77_LC_11_20_1 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i77_LC_11_20_1  (
            .in0(N__38326),
            .in1(_gnd_net_),
            .in2(N__45342),
            .in3(N__38346),
            .lcout(data_in_9_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50321),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i85_LC_11_20_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i85_LC_11_20_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i85_LC_11_20_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i85_LC_11_20_2  (
            .in0(N__38309),
            .in1(N__45213),
            .in2(_gnd_net_),
            .in3(N__38325),
            .lcout(data_in_10_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50321),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i93_LC_11_20_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i93_LC_11_20_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i93_LC_11_20_3 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i93_LC_11_20_3  (
            .in0(N__38597),
            .in1(_gnd_net_),
            .in2(N__45343),
            .in3(N__38308),
            .lcout(data_in_11_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50321),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i101_LC_11_20_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i101_LC_11_20_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i101_LC_11_20_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i101_LC_11_20_4  (
            .in0(N__38588),
            .in1(N__45210),
            .in2(_gnd_net_),
            .in3(N__38596),
            .lcout(data_in_12_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50321),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i109_LC_11_20_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i109_LC_11_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i109_LC_11_20_5 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_in_0___i109_LC_11_20_5  (
            .in0(N__38579),
            .in1(_gnd_net_),
            .in2(N__45341),
            .in3(N__38587),
            .lcout(data_in_13_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50321),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i117_LC_11_20_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i117_LC_11_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i117_LC_11_20_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i117_LC_11_20_6  (
            .in0(N__38558),
            .in1(N__45211),
            .in2(_gnd_net_),
            .in3(N__38578),
            .lcout(data_in_14_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50321),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i92_LC_11_21_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i92_LC_11_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i92_LC_11_21_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i92_LC_11_21_1  (
            .in0(N__45196),
            .in1(N__38569),
            .in2(_gnd_net_),
            .in3(N__38828),
            .lcout(data_in_11_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50332),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i125_LC_11_21_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i125_LC_11_21_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i125_LC_11_21_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i125_LC_11_21_4  (
            .in0(N__45209),
            .in1(N__38557),
            .in2(_gnd_net_),
            .in3(N__38525),
            .lcout(data_in_15_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50332),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i133_LC_11_22_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i133_LC_11_22_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i133_LC_11_22_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i133_LC_11_22_0  (
            .in0(N__45158),
            .in1(N__38524),
            .in2(_gnd_net_),
            .in3(N__38546),
            .lcout(data_in_16_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50341),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i34_LC_11_22_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i34_LC_11_22_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i34_LC_11_22_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_0___i34_LC_11_22_1  (
            .in0(N__39885),
            .in1(N__38493),
            .in2(_gnd_net_),
            .in3(N__45159),
            .lcout(data_in_4_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50341),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15747_2_lut_LC_11_22_2 .C_ON=1'b0;
    defparam \c0.i15747_2_lut_LC_11_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i15747_2_lut_LC_11_22_2 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \c0.i15747_2_lut_LC_11_22_2  (
            .in0(_gnd_net_),
            .in1(N__41797),
            .in2(_gnd_net_),
            .in3(N__48397),
            .lcout(),
            .ltout(\c0.n18089_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18426_bdd_4_lut_LC_11_22_3 .C_ON=1'b0;
    defparam \c0.n18426_bdd_4_lut_LC_11_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.n18426_bdd_4_lut_LC_11_22_3 .LUT_INIT=16'b1100110010111000;
    LogicCell40 \c0.n18426_bdd_4_lut_LC_11_22_3  (
            .in0(N__43973),
            .in1(N__38678),
            .in2(N__38477),
            .in3(N__48109),
            .lcout(),
            .ltout(\c0.n18429_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11402_4_lut_LC_11_22_4 .C_ON=1'b0;
    defparam \c0.i11402_4_lut_LC_11_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i11402_4_lut_LC_11_22_4 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \c0.i11402_4_lut_LC_11_22_4  (
            .in0(N__44063),
            .in1(N__48845),
            .in2(N__38693),
            .in3(N__48754),
            .lcout(tx_data_7_N_keep),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15753_2_lut_LC_11_22_6 .C_ON=1'b0;
    defparam \c0.i15753_2_lut_LC_11_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.i15753_2_lut_LC_11_22_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i15753_2_lut_LC_11_22_6  (
            .in0(_gnd_net_),
            .in1(N__45662),
            .in2(_gnd_net_),
            .in3(N__48396),
            .lcout(),
            .ltout(\c0.n18017_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_16021_LC_11_22_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_16021_LC_11_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_16021_LC_11_22_7 .LUT_INIT=16'b1011101111000000;
    LogicCell40 \c0.byte_transmit_counter_1__bdd_4_lut_16021_LC_11_22_7  (
            .in0(N__39395),
            .in1(N__48108),
            .in2(N__38681),
            .in3(N__47981),
            .lcout(\c0.n18426 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i140_LC_11_23_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i140_LC_11_23_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i140_LC_11_23_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i140_LC_11_23_0  (
            .in0(N__44950),
            .in1(N__38671),
            .in2(_gnd_net_),
            .in3(N__38852),
            .lcout(data_in_17_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50351),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15935_LC_11_23_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15935_LC_11_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15935_LC_11_23_1 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter_1__bdd_4_lut_15935_LC_11_23_1  (
            .in0(N__40874),
            .in1(N__48080),
            .in2(N__38660),
            .in3(N__47982),
            .lcout(),
            .ltout(\c0.n18378_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18378_bdd_4_lut_LC_11_23_2 .C_ON=1'b0;
    defparam \c0.n18378_bdd_4_lut_LC_11_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.n18378_bdd_4_lut_LC_11_23_2 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n18378_bdd_4_lut_LC_11_23_2  (
            .in0(N__48081),
            .in1(N__41351),
            .in2(N__38645),
            .in3(N__40655),
            .lcout(),
            .ltout(\c0.n18381_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11425_4_lut_LC_11_23_3 .C_ON=1'b0;
    defparam \c0.i11425_4_lut_LC_11_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i11425_4_lut_LC_11_23_3 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \c0.i11425_4_lut_LC_11_23_3  (
            .in0(N__43157),
            .in1(N__48844),
            .in2(N__38642),
            .in3(N__48759),
            .lcout(tx_data_2_N_keep),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i156_LC_11_23_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i156_LC_11_23_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i156_LC_11_23_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i156_LC_11_23_4  (
            .in0(N__44952),
            .in1(N__38633),
            .in2(_gnd_net_),
            .in3(N__38860),
            .lcout(data_in_19_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50351),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i110_LC_11_23_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i110_LC_11_23_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i110_LC_11_23_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i110_LC_11_23_5  (
            .in0(N__45204),
            .in1(N__38608),
            .in2(_gnd_net_),
            .in3(N__39335),
            .lcout(data_in_13_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50351),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i148_LC_11_23_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i148_LC_11_23_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i148_LC_11_23_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i148_LC_11_23_6  (
            .in0(N__44951),
            .in1(N__38851),
            .in2(_gnd_net_),
            .in3(N__38861),
            .lcout(data_in_18_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50351),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i97_LC_11_24_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i97_LC_11_24_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i97_LC_11_24_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i97_LC_11_24_0  (
            .in0(N__45051),
            .in1(N__38842),
            .in2(_gnd_net_),
            .in3(N__39068),
            .lcout(data_in_12_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50361),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i100_LC_11_24_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i100_LC_11_24_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i100_LC_11_24_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i100_LC_11_24_1  (
            .in0(N__38824),
            .in1(N__45052),
            .in2(_gnd_net_),
            .in3(N__38702),
            .lcout(data_in_12_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50361),
            .ce(),
            .sr(_gnd_net_));
    defparam n18462_bdd_4_lut_LC_11_24_2.C_ON=1'b0;
    defparam n18462_bdd_4_lut_LC_11_24_2.SEQ_MODE=4'b0000;
    defparam n18462_bdd_4_lut_LC_11_24_2.LUT_INIT=16'b1111101000001100;
    LogicCell40 n18462_bdd_4_lut_LC_11_24_2 (
            .in0(N__42206),
            .in1(N__39368),
            .in2(N__39137),
            .in3(N__38813),
            .lcout(n18465),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i71_LC_11_24_3 .C_ON=1'b0;
    defparam \c0.data_in_0___i71_LC_11_24_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i71_LC_11_24_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_0___i71_LC_11_24_3  (
            .in0(N__38800),
            .in1(N__38743),
            .in2(_gnd_net_),
            .in3(N__45053),
            .lcout(data_in_8_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50361),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i126_LC_11_24_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i126_LC_11_24_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i126_LC_11_24_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i126_LC_11_24_4  (
            .in0(N__45050),
            .in1(N__39349),
            .in2(_gnd_net_),
            .in3(N__38732),
            .lcout(data_in_15_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50361),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_i0_i9_LC_11_24_5 .C_ON=1'b0;
    defparam \c0.delay_counter_i0_i9_LC_11_24_5 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_i0_i9_LC_11_24_5 .LUT_INIT=16'b1110010010100000;
    LogicCell40 \c0.delay_counter_i0_i9_LC_11_24_5  (
            .in0(N__42438),
            .in1(N__40019),
            .in2(N__41936),
            .in3(N__42579),
            .lcout(\c0.delay_counter_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50361),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_i0_i6_LC_11_24_6 .C_ON=1'b0;
    defparam \c0.delay_counter_i0_i6_LC_11_24_6 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_i0_i6_LC_11_24_6 .LUT_INIT=16'b1010101011000000;
    LogicCell40 \c0.delay_counter_i0_i6_LC_11_24_6  (
            .in0(N__41964),
            .in1(N__39941),
            .in2(N__42581),
            .in3(N__42437),
            .lcout(\c0.delay_counter_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50361),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i108_LC_11_24_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i108_LC_11_24_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i108_LC_11_24_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i108_LC_11_24_7  (
            .in0(N__45054),
            .in1(N__38701),
            .in2(_gnd_net_),
            .in3(N__38714),
            .lcout(data_in_13_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50361),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i138_LC_11_25_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i138_LC_11_25_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i138_LC_11_25_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i138_LC_11_25_1  (
            .in0(N__45115),
            .in1(N__38983),
            .in2(_gnd_net_),
            .in3(N__38873),
            .lcout(data_in_17_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50372),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_adj_924_LC_11_25_2 .C_ON=1'b0;
    defparam \c0.i1_3_lut_adj_924_LC_11_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_adj_924_LC_11_25_2 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \c0.i1_3_lut_adj_924_LC_11_25_2  (
            .in0(N__39800),
            .in1(N__41900),
            .in2(_gnd_net_),
            .in3(N__38996),
            .lcout(\c0.n17349 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15288_2_lut_LC_11_25_3.C_ON=1'b0;
    defparam i15288_2_lut_LC_11_25_3.SEQ_MODE=4'b0000;
    defparam i15288_2_lut_LC_11_25_3.LUT_INIT=16'b1111111111001100;
    LogicCell40 i15288_2_lut_LC_11_25_3 (
            .in0(_gnd_net_),
            .in1(N__41018),
            .in2(_gnd_net_),
            .in3(N__41048),
            .lcout(),
            .ltout(n17737_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i4_4_lut_adj_1137_LC_11_25_4.C_ON=1'b0;
    defparam i4_4_lut_adj_1137_LC_11_25_4.SEQ_MODE=4'b0000;
    defparam i4_4_lut_adj_1137_LC_11_25_4.LUT_INIT=16'b0000000100000000;
    LogicCell40 i4_4_lut_adj_1137_LC_11_25_4 (
            .in0(N__40981),
            .in1(N__42884),
            .in2(N__38999),
            .in3(N__41159),
            .lcout(n17312),
            .ltout(n17312_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_1144_LC_11_25_5.C_ON=1'b0;
    defparam i1_2_lut_adj_1144_LC_11_25_5.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_1144_LC_11_25_5.LUT_INIT=16'b0000000011110000;
    LogicCell40 i1_2_lut_adj_1144_LC_11_25_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38990),
            .in3(N__42263),
            .lcout(n14_adj_2615),
            .ltout(n14_adj_2615_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i5_LC_11_25_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i5_LC_11_25_6 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i5_LC_11_25_6 .LUT_INIT=16'b0100111001000100;
    LogicCell40 \c0.byte_transmit_counter__i5_LC_11_25_6  (
            .in0(N__42697),
            .in1(N__41320),
            .in2(N__38987),
            .in3(N__41306),
            .lcout(byte_transmit_counter_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50372),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i2_LC_11_25_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i2_LC_11_25_7 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i2_LC_11_25_7 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \c0.byte_transmit_counter__i2_LC_11_25_7  (
            .in0(N__43034),
            .in1(N__42696),
            .in2(N__48164),
            .in3(N__42729),
            .lcout(byte_transmit_counter_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50372),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i130_LC_11_26_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i130_LC_11_26_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i130_LC_11_26_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i130_LC_11_26_0  (
            .in0(N__38984),
            .in1(N__45056),
            .in2(_gnd_net_),
            .in3(N__38965),
            .lcout(data_in_16_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50379),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_i0_LC_11_26_1 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_i0_LC_11_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Bit_Index_i0_LC_11_26_1 .LUT_INIT=16'b1010101001000100;
    LogicCell40 \c0.tx.r_Bit_Index_i0_LC_11_26_1  (
            .in0(N__38905),
            .in1(N__40154),
            .in2(_gnd_net_),
            .in3(N__38954),
            .lcout(r_Bit_Index_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50379),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i146_LC_11_26_2 .C_ON=1'b0;
    defparam \c0.data_in_0___i146_LC_11_26_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i146_LC_11_26_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i146_LC_11_26_2  (
            .in0(N__45113),
            .in1(N__38872),
            .in2(_gnd_net_),
            .in3(N__39029),
            .lcout(data_in_18_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50379),
            .ce(),
            .sr(_gnd_net_));
    defparam n18438_bdd_4_lut_LC_11_26_3.C_ON=1'b0;
    defparam n18438_bdd_4_lut_LC_11_26_3.SEQ_MODE=4'b0000;
    defparam n18438_bdd_4_lut_LC_11_26_3.LUT_INIT=16'b1010101011100100;
    LogicCell40 n18438_bdd_4_lut_LC_11_26_3 (
            .in0(N__39143),
            .in1(N__43181),
            .in2(N__42797),
            .in3(N__39130),
            .lcout(n18441),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i105_LC_11_26_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i105_LC_11_26_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i105_LC_11_26_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0___i105_LC_11_26_4  (
            .in0(N__39064),
            .in1(N__45055),
            .in2(_gnd_net_),
            .in3(N__39179),
            .lcout(data_in_13_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50379),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i3_LC_11_26_5 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i3_LC_11_26_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i3_LC_11_26_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.tx.r_Tx_Data_i3_LC_11_26_5  (
            .in0(N__48642),
            .in1(N__39053),
            .in2(_gnd_net_),
            .in3(N__40514),
            .lcout(r_Tx_Data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50379),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i154_LC_11_26_6 .C_ON=1'b0;
    defparam \c0.data_in_0___i154_LC_11_26_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i154_LC_11_26_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i154_LC_11_26_6  (
            .in0(N__45114),
            .in1(N__39040),
            .in2(_gnd_net_),
            .in3(N__39028),
            .lcout(data_in_19_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50379),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i0_LC_11_26_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i0_LC_11_26_7 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i0_LC_11_26_7 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \c0.byte_transmit_counter__i0_LC_11_26_7  (
            .in0(N__43073),
            .in1(N__48377),
            .in2(N__42708),
            .in3(N__40054),
            .lcout(\c0.byte_transmit_counter_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50379),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i121_LC_11_27_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i121_LC_11_27_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i121_LC_11_27_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0___i121_LC_11_27_1  (
            .in0(N__39008),
            .in1(N__44946),
            .in2(_gnd_net_),
            .in3(N__39190),
            .lcout(data_in_15_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50388),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15801_2_lut_LC_11_27_2 .C_ON=1'b0;
    defparam \c0.i15801_2_lut_LC_11_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.i15801_2_lut_LC_11_27_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i15801_2_lut_LC_11_27_2  (
            .in0(_gnd_net_),
            .in1(N__45713),
            .in2(_gnd_net_),
            .in3(N__48306),
            .lcout(\c0.n17937 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Bit_Index_i2_LC_11_27_3 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_i2_LC_11_27_3 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Bit_Index_i2_LC_11_27_3 .LUT_INIT=16'b0000000001101010;
    LogicCell40 \c0.rx.r_Bit_Index_i2_LC_11_27_3  (
            .in0(N__39290),
            .in1(N__39320),
            .in2(N__40502),
            .in3(N__40472),
            .lcout(r_Bit_Index_2_adj_2625),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50388),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i129_LC_11_27_4 .C_ON=1'b0;
    defparam \c0.data_in_0___i129_LC_11_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i129_LC_11_27_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i129_LC_11_27_4  (
            .in0(N__44945),
            .in1(N__39007),
            .in2(_gnd_net_),
            .in3(N__39020),
            .lcout(data_in_16_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50388),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11225_4_lut_LC_11_27_6 .C_ON=1'b0;
    defparam \c0.i11225_4_lut_LC_11_27_6 .SEQ_MODE=4'b0000;
    defparam \c0.i11225_4_lut_LC_11_27_6 .LUT_INIT=16'b0011001000000010;
    LogicCell40 \c0.i11225_4_lut_LC_11_27_6  (
            .in0(N__39377),
            .in1(N__48837),
            .in2(N__48761),
            .in3(N__43202),
            .lcout(),
            .ltout(tx_data_0_N_keep_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i0_LC_11_27_7 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i0_LC_11_27_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i0_LC_11_27_7 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \c0.tx.r_Tx_Data_i0_LC_11_27_7  (
            .in0(_gnd_net_),
            .in1(N__48648),
            .in2(N__39371),
            .in3(N__39367),
            .lcout(r_Tx_Data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50388),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i118_LC_11_28_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i118_LC_11_28_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i118_LC_11_28_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i118_LC_11_28_0  (
            .in0(N__44767),
            .in1(N__39353),
            .in2(_gnd_net_),
            .in3(N__39331),
            .lcout(data_in_14_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50395),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_868_LC_11_28_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_868_LC_11_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_868_LC_11_28_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_868_LC_11_28_1  (
            .in0(N__40741),
            .in1(N__48592),
            .in2(_gnd_net_),
            .in3(N__43940),
            .lcout(\c0.n17465 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2428_2_lut_LC_11_28_2 .C_ON=1'b0;
    defparam \c0.rx.i2428_2_lut_LC_11_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2428_2_lut_LC_11_28_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.rx.i2428_2_lut_LC_11_28_2  (
            .in0(_gnd_net_),
            .in1(N__40444),
            .in2(_gnd_net_),
            .in3(N__39228),
            .lcout(n4958),
            .ltout(n4958_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i7504_3_lut_4_lut_LC_11_28_3 .C_ON=1'b0;
    defparam \c0.rx.i7504_3_lut_4_lut_LC_11_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i7504_3_lut_4_lut_LC_11_28_3 .LUT_INIT=16'b1000000011001100;
    LogicCell40 \c0.rx.i7504_3_lut_4_lut_LC_11_28_3  (
            .in0(N__39285),
            .in1(N__40496),
            .in2(N__39251),
            .in3(N__39718),
            .lcout(n9920),
            .ltout(n9920_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Bit_Index_i1_LC_11_28_4 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_i1_LC_11_28_4 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Bit_Index_i1_LC_11_28_4 .LUT_INIT=16'b0000011100001000;
    LogicCell40 \c0.rx.r_Bit_Index_i1_LC_11_28_4  (
            .in0(N__40497),
            .in1(N__40445),
            .in2(N__39248),
            .in3(N__39229),
            .lcout(r_Bit_Index_1_adj_2626),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50395),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i113_LC_11_28_5 .C_ON=1'b0;
    defparam \c0.data_in_0___i113_LC_11_28_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i113_LC_11_28_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i113_LC_11_28_5  (
            .in0(N__44902),
            .in1(N__39175),
            .in2(_gnd_net_),
            .in3(N__39194),
            .lcout(data_in_14_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50395),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_8__1__3532_LC_11_29_1 .C_ON=1'b0;
    defparam \c0.data_out_8__1__3532_LC_11_29_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_8__1__3532_LC_11_29_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \c0.data_out_8__1__3532_LC_11_29_1  (
            .in0(N__46031),
            .in1(_gnd_net_),
            .in2(N__39164),
            .in3(N__44481),
            .lcout(data_out_8_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50400),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_8__0__3533_LC_11_29_2 .C_ON=1'b0;
    defparam \c0.data_out_8__0__3533_LC_11_29_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_8__0__3533_LC_11_29_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_out_8__0__3533_LC_11_29_2  (
            .in0(N__47826),
            .in1(N__46030),
            .in2(_gnd_net_),
            .in3(N__39437),
            .lcout(data_out_8_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50400),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1062_LC_11_29_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1062_LC_11_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1062_LC_11_29_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1062_LC_11_29_3  (
            .in0(N__44474),
            .in1(N__47825),
            .in2(_gnd_net_),
            .in3(N__39484),
            .lcout(\c0.n8953 ),
            .ltout(\c0.n8953_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1044_LC_11_29_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1044_LC_11_29_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1044_LC_11_29_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1044_LC_11_29_4  (
            .in0(_gnd_net_),
            .in1(N__41657),
            .in2(N__39419),
            .in3(N__45597),
            .lcout(\c0.n17626 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_8__5__3528_LC_11_29_5 .C_ON=1'b0;
    defparam \c0.data_out_8__5__3528_LC_11_29_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_8__5__3528_LC_11_29_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_8__5__3528_LC_11_29_5  (
            .in0(N__46032),
            .in1(N__39416),
            .in2(_gnd_net_),
            .in3(N__49697),
            .lcout(data_out_8_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50400),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i5_3_lut_LC_11_29_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i5_3_lut_LC_11_29_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i5_3_lut_LC_11_29_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_7_i5_3_lut_LC_11_29_6  (
            .in0(N__48394),
            .in1(N__43527),
            .in2(_gnd_net_),
            .in3(N__47800),
            .lcout(\c0.n5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_882_LC_11_29_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_882_LC_11_29_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_882_LC_11_29_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_882_LC_11_29_7  (
            .in0(N__40693),
            .in1(N__47669),
            .in2(_gnd_net_),
            .in3(N__40740),
            .lcout(\c0.n17400 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_5__6__3551_LC_11_30_0 .C_ON=1'b0;
    defparam \c0.data_out_5__6__3551_LC_11_30_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_5__6__3551_LC_11_30_0 .LUT_INIT=16'b1111101100001011;
    LogicCell40 \c0.data_out_5__6__3551_LC_11_30_0  (
            .in0(N__49446),
            .in1(N__40643),
            .in2(N__46916),
            .in3(N__39383),
            .lcout(\c0.data_out_7__6__N_530 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50406),
            .ce(N__46546),
            .sr(_gnd_net_));
    defparam \c0.data_out_5__7__I_0_3654_2_lut_LC_11_30_1 .C_ON=1'b0;
    defparam \c0.data_out_5__7__I_0_3654_2_lut_LC_11_30_1 .SEQ_MODE=4'b0000;
    defparam \c0.data_out_5__7__I_0_3654_2_lut_LC_11_30_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.data_out_5__7__I_0_3654_2_lut_LC_11_30_1  (
            .in0(_gnd_net_),
            .in1(N__48569),
            .in2(_gnd_net_),
            .in3(N__45653),
            .lcout(\c0.data_out_7__1__N_626 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1003_LC_11_30_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1003_LC_11_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1003_LC_11_30_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1003_LC_11_30_2  (
            .in0(N__45654),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45914),
            .lcout(\c0.n17665 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i13_4_lut_4_lut_LC_11_30_3 .C_ON=1'b0;
    defparam \c0.rx.i13_4_lut_4_lut_LC_11_30_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i13_4_lut_4_lut_LC_11_30_3 .LUT_INIT=16'b0100000000001111;
    LogicCell40 \c0.rx.i13_4_lut_4_lut_LC_11_30_3  (
            .in0(N__39773),
            .in1(N__39641),
            .in2(N__39719),
            .in3(N__39588),
            .lcout(\c0.rx.n9553 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_4_lut_4_lut_LC_11_30_4 .C_ON=1'b0;
    defparam \c0.rx.i1_4_lut_4_lut_LC_11_30_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_4_lut_4_lut_LC_11_30_4 .LUT_INIT=16'b0001000000010001;
    LogicCell40 \c0.rx.i1_4_lut_4_lut_LC_11_30_4  (
            .in0(N__39587),
            .in1(N__39772),
            .in2(N__39650),
            .in3(N__39713),
            .lcout(n9646),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i15891_2_lut_3_lut_LC_11_30_6 .C_ON=1'b0;
    defparam \c0.rx.i15891_2_lut_3_lut_LC_11_30_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i15891_2_lut_3_lut_LC_11_30_6 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \c0.rx.i15891_2_lut_3_lut_LC_11_30_6  (
            .in0(N__39589),
            .in1(N__39774),
            .in2(_gnd_net_),
            .in3(N__39712),
            .lcout(\c0.rx.n17351 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_adj_815_LC_11_30_7 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_adj_815_LC_11_30_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_adj_815_LC_11_30_7 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \c0.rx.i1_2_lut_adj_815_LC_11_30_7  (
            .in0(_gnd_net_),
            .in1(N__39710),
            .in2(_gnd_net_),
            .in3(N__39586),
            .lcout(\c0.rx.n17376 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__2__I_596_2_lut_LC_11_31_0 .C_ON=1'b0;
    defparam \c0.data_out_6__2__I_596_2_lut_LC_11_31_0 .SEQ_MODE=4'b0000;
    defparam \c0.data_out_6__2__I_596_2_lut_LC_11_31_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.data_out_6__2__I_596_2_lut_LC_11_31_0  (
            .in0(N__44139),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43803),
            .lcout(\c0.data_out_6__2__N_803 ),
            .ltout(\c0.data_out_6__2__N_803_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.mux_832_i1_4_lut_LC_11_31_1 .C_ON=1'b0;
    defparam \c0.mux_832_i1_4_lut_LC_11_31_1 .SEQ_MODE=4'b0000;
    defparam \c0.mux_832_i1_4_lut_LC_11_31_1 .LUT_INIT=16'b0000111101100110;
    LogicCell40 \c0.mux_832_i1_4_lut_LC_11_31_1  (
            .in0(N__49790),
            .in1(N__43132),
            .in2(N__39509),
            .in3(N__49447),
            .lcout(),
            .ltout(\c0.n2216_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__2__3547_LC_11_31_2 .C_ON=1'b0;
    defparam \c0.data_out_6__2__3547_LC_11_31_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__2__3547_LC_11_31_2 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \c0.data_out_6__2__3547_LC_11_31_2  (
            .in0(N__47415),
            .in1(N__39506),
            .in2(N__39488),
            .in3(N__46889),
            .lcout(\c0.data_out_6_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50412),
            .ce(N__46538),
            .sr(_gnd_net_));
    defparam \c0.i15712_2_lut_LC_11_31_3 .C_ON=1'b0;
    defparam \c0.i15712_2_lut_LC_11_31_3 .SEQ_MODE=4'b0000;
    defparam \c0.i15712_2_lut_LC_11_31_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i15712_2_lut_LC_11_31_3  (
            .in0(_gnd_net_),
            .in1(N__39467),
            .in2(_gnd_net_),
            .in3(N__47414),
            .lcout(),
            .ltout(\c0.n17964_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_5__2__3555_LC_11_31_4 .C_ON=1'b0;
    defparam \c0.data_out_5__2__3555_LC_11_31_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_5__2__3555_LC_11_31_4 .LUT_INIT=16'b1111000011101110;
    LogicCell40 \c0.data_out_5__2__3555_LC_11_31_4  (
            .in0(N__49448),
            .in1(N__39446),
            .in2(N__39440),
            .in3(N__46888),
            .lcout(\c0.data_out_5_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50412),
            .ce(N__46538),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_855_LC_11_31_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_855_LC_11_31_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_855_LC_11_31_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_855_LC_11_31_5  (
            .in0(N__46979),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41237),
            .lcout(\c0.n17525 ),
            .ltout(\c0.n17525_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_856_LC_11_31_6 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_856_LC_11_31_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_856_LC_11_31_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_856_LC_11_31_6  (
            .in0(N__40702),
            .in1(N__47644),
            .in2(N__39791),
            .in3(N__47579),
            .lcout(\c0.n17644 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_904_LC_11_31_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_904_LC_11_31_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_904_LC_11_31_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_904_LC_11_31_7  (
            .in0(N__46954),
            .in1(N__49846),
            .in2(_gnd_net_),
            .in3(N__43561),
            .lcout(\c0.n6_adj_2467 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_1__4__3585_LC_11_32_0 .C_ON=1'b0;
    defparam \c0.data_out_1__4__3585_LC_11_32_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_1__4__3585_LC_11_32_0 .LUT_INIT=16'b0000110001011100;
    LogicCell40 \c0.data_out_1__4__3585_LC_11_32_0  (
            .in0(N__49450),
            .in1(N__49867),
            .in2(N__46502),
            .in3(N__46884),
            .lcout(\c0.data_out_5__5__N_950 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50417),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_1__2__3587_LC_11_32_1 .C_ON=1'b0;
    defparam \c0.data_out_1__2__3587_LC_11_32_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_1__2__3587_LC_11_32_1 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \c0.data_out_1__2__3587_LC_11_32_1  (
            .in0(N__46882),
            .in1(N__46484),
            .in2(N__43770),
            .in3(N__49451),
            .lcout(data_out_1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50417),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_1__7__3582_LC_11_32_2 .C_ON=1'b0;
    defparam \c0.data_out_1__7__3582_LC_11_32_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_1__7__3582_LC_11_32_2 .LUT_INIT=16'b1111000001110010;
    LogicCell40 \c0.data_out_1__7__3582_LC_11_32_2  (
            .in0(N__47453),
            .in1(N__46883),
            .in2(N__41793),
            .in3(N__47136),
            .lcout(data_out_1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50417),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1061_LC_11_32_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1061_LC_11_32_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1061_LC_11_32_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1061_LC_11_32_4  (
            .in0(N__49615),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49651),
            .lcout(\c0.n8970 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_3__4__3569_LC_11_32_5 .C_ON=1'b0;
    defparam \c0.data_out_3__4__3569_LC_11_32_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_3__4__3569_LC_11_32_5 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \c0.data_out_3__4__3569_LC_11_32_5  (
            .in0(N__47137),
            .in1(N__41244),
            .in2(N__47498),
            .in3(N__47454),
            .lcout(data_out_3_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50417),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__5__3592_LC_11_32_6 .C_ON=1'b0;
    defparam \c0.data_out_0__5__3592_LC_11_32_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__5__3592_LC_11_32_6 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \c0.data_out_0__5__3592_LC_11_32_6  (
            .in0(N__47452),
            .in1(N__47135),
            .in2(N__43946),
            .in3(N__47494),
            .lcout(data_out_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50417),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_DV_52_LC_11_32_7 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_DV_52_LC_11_32_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_DV_52_LC_11_32_7 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \c0.rx.r_Rx_DV_52_LC_11_32_7  (
            .in0(N__39788),
            .in1(N__39779),
            .in2(N__44768),
            .in3(N__39717),
            .lcout(rx_data_ready),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50417),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i42_LC_12_19_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i42_LC_12_19_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i42_LC_12_19_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i42_LC_12_19_0  (
            .in0(N__45293),
            .in1(N__39878),
            .in2(_gnd_net_),
            .in3(N__39931),
            .lcout(data_in_5_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50322),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i87_LC_12_22_0 .C_ON=1'b0;
    defparam \c0.data_in_0___i87_LC_12_22_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i87_LC_12_22_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i87_LC_12_22_0  (
            .in0(N__45157),
            .in1(N__39812),
            .in2(_gnd_net_),
            .in3(N__39834),
            .lcout(data_in_10_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50352),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i43_4_lut_LC_12_22_1 .C_ON=1'b0;
    defparam \c0.i43_4_lut_LC_12_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i43_4_lut_LC_12_22_1 .LUT_INIT=16'b0011000000111010;
    LogicCell40 \c0.i43_4_lut_LC_12_22_1  (
            .in0(N__46795),
            .in1(N__40928),
            .in2(N__49308),
            .in3(N__42155),
            .lcout(\c0.n25_adj_2517 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_2_lut_3_lut_LC_12_22_5 .C_ON=1'b0;
    defparam \c0.i6_2_lut_3_lut_LC_12_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i6_2_lut_3_lut_LC_12_22_5 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \c0.i6_2_lut_3_lut_LC_12_22_5  (
            .in0(N__49244),
            .in1(N__46794),
            .in2(_gnd_net_),
            .in3(N__47342),
            .lcout(n9631),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_i0_i8_LC_12_23_0 .C_ON=1'b0;
    defparam \c0.delay_counter_i0_i8_LC_12_23_0 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_i0_i8_LC_12_23_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.delay_counter_i0_i8_LC_12_23_0  (
            .in0(N__40031),
            .in1(N__42329),
            .in2(_gnd_net_),
            .in3(N__42429),
            .lcout(\c0.delay_counter_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50362),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i95_LC_12_23_1 .C_ON=1'b0;
    defparam \c0.data_in_0___i95_LC_12_23_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i95_LC_12_23_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i95_LC_12_23_1  (
            .in0(N__45203),
            .in1(N__39811),
            .in2(_gnd_net_),
            .in3(N__40943),
            .lcout(data_in_11_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50362),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15306_4_lut_LC_12_23_3 .C_ON=1'b0;
    defparam \c0.i15306_4_lut_LC_12_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i15306_4_lut_LC_12_23_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i15306_4_lut_LC_12_23_3  (
            .in0(N__42300),
            .in1(N__42083),
            .in2(N__42334),
            .in3(N__41738),
            .lcout(\c0.n17755 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_i0_i10_LC_12_23_4 .C_ON=1'b0;
    defparam \c0.delay_counter_i0_i10_LC_12_23_4 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_i0_i10_LC_12_23_4 .LUT_INIT=16'b1010101011000000;
    LogicCell40 \c0.delay_counter_i0_i10_LC_12_23_4  (
            .in0(N__41739),
            .in1(N__42562),
            .in2(N__40010),
            .in3(N__42427),
            .lcout(\c0.delay_counter_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50362),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_i0_i3_LC_12_23_5 .C_ON=1'b0;
    defparam \c0.delay_counter_i0_i3_LC_12_23_5 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_i0_i3_LC_12_23_5 .LUT_INIT=16'b1101100010001000;
    LogicCell40 \c0.delay_counter_i0_i3_LC_12_23_5  (
            .in0(N__42428),
            .in1(N__41123),
            .in2(N__39959),
            .in3(N__42569),
            .lcout(\c0.delay_counter_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50362),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_adj_1021_LC_12_23_6 .C_ON=1'b0;
    defparam \c0.i1_3_lut_adj_1021_LC_12_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_adj_1021_LC_12_23_6 .LUT_INIT=16'b0101010111011101;
    LogicCell40 \c0.i1_3_lut_adj_1021_LC_12_23_6  (
            .in0(N__42656),
            .in1(N__39983),
            .in2(_gnd_net_),
            .in3(N__47283),
            .lcout(\c0.n1314 ),
            .ltout(\c0.n1314_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_i0_i2_LC_12_23_7 .C_ON=1'b0;
    defparam \c0.delay_counter_i0_i2_LC_12_23_7 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_i0_i2_LC_12_23_7 .LUT_INIT=16'b1111100000001000;
    LogicCell40 \c0.delay_counter_i0_i2_LC_12_23_7  (
            .in0(N__42561),
            .in1(N__39968),
            .in2(N__39977),
            .in3(N__41086),
            .lcout(\c0.delay_counter_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50362),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_3777_2_lut_LC_12_24_0 .C_ON=1'b1;
    defparam \c0.add_3777_2_lut_LC_12_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.add_3777_2_lut_LC_12_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_3777_2_lut_LC_12_24_0  (
            .in0(_gnd_net_),
            .in1(N__41043),
            .in2(_gnd_net_),
            .in3(N__39974),
            .lcout(\c0.n7275 ),
            .ltout(),
            .carryin(bfn_12_24_0_),
            .carryout(\c0.n16305 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_3777_3_lut_LC_12_24_1 .C_ON=1'b1;
    defparam \c0.add_3777_3_lut_LC_12_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_3777_3_lut_LC_12_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_3777_3_lut_LC_12_24_1  (
            .in0(_gnd_net_),
            .in1(N__41102),
            .in2(_gnd_net_),
            .in3(N__39971),
            .lcout(\c0.n7274 ),
            .ltout(),
            .carryin(\c0.n16305 ),
            .carryout(\c0.n16306 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_3777_4_lut_LC_12_24_2 .C_ON=1'b1;
    defparam \c0.add_3777_4_lut_LC_12_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_3777_4_lut_LC_12_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_3777_4_lut_LC_12_24_2  (
            .in0(_gnd_net_),
            .in1(N__41085),
            .in2(_gnd_net_),
            .in3(N__39962),
            .lcout(\c0.n7273 ),
            .ltout(),
            .carryin(\c0.n16306 ),
            .carryout(\c0.n16307 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_3777_5_lut_LC_12_24_3 .C_ON=1'b1;
    defparam \c0.add_3777_5_lut_LC_12_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_3777_5_lut_LC_12_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_3777_5_lut_LC_12_24_3  (
            .in0(_gnd_net_),
            .in1(N__41121),
            .in2(_gnd_net_),
            .in3(N__39950),
            .lcout(\c0.n7272 ),
            .ltout(),
            .carryin(\c0.n16307 ),
            .carryout(\c0.n16308 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_3777_6_lut_LC_12_24_4 .C_ON=1'b1;
    defparam \c0.add_3777_6_lut_LC_12_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_3777_6_lut_LC_12_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_3777_6_lut_LC_12_24_4  (
            .in0(_gnd_net_),
            .in1(N__41065),
            .in2(_gnd_net_),
            .in3(N__39947),
            .lcout(\c0.n7271 ),
            .ltout(),
            .carryin(\c0.n16308 ),
            .carryout(\c0.n16309 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_3777_7_lut_LC_12_24_5 .C_ON=1'b1;
    defparam \c0.add_3777_7_lut_LC_12_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_3777_7_lut_LC_12_24_5 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.add_3777_7_lut_LC_12_24_5  (
            .in0(N__42555),
            .in1(_gnd_net_),
            .in2(N__42302),
            .in3(N__39944),
            .lcout(\c0.n18012 ),
            .ltout(),
            .carryin(\c0.n16309 ),
            .carryout(\c0.n16310 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_3777_8_lut_LC_12_24_6 .C_ON=1'b1;
    defparam \c0.add_3777_8_lut_LC_12_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_3777_8_lut_LC_12_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_3777_8_lut_LC_12_24_6  (
            .in0(_gnd_net_),
            .in1(N__41960),
            .in2(_gnd_net_),
            .in3(N__39935),
            .lcout(\c0.n7269 ),
            .ltout(),
            .carryin(\c0.n16310 ),
            .carryout(\c0.n16311 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_3777_9_lut_LC_12_24_7 .C_ON=1'b1;
    defparam \c0.add_3777_9_lut_LC_12_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_3777_9_lut_LC_12_24_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_3777_9_lut_LC_12_24_7  (
            .in0(_gnd_net_),
            .in1(N__42380),
            .in2(_gnd_net_),
            .in3(N__40034),
            .lcout(\c0.n7268 ),
            .ltout(),
            .carryin(\c0.n16311 ),
            .carryout(\c0.n16312 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_3777_10_lut_LC_12_25_0 .C_ON=1'b1;
    defparam \c0.add_3777_10_lut_LC_12_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.add_3777_10_lut_LC_12_25_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.add_3777_10_lut_LC_12_25_0  (
            .in0(N__42575),
            .in1(N__42333),
            .in2(_gnd_net_),
            .in3(N__40022),
            .lcout(\c0.n18011 ),
            .ltout(),
            .carryin(bfn_12_25_0_),
            .carryout(\c0.n16313 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_3777_11_lut_LC_12_25_1 .C_ON=1'b1;
    defparam \c0.add_3777_11_lut_LC_12_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_3777_11_lut_LC_12_25_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_3777_11_lut_LC_12_25_1  (
            .in0(_gnd_net_),
            .in1(N__41927),
            .in2(_gnd_net_),
            .in3(N__40013),
            .lcout(\c0.n7266 ),
            .ltout(),
            .carryin(\c0.n16313 ),
            .carryout(\c0.n16314 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_3777_12_lut_LC_12_25_2 .C_ON=1'b1;
    defparam \c0.add_3777_12_lut_LC_12_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_3777_12_lut_LC_12_25_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_3777_12_lut_LC_12_25_2  (
            .in0(_gnd_net_),
            .in1(N__41743),
            .in2(_gnd_net_),
            .in3(N__39998),
            .lcout(\c0.n7265 ),
            .ltout(),
            .carryin(\c0.n16314 ),
            .carryout(\c0.n16315 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_3777_13_lut_LC_12_25_3 .C_ON=1'b1;
    defparam \c0.add_3777_13_lut_LC_12_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_3777_13_lut_LC_12_25_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_3777_13_lut_LC_12_25_3  (
            .in0(_gnd_net_),
            .in1(N__42355),
            .in2(_gnd_net_),
            .in3(N__39995),
            .lcout(\c0.n7264 ),
            .ltout(),
            .carryin(\c0.n16315 ),
            .carryout(\c0.n16316 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_3777_14_lut_LC_12_25_4 .C_ON=1'b1;
    defparam \c0.add_3777_14_lut_LC_12_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_3777_14_lut_LC_12_25_4 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.add_3777_14_lut_LC_12_25_4  (
            .in0(N__42574),
            .in1(N__42082),
            .in2(_gnd_net_),
            .in3(N__39992),
            .lcout(\c0.n18009 ),
            .ltout(),
            .carryin(\c0.n16316 ),
            .carryout(\c0.n16317 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_3777_15_lut_LC_12_25_5 .C_ON=1'b1;
    defparam \c0.add_3777_15_lut_LC_12_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_3777_15_lut_LC_12_25_5 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.add_3777_15_lut_LC_12_25_5  (
            .in0(N__42551),
            .in1(N__41009),
            .in2(_gnd_net_),
            .in3(N__39989),
            .lcout(\c0.n18008 ),
            .ltout(),
            .carryin(\c0.n16317 ),
            .carryout(\c0.n16318 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_3777_16_lut_LC_12_25_6 .C_ON=1'b0;
    defparam \c0.add_3777_16_lut_LC_12_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_3777_16_lut_LC_12_25_6 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \c0.add_3777_16_lut_LC_12_25_6  (
            .in0(N__40982),
            .in1(N__42552),
            .in2(_gnd_net_),
            .in3(N__39986),
            .lcout(\c0.n18105 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i7_LC_12_25_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i7_LC_12_25_7 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i7_LC_12_25_7 .LUT_INIT=16'b0011101000001010;
    LogicCell40 \c0.byte_transmit_counter__i7_LC_12_25_7  (
            .in0(N__41282),
            .in1(N__42730),
            .in2(N__42692),
            .in3(N__41267),
            .lcout(byte_transmit_counter_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50380),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i15852_3_lut_4_lut_4_lut_LC_12_26_0 .C_ON=1'b0;
    defparam \c0.tx.i15852_3_lut_4_lut_4_lut_LC_12_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i15852_3_lut_4_lut_4_lut_LC_12_26_0 .LUT_INIT=16'b1000001110000000;
    LogicCell40 \c0.tx.i15852_3_lut_4_lut_4_lut_LC_12_26_0  (
            .in0(N__40413),
            .in1(N__40239),
            .in2(N__40162),
            .in3(N__42984),
            .lcout(),
            .ltout(n4_adj_2653_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Active_47_LC_12_26_1 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Active_47_LC_12_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Active_47_LC_12_26_1 .LUT_INIT=16'b1010101000111010;
    LogicCell40 \c0.tx.r_Tx_Active_47_LC_12_26_1  (
            .in0(N__42914),
            .in1(N__40153),
            .in2(N__40379),
            .in3(N__40338),
            .lcout(tx_active),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50389),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i241_2_lut_LC_12_26_2 .C_ON=1'b0;
    defparam \c0.i241_2_lut_LC_12_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.i241_2_lut_LC_12_26_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.i241_2_lut_LC_12_26_2  (
            .in0(_gnd_net_),
            .in1(N__40061),
            .in2(_gnd_net_),
            .in3(N__42913),
            .lcout(\c0.n251 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i2_2_lut_3_lut_4_lut_LC_12_26_4 .C_ON=1'b0;
    defparam \c0.tx.i2_2_lut_3_lut_4_lut_LC_12_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i2_2_lut_3_lut_4_lut_LC_12_26_4 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \c0.tx.i2_2_lut_3_lut_4_lut_LC_12_26_4  (
            .in0(N__40337),
            .in1(N__40238),
            .in2(N__40161),
            .in3(N__42983),
            .lcout(n7734),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_active_prev_3508_LC_12_26_5 .C_ON=1'b0;
    defparam \c0.tx_active_prev_3508_LC_12_26_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx_active_prev_3508_LC_12_26_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \c0.tx_active_prev_3508_LC_12_26_5  (
            .in0(N__42915),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.tx_active_prev ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50389),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i1_LC_12_26_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i1_LC_12_26_6 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i1_LC_12_26_6 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \c0.byte_transmit_counter__i1_LC_12_26_6  (
            .in0(N__43052),
            .in1(N__47930),
            .in2(N__42707),
            .in3(N__40055),
            .lcout(\c0.byte_transmit_counter_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50389),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i2_3_lut_LC_12_26_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i2_3_lut_LC_12_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i2_3_lut_LC_12_26_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_5_i2_3_lut_LC_12_26_7  (
            .in0(N__46950),
            .in1(N__40847),
            .in2(_gnd_net_),
            .in3(N__48376),
            .lcout(\c0.n2_adj_2476 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15940_LC_12_27_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15940_LC_12_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15940_LC_12_27_0 .LUT_INIT=16'b1111100000111000;
    LogicCell40 \c0.byte_transmit_counter_1__bdd_4_lut_15940_LC_12_27_0  (
            .in0(N__40043),
            .in1(N__48106),
            .in2(N__47969),
            .in3(N__41384),
            .lcout(),
            .ltout(\c0.n18390_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18390_bdd_4_lut_LC_12_27_1 .C_ON=1'b0;
    defparam \c0.n18390_bdd_4_lut_LC_12_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.n18390_bdd_4_lut_LC_12_27_1 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n18390_bdd_4_lut_LC_12_27_1  (
            .in0(N__48107),
            .in1(N__41360),
            .in2(N__40037),
            .in3(N__40508),
            .lcout(),
            .ltout(\c0.n18393_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11421_4_lut_LC_12_27_2 .C_ON=1'b0;
    defparam \c0.i11421_4_lut_LC_12_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.i11421_4_lut_LC_12_27_2 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \c0.i11421_4_lut_LC_12_27_2  (
            .in0(N__45524),
            .in1(N__48815),
            .in2(N__40517),
            .in3(N__48755),
            .lcout(tx_data_3_N_keep),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15744_2_lut_LC_12_27_4 .C_ON=1'b0;
    defparam \c0.i15744_2_lut_LC_12_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.i15744_2_lut_LC_12_27_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \c0.i15744_2_lut_LC_12_27_4  (
            .in0(N__48313),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43408),
            .lcout(\c0.n18095 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i5_3_lut_LC_12_27_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i5_3_lut_LC_12_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i5_3_lut_LC_12_27_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_4_i5_3_lut_LC_12_27_5  (
            .in0(N__41656),
            .in1(N__43300),
            .in2(_gnd_net_),
            .in3(N__48312),
            .lcout(\c0.n5_adj_2447 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_LC_12_28_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_LC_12_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_LC_12_28_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_LC_12_28_0  (
            .in0(N__43407),
            .in1(N__40728),
            .in2(N__40697),
            .in3(N__46441),
            .lcout(\c0.n17641 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__1__I_638_2_lut_LC_12_28_1 .C_ON=1'b0;
    defparam \c0.data_out_6__1__I_638_2_lut_LC_12_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.data_out_6__1__I_638_2_lut_LC_12_28_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.data_out_6__1__I_638_2_lut_LC_12_28_1  (
            .in0(N__40848),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44013),
            .lcout(\c0.data_out_6__1__N_849 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Bit_Index_i0_LC_12_28_2 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_i0_LC_12_28_2 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Bit_Index_i0_LC_12_28_2 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \c0.rx.r_Bit_Index_i0_LC_12_28_2  (
            .in0(N__40501),
            .in1(N__40451),
            .in2(_gnd_net_),
            .in3(N__40471),
            .lcout(r_Bit_Index_0_adj_2627),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50401),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_2__0__3581_LC_12_28_3 .C_ON=1'b0;
    defparam \c0.data_out_2__0__3581_LC_12_28_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_2__0__3581_LC_12_28_3 .LUT_INIT=16'b1011111100010000;
    LogicCell40 \c0.data_out_2__0__3581_LC_12_28_3  (
            .in0(N__47039),
            .in1(N__46872),
            .in2(N__47465),
            .in3(N__40686),
            .lcout(data_out_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50401),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_834_LC_12_28_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_834_LC_12_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_834_LC_12_28_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_834_LC_12_28_4  (
            .in0(N__44014),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40849),
            .lcout(\c0.n17445 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15782_2_lut_LC_12_28_5 .C_ON=1'b0;
    defparam \c0.i15782_2_lut_LC_12_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.i15782_2_lut_LC_12_28_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.i15782_2_lut_LC_12_28_5  (
            .in0(_gnd_net_),
            .in1(N__40526),
            .in2(_gnd_net_),
            .in3(N__48395),
            .lcout(\c0.n18062 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_2__2__3579_LC_12_28_6 .C_ON=1'b0;
    defparam \c0.data_out_2__2__3579_LC_12_28_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_2__2__3579_LC_12_28_6 .LUT_INIT=16'b1100110001001110;
    LogicCell40 \c0.data_out_2__2__3579_LC_12_28_6  (
            .in0(N__47434),
            .in1(N__40729),
            .in2(N__46915),
            .in3(N__47040),
            .lcout(data_out_6__6__N_729),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50401),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_3__5__3568_LC_12_28_7 .C_ON=1'b0;
    defparam \c0.data_out_3__5__3568_LC_12_28_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_3__5__3568_LC_12_28_7 .LUT_INIT=16'b1010110010101010;
    LogicCell40 \c0.data_out_3__5__3568_LC_12_28_7  (
            .in0(N__46949),
            .in1(N__46873),
            .in2(N__47078),
            .in3(N__47435),
            .lcout(data_out_3_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50401),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_895_LC_12_29_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_895_LC_12_29_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_895_LC_12_29_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_895_LC_12_29_0  (
            .in0(N__47767),
            .in1(N__43949),
            .in2(N__43421),
            .in3(N__40850),
            .lcout(\c0.data_out_6__7__N_675 ),
            .ltout(\c0.data_out_6__7__N_675_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15683_3_lut_LC_12_29_1 .C_ON=1'b0;
    defparam \c0.i15683_3_lut_LC_12_29_1 .SEQ_MODE=4'b0000;
    defparam \c0.i15683_3_lut_LC_12_29_1 .LUT_INIT=16'b1000001010000010;
    LogicCell40 \c0.i15683_3_lut_LC_12_29_1  (
            .in0(N__49435),
            .in1(N__45658),
            .in2(N__40595),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\c0.n17928_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__7__3534_LC_12_29_2 .C_ON=1'b0;
    defparam \c0.data_out_7__7__3534_LC_12_29_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__7__3534_LC_12_29_2 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \c0.data_out_7__7__3534_LC_12_29_2  (
            .in0(N__47398),
            .in1(N__40592),
            .in2(N__40571),
            .in3(N__46871),
            .lcout(\c0.data_out_7_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50407),
            .ce(N__44187),
            .sr(_gnd_net_));
    defparam \c0.i15763_2_lut_LC_12_29_3 .C_ON=1'b0;
    defparam \c0.i15763_2_lut_LC_12_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.i15763_2_lut_LC_12_29_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i15763_2_lut_LC_12_29_3  (
            .in0(N__40568),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47397),
            .lcout(),
            .ltout(\c0.n17906_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__6__3535_LC_12_29_4 .C_ON=1'b0;
    defparam \c0.data_out_7__6__3535_LC_12_29_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__6__3535_LC_12_29_4 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \c0.data_out_7__6__3535_LC_12_29_4  (
            .in0(N__49383),
            .in1(N__40550),
            .in2(N__40541),
            .in3(N__46870),
            .lcout(\c0.data_out_7_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50407),
            .ce(N__44187),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_878_LC_12_29_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_878_LC_12_29_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_878_LC_12_29_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_878_LC_12_29_5  (
            .in0(N__48198),
            .in1(N__47799),
            .in2(_gnd_net_),
            .in3(N__41821),
            .lcout(\c0.n8950 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__2__3539_LC_12_29_7 .C_ON=1'b0;
    defparam \c0.data_out_7__2__3539_LC_12_29_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__2__3539_LC_12_29_7 .LUT_INIT=16'b1110101001000000;
    LogicCell40 \c0.data_out_7__2__3539_LC_12_29_7  (
            .in0(N__46869),
            .in1(N__43121),
            .in2(N__49449),
            .in3(N__40538),
            .lcout(\c0.data_out_7_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50407),
            .ce(N__44187),
            .sr(_gnd_net_));
    defparam \c0.data_out_10__6__3511_LC_12_30_0 .C_ON=1'b0;
    defparam \c0.data_out_10__6__3511_LC_12_30_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_10__6__3511_LC_12_30_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_10__6__3511_LC_12_30_0  (
            .in0(N__43945),
            .in1(N__40745),
            .in2(N__46219),
            .in3(N__48570),
            .lcout(\c0.data_out_10_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50413),
            .ce(N__46047),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_2_i2_3_lut_LC_12_30_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_2_i2_3_lut_LC_12_30_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_2_i2_3_lut_LC_12_30_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_2_i2_3_lut_LC_12_30_3  (
            .in0(N__40743),
            .in1(N__41623),
            .in2(_gnd_net_),
            .in3(N__48460),
            .lcout(\c0.n2_adj_2483 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_835_LC_12_30_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_835_LC_12_30_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_835_LC_12_30_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_835_LC_12_30_4  (
            .in0(_gnd_net_),
            .in1(N__44268),
            .in2(_gnd_net_),
            .in3(N__43651),
            .lcout(\c0.n8634 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1104_LC_12_30_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1104_LC_12_30_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1104_LC_12_30_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i2_3_lut_adj_1104_LC_12_30_5  (
            .in0(N__49866),
            .in1(_gnd_net_),
            .in2(N__41254),
            .in3(N__41624),
            .lcout(\c0.n17389 ),
            .ltout(\c0.n17389_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1052_LC_12_30_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1052_LC_12_30_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1052_LC_12_30_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1052_LC_12_30_6  (
            .in0(N__41541),
            .in1(N__43562),
            .in2(N__40637),
            .in3(N__45717),
            .lcout(\c0.n17600 ),
            .ltout(\c0.n17600_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.mux_728_i1_4_lut_LC_12_30_7 .C_ON=1'b0;
    defparam \c0.mux_728_i1_4_lut_LC_12_30_7 .SEQ_MODE=4'b0000;
    defparam \c0.mux_728_i1_4_lut_LC_12_30_7 .LUT_INIT=16'b1111000001100110;
    LogicCell40 \c0.mux_728_i1_4_lut_LC_12_30_7  (
            .in0(N__40744),
            .in1(N__43944),
            .in2(N__40634),
            .in3(N__49417),
            .lcout(\c0.n9658 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1060_LC_12_31_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1060_LC_12_31_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1060_LC_12_31_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1060_LC_12_31_0  (
            .in0(N__43750),
            .in1(N__41621),
            .in2(N__41546),
            .in3(N__44140),
            .lcout(\c0.n17398 ),
            .ltout(\c0.n17398_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.mux_780_i1_4_lut_LC_12_31_1 .C_ON=1'b0;
    defparam \c0.mux_780_i1_4_lut_LC_12_31_1 .SEQ_MODE=4'b0000;
    defparam \c0.mux_780_i1_4_lut_LC_12_31_1 .LUT_INIT=16'b0000111101100110;
    LogicCell40 \c0.mux_780_i1_4_lut_LC_12_31_1  (
            .in0(N__41689),
            .in1(N__46382),
            .in2(N__40619),
            .in3(N__49420),
            .lcout(),
            .ltout(\c0.n2146_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__4__3545_LC_12_31_2 .C_ON=1'b0;
    defparam \c0.data_out_6__4__3545_LC_12_31_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__4__3545_LC_12_31_2 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \c0.data_out_6__4__3545_LC_12_31_2  (
            .in0(N__47436),
            .in1(N__40616),
            .in2(N__40598),
            .in3(N__46896),
            .lcout(\c0.data_out_6_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50418),
            .ce(N__46557),
            .sr(_gnd_net_));
    defparam \c0.data_out_1__1__3588_LC_12_31_3 .C_ON=1'b0;
    defparam \c0.data_out_1__1__3588_LC_12_31_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_1__1__3588_LC_12_31_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \c0.data_out_1__1__3588_LC_12_31_3  (
            .in0(N__46894),
            .in1(N__49421),
            .in2(_gnd_net_),
            .in3(N__47437),
            .lcout(\c0.data_out_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50418),
            .ce(N__46557),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1088_LC_12_31_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1088_LC_12_31_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1088_LC_12_31_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1088_LC_12_31_4  (
            .in0(N__43749),
            .in1(N__43796),
            .in2(_gnd_net_),
            .in3(N__44000),
            .lcout(\c0.data_out_5__3__N_964 ),
            .ltout(\c0.data_out_5__3__N_964_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1069_LC_12_31_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1069_LC_12_31_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1069_LC_12_31_5 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \c0.i1_2_lut_adj_1069_LC_12_31_5  (
            .in0(_gnd_net_),
            .in1(N__43647),
            .in2(N__40772),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\c0.data_out_6__3__N_785_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.mux_806_i1_4_lut_LC_12_31_6 .C_ON=1'b0;
    defparam \c0.mux_806_i1_4_lut_LC_12_31_6 .SEQ_MODE=4'b0000;
    defparam \c0.mux_806_i1_4_lut_LC_12_31_6 .LUT_INIT=16'b1011000111100100;
    LogicCell40 \c0.mux_806_i1_4_lut_LC_12_31_6  (
            .in0(N__49419),
            .in1(N__45749),
            .in2(N__40769),
            .in3(N__49791),
            .lcout(),
            .ltout(\c0.n2181_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__3__3546_LC_12_31_7 .C_ON=1'b0;
    defparam \c0.data_out_6__3__3546_LC_12_31_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__3__3546_LC_12_31_7 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \c0.data_out_6__3__3546_LC_12_31_7  (
            .in0(N__46895),
            .in1(N__40766),
            .in2(N__40748),
            .in3(N__47438),
            .lcout(\c0.data_out_6_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50418),
            .ce(N__46557),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__6__3591_LC_12_32_0 .C_ON=1'b0;
    defparam \c0.data_out_0__6__3591_LC_12_32_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__6__3591_LC_12_32_0 .LUT_INIT=16'b0000010111001100;
    LogicCell40 \c0.data_out_0__6__3591_LC_12_32_0  (
            .in0(N__49422),
            .in1(N__47766),
            .in2(N__46918),
            .in3(N__46523),
            .lcout(\c0.data_out_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50423),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_3__2__3571_LC_12_32_1 .C_ON=1'b0;
    defparam \c0.data_out_3__2__3571_LC_12_32_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_3__2__3571_LC_12_32_1 .LUT_INIT=16'b1101110010001100;
    LogicCell40 \c0.data_out_3__2__3571_LC_12_32_1  (
            .in0(N__47126),
            .in1(N__41615),
            .in2(N__47461),
            .in3(N__47488),
            .lcout(data_out_5__4__N_959),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50423),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1067_LC_12_32_2 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1067_LC_12_32_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1067_LC_12_32_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1067_LC_12_32_2  (
            .in0(N__40742),
            .in1(N__43394),
            .in2(N__40703),
            .in3(N__41755),
            .lcout(\c0.n17653 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_2__3__3578_LC_12_32_3 .C_ON=1'b0;
    defparam \c0.data_out_2__3__3578_LC_12_32_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_2__3__3578_LC_12_32_3 .LUT_INIT=16'b0101000001110010;
    LogicCell40 \c0.data_out_2__3__3578_LC_12_32_3  (
            .in0(N__46524),
            .in1(N__46907),
            .in2(N__43409),
            .in3(N__49423),
            .lcout(\c0.data_out_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50423),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_2__7__3574_LC_12_32_4 .C_ON=1'b0;
    defparam \c0.data_out_2__7__3574_LC_12_32_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_2__7__3574_LC_12_32_4 .LUT_INIT=16'b1100010011001110;
    LogicCell40 \c0.data_out_2__7__3574_LC_12_32_4  (
            .in0(N__47450),
            .in1(N__43994),
            .in2(N__47141),
            .in3(N__46898),
            .lcout(data_out_6__1__N_850),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50423),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_2__5__3576_LC_12_32_5 .C_ON=1'b0;
    defparam \c0.data_out_2__5__3576_LC_12_32_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_2__5__3576_LC_12_32_5 .LUT_INIT=16'b1101000111110000;
    LogicCell40 \c0.data_out_2__5__3576_LC_12_32_5  (
            .in0(N__46897),
            .in1(N__47122),
            .in2(N__40846),
            .in3(N__47451),
            .lcout(data_out_6__7__N_678),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50423),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_990_LC_12_32_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_990_LC_12_32_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_990_LC_12_32_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_990_LC_12_32_7  (
            .in0(N__40831),
            .in1(N__44128),
            .in2(N__44001),
            .in3(N__41614),
            .lcout(\c0.n8964 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15704_4_lut_LC_13_21_0.C_ON=1'b0;
    defparam i15704_4_lut_LC_13_21_0.SEQ_MODE=4'b0000;
    defparam i15704_4_lut_LC_13_21_0.LUT_INIT=16'b0101010001010101;
    LogicCell40 i15704_4_lut_LC_13_21_0 (
            .in0(N__47295),
            .in1(N__42571),
            .in2(N__42893),
            .in3(N__42050),
            .lcout(n17958),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_889_LC_13_21_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_889_LC_13_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_889_LC_13_21_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i1_2_lut_adj_889_LC_13_21_4  (
            .in0(N__47296),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46799),
            .lcout(n2615),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1007_LC_13_22_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1007_LC_13_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1007_LC_13_22_0 .LUT_INIT=16'b1110000011110000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1007_LC_13_22_0  (
            .in0(N__42888),
            .in1(N__42570),
            .in2(N__41453),
            .in3(N__42049),
            .lcout(n8488),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1025_LC_13_22_1 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1025_LC_13_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1025_LC_13_22_1 .LUT_INIT=16'b0000111100001110;
    LogicCell40 \c0.i1_4_lut_adj_1025_LC_13_22_1  (
            .in0(N__43010),
            .in1(N__42839),
            .in2(N__42892),
            .in3(N__42184),
            .lcout(n96),
            .ltout(n96_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_LC_13_22_2 .C_ON=1'b0;
    defparam \c0.i13_4_lut_LC_13_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_LC_13_22_2 .LUT_INIT=16'b1111111001010100;
    LogicCell40 \c0.i13_4_lut_LC_13_22_2  (
            .in0(N__49253),
            .in1(N__47229),
            .in2(N__40814),
            .in3(N__42126),
            .lcout(n17709),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_1147_LC_13_22_3.C_ON=1'b0;
    defparam i1_3_lut_adj_1147_LC_13_22_3.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_1147_LC_13_22_3.LUT_INIT=16'b1010101000100010;
    LogicCell40 i1_3_lut_adj_1147_LC_13_22_3 (
            .in0(N__46788),
            .in1(N__41988),
            .in2(_gnd_net_),
            .in3(N__42108),
            .lcout(),
            .ltout(n47_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_1148_LC_13_22_4.C_ON=1'b0;
    defparam i1_4_lut_adj_1148_LC_13_22_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_1148_LC_13_22_4.LUT_INIT=16'b0101010101010001;
    LogicCell40 i1_4_lut_adj_1148_LC_13_22_4 (
            .in0(N__49254),
            .in1(N__40807),
            .in2(N__40811),
            .in3(N__42003),
            .lcout(),
            .ltout(n41_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.UART_TRANSMITTER_state_i0_i2_LC_13_22_5 .C_ON=1'b0;
    defparam \c0.UART_TRANSMITTER_state_i0_i2_LC_13_22_5 .SEQ_MODE=4'b1000;
    defparam \c0.UART_TRANSMITTER_state_i0_i2_LC_13_22_5 .LUT_INIT=16'b0000111000001111;
    LogicCell40 \c0.UART_TRANSMITTER_state_i0_i2_LC_13_22_5  (
            .in0(N__42004),
            .in1(N__40808),
            .in2(N__40796),
            .in3(N__40907),
            .lcout(UART_TRANSMITTER_state_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50363),
            .ce(),
            .sr(_gnd_net_));
    defparam i64_4_lut_LC_13_22_6.C_ON=1'b0;
    defparam i64_4_lut_LC_13_22_6.SEQ_MODE=4'b0000;
    defparam i64_4_lut_LC_13_22_6.LUT_INIT=16'b0011000010111000;
    LogicCell40 i64_4_lut_LC_13_22_6 (
            .in0(N__41989),
            .in1(N__46787),
            .in2(N__40916),
            .in3(N__42142),
            .lcout(n43),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_i0_i4_LC_13_23_0 .C_ON=1'b0;
    defparam \c0.delay_counter_i0_i4_LC_13_23_0 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_i0_i4_LC_13_23_0 .LUT_INIT=16'b1010101011000000;
    LogicCell40 \c0.delay_counter_i0_i4_LC_13_23_0  (
            .in0(N__41066),
            .in1(N__42567),
            .in2(N__40901),
            .in3(N__42430),
            .lcout(\c0.delay_counter_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50373),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__1__3596_LC_13_23_1 .C_ON=1'b0;
    defparam \c0.data_out_0__1__3596_LC_13_23_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__1__3596_LC_13_23_1 .LUT_INIT=16'b1010001110101010;
    LogicCell40 \c0.data_out_0__1__3596_LC_13_23_1  (
            .in0(N__47619),
            .in1(N__46789),
            .in2(N__47127),
            .in3(N__47241),
            .lcout(data_out_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50373),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_i0_i14_LC_13_23_3 .C_ON=1'b0;
    defparam \c0.delay_counter_i0_i14_LC_13_23_3 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_i0_i14_LC_13_23_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \c0.delay_counter_i0_i14_LC_13_23_3  (
            .in0(N__42431),
            .in1(_gnd_net_),
            .in2(N__40892),
            .in3(N__40974),
            .lcout(delay_counter_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50373),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_i0_i5_LC_13_23_4 .C_ON=1'b0;
    defparam \c0.delay_counter_i0_i5_LC_13_23_4 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_i0_i5_LC_13_23_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.delay_counter_i0_i5_LC_13_23_4  (
            .in0(N__40880),
            .in1(N__42301),
            .in2(_gnd_net_),
            .in3(N__42432),
            .lcout(\c0.delay_counter_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50373),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_1001_LC_13_23_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_1001_LC_13_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_1001_LC_13_23_5 .LUT_INIT=16'b0000000000001110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_1001_LC_13_23_5  (
            .in0(N__42838),
            .in1(N__42185),
            .in2(N__42985),
            .in3(N__42930),
            .lcout(\c0.n113 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15731_2_lut_LC_13_23_6 .C_ON=1'b0;
    defparam \c0.i15731_2_lut_LC_13_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i15731_2_lut_LC_13_23_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i15731_2_lut_LC_13_23_6  (
            .in0(_gnd_net_),
            .in1(N__43588),
            .in2(_gnd_net_),
            .in3(N__48426),
            .lcout(\c0.n17936 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_i0_i0_LC_13_24_1 .C_ON=1'b0;
    defparam \c0.delay_counter_i0_i0_LC_13_24_1 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_i0_i0_LC_13_24_1 .LUT_INIT=16'b1010101011001111;
    LogicCell40 \c0.delay_counter_i0_i0_LC_13_24_1  (
            .in0(N__41047),
            .in1(N__40865),
            .in2(N__42580),
            .in3(N__42433),
            .lcout(delay_counter_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50381),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_i0_i1_LC_13_24_2 .C_ON=1'b0;
    defparam \c0.delay_counter_i0_i1_LC_13_24_2 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_i0_i1_LC_13_24_2 .LUT_INIT=16'b1101100010001000;
    LogicCell40 \c0.delay_counter_i0_i1_LC_13_24_2  (
            .in0(N__42435),
            .in1(N__41101),
            .in2(N__40859),
            .in3(N__42566),
            .lcout(\c0.delay_counter_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50381),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_i0_i13_LC_13_24_3 .C_ON=1'b0;
    defparam \c0.delay_counter_i0_i13_LC_13_24_3 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_i0_i13_LC_13_24_3 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \c0.delay_counter_i0_i13_LC_13_24_3  (
            .in0(N__41132),
            .in1(_gnd_net_),
            .in2(N__41011),
            .in3(N__42436),
            .lcout(delay_counter_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50381),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_912_LC_13_24_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_912_LC_13_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_912_LC_13_24_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i3_4_lut_adj_912_LC_13_24_4  (
            .in0(N__41122),
            .in1(N__41100),
            .in2(N__41087),
            .in3(N__41064),
            .lcout(\c0.n17387 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1042_LC_13_24_5 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1042_LC_13_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1042_LC_13_24_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i4_4_lut_adj_1042_LC_13_24_5  (
            .in0(N__42224),
            .in1(N__41036),
            .in2(N__41010),
            .in3(N__40968),
            .lcout(n29),
            .ltout(n29_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_i0_i11_LC_13_24_6 .C_ON=1'b0;
    defparam \c0.delay_counter_i0_i11_LC_13_24_6 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_i0_i11_LC_13_24_6 .LUT_INIT=16'b1110101001000000;
    LogicCell40 \c0.delay_counter_i0_i11_LC_13_24_6  (
            .in0(N__42434),
            .in1(N__40952),
            .in2(N__40946),
            .in3(N__42356),
            .lcout(\c0.delay_counter_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50381),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i103_LC_13_24_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i103_LC_13_24_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i103_LC_13_24_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0___i103_LC_13_24_7  (
            .in0(N__45495),
            .in1(N__44540),
            .in2(_gnd_net_),
            .in3(N__40942),
            .lcout(data_in_12_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50381),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i149_2_lut_3_lut_LC_13_25_0 .C_ON=1'b0;
    defparam \c0.i149_2_lut_3_lut_LC_13_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.i149_2_lut_3_lut_LC_13_25_0 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \c0.i149_2_lut_3_lut_LC_13_25_0  (
            .in0(N__43069),
            .in1(N__43051),
            .in2(_gnd_net_),
            .in3(N__43027),
            .lcout(\c0.n149 ),
            .ltout(\c0.n149_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_adj_915_LC_13_25_1 .C_ON=1'b0;
    defparam \c0.i1_3_lut_adj_915_LC_13_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_adj_915_LC_13_25_1 .LUT_INIT=16'b1111111110100000;
    LogicCell40 \c0.i1_3_lut_adj_915_LC_13_25_1  (
            .in0(N__42828),
            .in1(_gnd_net_),
            .in2(N__40931),
            .in3(N__42175),
            .lcout(n119),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1019_LC_13_25_2 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1019_LC_13_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1019_LC_13_25_2 .LUT_INIT=16'b0011001000100010;
    LogicCell40 \c0.i1_4_lut_adj_1019_LC_13_25_2  (
            .in0(N__42176),
            .in1(N__42870),
            .in2(N__42590),
            .in3(N__42829),
            .lcout(\c0.n93 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1126_LC_13_25_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1126_LC_13_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1126_LC_13_25_3 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1126_LC_13_25_3  (
            .in0(N__46627),
            .in1(N__47242),
            .in2(_gnd_net_),
            .in3(N__42240),
            .lcout(n8529),
            .ltout(n8529_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_917_LC_13_25_4 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_917_LC_13_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_917_LC_13_25_4 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \c0.i2_4_lut_adj_917_LC_13_25_4  (
            .in0(N__49255),
            .in1(N__43002),
            .in2(N__41180),
            .in3(N__41174),
            .lcout(\c0.n16450 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_905_LC_13_25_5 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_905_LC_13_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_905_LC_13_25_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i3_4_lut_adj_905_LC_13_25_5  (
            .in0(N__41299),
            .in1(N__42628),
            .in2(N__41210),
            .in3(N__41266),
            .lcout(\c0.n8550 ),
            .ltout(\c0.n8550_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_908_LC_13_25_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_908_LC_13_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_908_LC_13_25_6 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \c0.i1_2_lut_adj_908_LC_13_25_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__41177),
            .in3(N__42827),
            .lcout(n121_adj_2606),
            .ltout(n121_adj_2606_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_LC_13_25_7.C_ON=1'b0;
    defparam i1_4_lut_LC_13_25_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_LC_13_25_7.LUT_INIT=16'b1110101010101010;
    LogicCell40 i1_4_lut_LC_13_25_7 (
            .in0(N__41423),
            .in1(N__41168),
            .in2(N__41162),
            .in3(N__49256),
            .lcout(n13_adj_2652),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_3776_2_lut_LC_13_26_0 .C_ON=1'b1;
    defparam \c0.add_3776_2_lut_LC_13_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.add_3776_2_lut_LC_13_26_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_3776_2_lut_LC_13_26_0  (
            .in0(_gnd_net_),
            .in1(N__41150),
            .in2(N__48398),
            .in3(_gnd_net_),
            .lcout(\c0.tx_transmit_N_2239_0 ),
            .ltout(),
            .carryin(bfn_13_26_0_),
            .carryout(\c0.n16350 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_3776_3_lut_LC_13_26_1 .C_ON=1'b1;
    defparam \c0.add_3776_3_lut_LC_13_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_3776_3_lut_LC_13_26_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_3776_3_lut_LC_13_26_1  (
            .in0(_gnd_net_),
            .in1(N__47890),
            .in2(_gnd_net_),
            .in3(N__41144),
            .lcout(\c0.tx_transmit_N_2239_1 ),
            .ltout(),
            .carryin(\c0.n16350 ),
            .carryout(\c0.n16351 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_3776_4_lut_LC_13_26_2 .C_ON=1'b1;
    defparam \c0.add_3776_4_lut_LC_13_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_3776_4_lut_LC_13_26_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_3776_4_lut_LC_13_26_2  (
            .in0(_gnd_net_),
            .in1(N__48112),
            .in2(_gnd_net_),
            .in3(N__41141),
            .lcout(tx_transmit_N_2239_2),
            .ltout(),
            .carryin(\c0.n16351 ),
            .carryout(\c0.n16352 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_3776_5_lut_LC_13_26_3 .C_ON=1'b1;
    defparam \c0.add_3776_5_lut_LC_13_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_3776_5_lut_LC_13_26_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_3776_5_lut_LC_13_26_3  (
            .in0(_gnd_net_),
            .in1(N__48720),
            .in2(_gnd_net_),
            .in3(N__41138),
            .lcout(tx_transmit_N_2239_3),
            .ltout(),
            .carryin(\c0.n16352 ),
            .carryout(\c0.n16353 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_3776_6_lut_LC_13_26_4 .C_ON=1'b1;
    defparam \c0.add_3776_6_lut_LC_13_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_3776_6_lut_LC_13_26_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_3776_6_lut_LC_13_26_4  (
            .in0(_gnd_net_),
            .in1(N__48804),
            .in2(_gnd_net_),
            .in3(N__41135),
            .lcout(tx_transmit_N_2239_4),
            .ltout(),
            .carryin(\c0.n16353 ),
            .carryout(\c0.n16354 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_3776_7_lut_LC_13_26_5 .C_ON=1'b1;
    defparam \c0.add_3776_7_lut_LC_13_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_3776_7_lut_LC_13_26_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_3776_7_lut_LC_13_26_5  (
            .in0(_gnd_net_),
            .in1(N__41324),
            .in2(_gnd_net_),
            .in3(N__41288),
            .lcout(tx_transmit_N_2239_5),
            .ltout(),
            .carryin(\c0.n16354 ),
            .carryout(\c0.n16355 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_3776_8_lut_LC_13_26_6 .C_ON=1'b1;
    defparam \c0.add_3776_8_lut_LC_13_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_3776_8_lut_LC_13_26_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_3776_8_lut_LC_13_26_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42617),
            .in3(N__41285),
            .lcout(tx_transmit_N_2239_6),
            .ltout(),
            .carryin(\c0.n16355 ),
            .carryout(\c0.n16356 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_3776_9_lut_LC_13_26_7 .C_ON=1'b0;
    defparam \c0.add_3776_9_lut_LC_13_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_3776_9_lut_LC_13_26_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_3776_9_lut_LC_13_26_7  (
            .in0(_gnd_net_),
            .in1(N__41281),
            .in2(_gnd_net_),
            .in3(N__41270),
            .lcout(tx_transmit_N_2239_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15743_2_lut_LC_13_27_0 .C_ON=1'b0;
    defparam \c0.i15743_2_lut_LC_13_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.i15743_2_lut_LC_13_27_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i15743_2_lut_LC_13_27_0  (
            .in0(N__48401),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41255),
            .lcout(),
            .ltout(\c0.n18093_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18396_bdd_4_lut_LC_13_27_1 .C_ON=1'b0;
    defparam \c0.n18396_bdd_4_lut_LC_13_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.n18396_bdd_4_lut_LC_13_27_1 .LUT_INIT=16'b1100110011100010;
    LogicCell40 \c0.n18396_bdd_4_lut_LC_13_27_1  (
            .in0(N__41366),
            .in1(N__41186),
            .in2(N__41216),
            .in3(N__48133),
            .lcout(),
            .ltout(\c0.n18399_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11416_4_lut_LC_13_27_2 .C_ON=1'b0;
    defparam \c0.i11416_4_lut_LC_13_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.i11416_4_lut_LC_13_27_2 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \c0.i11416_4_lut_LC_13_27_2  (
            .in0(N__41390),
            .in1(N__48811),
            .in2(N__41213),
            .in3(N__48724),
            .lcout(tx_data_4_N_keep),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i4_LC_13_27_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i4_LC_13_27_3 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i4_LC_13_27_3 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \c0.byte_transmit_counter__i4_LC_13_27_3  (
            .in0(N__42749),
            .in1(N__42706),
            .in2(N__48833),
            .in3(N__41209),
            .lcout(byte_transmit_counter_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50402),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15689_2_lut_LC_13_27_4 .C_ON=1'b0;
    defparam \c0.i15689_2_lut_LC_13_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.i15689_2_lut_LC_13_27_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i15689_2_lut_LC_13_27_4  (
            .in0(N__48399),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43231),
            .lcout(),
            .ltout(\c0.n17941_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15945_LC_13_27_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15945_LC_13_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15945_LC_13_27_5 .LUT_INIT=16'b1011101111000000;
    LogicCell40 \c0.byte_transmit_counter_1__bdd_4_lut_15945_LC_13_27_5  (
            .in0(N__41195),
            .in1(N__48129),
            .in2(N__41189),
            .in3(N__47956),
            .lcout(\c0.n18396 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15796_4_lut_LC_13_27_6 .C_ON=1'b0;
    defparam \c0.i15796_4_lut_LC_13_27_6 .SEQ_MODE=4'b0000;
    defparam \c0.i15796_4_lut_LC_13_27_6 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \c0.i15796_4_lut_LC_13_27_6  (
            .in0(N__47957),
            .in1(N__41372),
            .in2(N__48156),
            .in3(N__44447),
            .lcout(\c0.n18068 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_3_i5_3_lut_LC_13_27_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_3_i5_3_lut_LC_13_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_3_i5_3_lut_LC_13_27_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_3_i5_3_lut_LC_13_27_7  (
            .in0(N__46086),
            .in1(N__43269),
            .in2(_gnd_net_),
            .in3(N__48400),
            .lcout(\c0.n5_adj_2490 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_10__4__3513_LC_13_28_0 .C_ON=1'b0;
    defparam \c0.data_out_10__4__3513_LC_13_28_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_10__4__3513_LC_13_28_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_10__4__3513_LC_13_28_0  (
            .in0(N__46087),
            .in1(N__41672),
            .in2(N__46365),
            .in3(N__43461),
            .lcout(\c0.data_out_10_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50408),
            .ce(N__46029),
            .sr(_gnd_net_));
    defparam \c0.i15822_2_lut_LC_13_28_1 .C_ON=1'b0;
    defparam \c0.i15822_2_lut_LC_13_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.i15822_2_lut_LC_13_28_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \c0.i15822_2_lut_LC_13_28_1  (
            .in0(N__48414),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41378),
            .lcout(\c0.n18067 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15742_2_lut_LC_13_28_2 .C_ON=1'b0;
    defparam \c0.i15742_2_lut_LC_13_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.i15742_2_lut_LC_13_28_2 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \c0.i15742_2_lut_LC_13_28_2  (
            .in0(_gnd_net_),
            .in1(N__49874),
            .in2(_gnd_net_),
            .in3(N__48411),
            .lcout(\c0.n18092 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15794_2_lut_LC_13_28_4 .C_ON=1'b0;
    defparam \c0.i15794_2_lut_LC_13_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.i15794_2_lut_LC_13_28_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \c0.i15794_2_lut_LC_13_28_4  (
            .in0(N__47696),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48412),
            .lcout(\c0.n18094 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15798_2_lut_LC_13_28_5 .C_ON=1'b0;
    defparam \c0.i15798_2_lut_LC_13_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.i15798_2_lut_LC_13_28_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i15798_2_lut_LC_13_28_5  (
            .in0(N__48413),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43772),
            .lcout(\c0.n18096 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15815_2_lut_LC_13_28_6 .C_ON=1'b0;
    defparam \c0.i15815_2_lut_LC_13_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.i15815_2_lut_LC_13_28_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i15815_2_lut_LC_13_28_6  (
            .in0(_gnd_net_),
            .in1(N__47577),
            .in2(_gnd_net_),
            .in3(N__48415),
            .lcout(\c0.n18088 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15875_2_lut_3_lut_4_lut_LC_13_29_0 .C_ON=1'b0;
    defparam \c0.i15875_2_lut_3_lut_4_lut_LC_13_29_0 .SEQ_MODE=4'b0000;
    defparam \c0.i15875_2_lut_3_lut_4_lut_LC_13_29_0 .LUT_INIT=16'b0000111000000000;
    LogicCell40 \c0.i15875_2_lut_3_lut_4_lut_LC_13_29_0  (
            .in0(N__46696),
            .in1(N__49322),
            .in2(N__47077),
            .in3(N__47300),
            .lcout(\c0.n9518 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11502_2_lut_3_lut_LC_13_29_1 .C_ON=1'b0;
    defparam \c0.i11502_2_lut_3_lut_LC_13_29_1 .SEQ_MODE=4'b0000;
    defparam \c0.i11502_2_lut_3_lut_LC_13_29_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.i11502_2_lut_3_lut_LC_13_29_1  (
            .in0(N__47299),
            .in1(N__49324),
            .in2(_gnd_net_),
            .in3(N__46695),
            .lcout(n4430),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_LC_13_29_2 .C_ON=1'b0;
    defparam \c0.i3_4_lut_LC_13_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_LC_13_29_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_LC_13_29_2  (
            .in0(N__43708),
            .in1(N__44046),
            .in2(N__48527),
            .in3(N__41759),
            .lcout(\c0.n9276 ),
            .ltout(\c0.n9276_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_827_LC_13_29_3 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_827_LC_13_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_827_LC_13_29_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_827_LC_13_29_3  (
            .in0(N__41545),
            .in1(N__44084),
            .in2(N__41525),
            .in3(N__45722),
            .lcout(\c0.n17623 ),
            .ltout(\c0.n17623_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15771_4_lut_LC_13_29_4 .C_ON=1'b0;
    defparam \c0.i15771_4_lut_LC_13_29_4 .SEQ_MODE=4'b0000;
    defparam \c0.i15771_4_lut_LC_13_29_4 .LUT_INIT=16'b0110100100000000;
    LogicCell40 \c0.i15771_4_lut_LC_13_29_4  (
            .in0(N__47529),
            .in1(N__41522),
            .in2(N__41510),
            .in3(N__49323),
            .lcout(),
            .ltout(\c0.n17916_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__0__3541_LC_13_29_5 .C_ON=1'b0;
    defparam \c0.data_out_7__0__3541_LC_13_29_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__0__3541_LC_13_29_5 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \c0.data_out_7__0__3541_LC_13_29_5  (
            .in0(N__47301),
            .in1(N__41507),
            .in2(N__41483),
            .in3(N__46697),
            .lcout(\c0.data_out_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50414),
            .ce(N__44173),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1055_LC_13_29_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1055_LC_13_29_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1055_LC_13_29_6 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1055_LC_13_29_6  (
            .in0(N__46694),
            .in1(N__49321),
            .in2(_gnd_net_),
            .in3(N__47298),
            .lcout(\c0.n8486 ),
            .ltout(\c0.n8486_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_920_LC_13_29_7 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_920_LC_13_29_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_920_LC_13_29_7 .LUT_INIT=16'b1111111101000000;
    LogicCell40 \c0.i1_4_lut_adj_920_LC_13_29_7  (
            .in0(N__42248),
            .in1(N__42047),
            .in2(N__41435),
            .in3(N__41432),
            .lcout(n4_adj_2612),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15690_2_lut_LC_13_30_0 .C_ON=1'b0;
    defparam \c0.i15690_2_lut_LC_13_30_0 .SEQ_MODE=4'b0000;
    defparam \c0.i15690_2_lut_LC_13_30_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i15690_2_lut_LC_13_30_0  (
            .in0(N__41411),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47402),
            .lcout(),
            .ltout(\c0.n17925_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__5__3536_LC_13_30_1 .C_ON=1'b0;
    defparam \c0.data_out_7__5__3536_LC_13_30_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__5__3536_LC_13_30_1 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \c0.data_out_7__5__3536_LC_13_30_1  (
            .in0(N__44368),
            .in1(N__49328),
            .in2(N__41393),
            .in3(N__46878),
            .lcout(\c0.data_out_7_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50419),
            .ce(N__44188),
            .sr(_gnd_net_));
    defparam \c0.i15673_2_lut_LC_13_30_2 .C_ON=1'b0;
    defparam \c0.i15673_2_lut_LC_13_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.i15673_2_lut_LC_13_30_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i15673_2_lut_LC_13_30_2  (
            .in0(_gnd_net_),
            .in1(N__41717),
            .in2(_gnd_net_),
            .in3(N__47401),
            .lcout(),
            .ltout(\c0.n17931_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__4__3537_LC_13_30_3 .C_ON=1'b0;
    defparam \c0.data_out_7__4__3537_LC_13_30_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__4__3537_LC_13_30_3 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \c0.data_out_7__4__3537_LC_13_30_3  (
            .in0(N__41668),
            .in1(N__49327),
            .in2(N__41699),
            .in3(N__46877),
            .lcout(\c0.data_out_7_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50419),
            .ce(N__44188),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_833_LC_13_30_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_833_LC_13_30_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_833_LC_13_30_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_833_LC_13_30_4  (
            .in0(_gnd_net_),
            .in1(N__41648),
            .in2(_gnd_net_),
            .in3(N__45590),
            .lcout(\c0.n8812 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_LC_13_30_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_LC_13_30_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_LC_13_30_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_LC_13_30_5  (
            .in0(N__43413),
            .in1(N__46448),
            .in2(N__47711),
            .in3(N__44051),
            .lcout(\c0.n17499 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_871_LC_13_30_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_871_LC_13_30_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_871_LC_13_30_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_871_LC_13_30_6  (
            .in0(N__46449),
            .in1(N__43230),
            .in2(N__41696),
            .in3(N__48526),
            .lcout(\c0.data_out_7__4__N_550 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_890_LC_13_30_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_890_LC_13_30_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_890_LC_13_30_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_890_LC_13_30_7  (
            .in0(N__41649),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46079),
            .lcout(\c0.n6_adj_2451 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15713_4_lut_LC_13_31_0 .C_ON=1'b0;
    defparam \c0.i15713_4_lut_LC_13_31_0 .SEQ_MODE=4'b0000;
    defparam \c0.i15713_4_lut_LC_13_31_0 .LUT_INIT=16'b1111011011111001;
    LogicCell40 \c0.i15713_4_lut_LC_13_31_0  (
            .in0(N__44123),
            .in1(N__41622),
            .in2(N__49445),
            .in3(N__43769),
            .lcout(),
            .ltout(\c0.n17967_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_5__4__3553_LC_13_31_1 .C_ON=1'b0;
    defparam \c0.data_out_5__4__3553_LC_13_31_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_5__4__3553_LC_13_31_1 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \c0.data_out_5__4__3553_LC_13_31_1  (
            .in0(N__41591),
            .in1(N__46899),
            .in2(N__41570),
            .in3(N__47404),
            .lcout(\c0.data_out_7__4__N_556 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50424),
            .ce(N__46564),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_1114_LC_13_31_2 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_1114_LC_13_31_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_1114_LC_13_31_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_1114_LC_13_31_2  (
            .in0(N__49808),
            .in1(N__43648),
            .in2(N__41567),
            .in3(N__41555),
            .lcout(\c0.n17662 ),
            .ltout(\c0.n17662_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.mux_702_i1_4_lut_LC_13_31_3 .C_ON=1'b0;
    defparam \c0.mux_702_i1_4_lut_LC_13_31_3 .SEQ_MODE=4'b0000;
    defparam \c0.mux_702_i1_4_lut_LC_13_31_3 .LUT_INIT=16'b0100111011100100;
    LogicCell40 \c0.mux_702_i1_4_lut_LC_13_31_3  (
            .in0(N__49418),
            .in1(N__45779),
            .in2(N__41888),
            .in3(N__49519),
            .lcout(),
            .ltout(\c0.n2041_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__7__3542_LC_13_31_4 .C_ON=1'b0;
    defparam \c0.data_out_6__7__3542_LC_13_31_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__7__3542_LC_13_31_4 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \c0.data_out_6__7__3542_LC_13_31_4  (
            .in0(N__47403),
            .in1(N__41885),
            .in2(N__41864),
            .in3(N__46914),
            .lcout(\c0.data_out_6_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50424),
            .ce(N__46564),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1084_LC_13_31_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1084_LC_13_31_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1084_LC_13_31_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1084_LC_13_31_5  (
            .in0(N__45625),
            .in1(N__48590),
            .in2(_gnd_net_),
            .in3(N__43226),
            .lcout(\c0.n17611 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_5__7__3550_LC_13_32_1 .C_ON=1'b0;
    defparam \c0.data_out_5__7__3550_LC_13_32_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_5__7__3550_LC_13_32_1 .LUT_INIT=16'b1111111000001110;
    LogicCell40 \c0.data_out_5__7__3550_LC_13_32_1  (
            .in0(N__49326),
            .in1(N__49730),
            .in2(N__46919),
            .in3(N__41861),
            .lcout(\c0.data_out_7__7__N_519 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50427),
            .ce(N__46565),
            .sr(_gnd_net_));
    defparam \c0.mux_884_i1_4_lut_LC_13_32_4 .C_ON=1'b0;
    defparam \c0.mux_884_i1_4_lut_LC_13_32_4 .SEQ_MODE=4'b0000;
    defparam \c0.mux_884_i1_4_lut_LC_13_32_4 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \c0.mux_884_i1_4_lut_LC_13_32_4  (
            .in0(N__47753),
            .in1(N__49325),
            .in2(N__47537),
            .in3(N__44069),
            .lcout(),
            .ltout(\c0.n17693_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__0__3549_LC_13_32_5 .C_ON=1'b0;
    defparam \c0.data_out_6__0__3549_LC_13_32_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__0__3549_LC_13_32_5 .LUT_INIT=16'b1000100000001111;
    LogicCell40 \c0.data_out_6__0__3549_LC_13_32_5  (
            .in0(N__47405),
            .in1(N__41849),
            .in2(N__41828),
            .in3(N__46900),
            .lcout(\c0.data_out_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50427),
            .ce(N__46565),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1123_LC_13_32_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1123_LC_13_32_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1123_LC_13_32_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_1123_LC_13_32_6  (
            .in0(N__41792),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43672),
            .lcout(\c0.n17578 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4518_2_lut_LC_14_22_0 .C_ON=1'b0;
    defparam \c0.i4518_2_lut_LC_14_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i4518_2_lut_LC_14_22_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i4518_2_lut_LC_14_22_0  (
            .in0(N__42573),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42127),
            .lcout(n6878),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_1039_LC_14_22_1 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_1039_LC_14_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_1039_LC_14_22_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i6_4_lut_adj_1039_LC_14_22_1  (
            .in0(N__42065),
            .in1(N__41935),
            .in2(N__41975),
            .in3(N__41744),
            .lcout(\c0.n14_adj_2533 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_3_lut_adj_1152_LC_14_22_3.C_ON=1'b0;
    defparam i2_3_lut_adj_1152_LC_14_22_3.SEQ_MODE=4'b0000;
    defparam i2_3_lut_adj_1152_LC_14_22_3.LUT_INIT=16'b0100010000000000;
    LogicCell40 i2_3_lut_adj_1152_LC_14_22_3 (
            .in0(N__47235),
            .in1(N__42572),
            .in2(_gnd_net_),
            .in3(N__42154),
            .lcout(n17364),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1030_LC_14_23_0 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1030_LC_14_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1030_LC_14_23_0 .LUT_INIT=16'b0111010101111111;
    LogicCell40 \c0.i1_4_lut_adj_1030_LC_14_23_0  (
            .in0(N__46785),
            .in1(N__42143),
            .in2(N__49364),
            .in3(N__42110),
            .lcout(),
            .ltout(n17672_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.UART_TRANSMITTER_state_i0_i0_LC_14_23_1 .C_ON=1'b0;
    defparam \c0.UART_TRANSMITTER_state_i0_i0_LC_14_23_1 .SEQ_MODE=4'b1000;
    defparam \c0.UART_TRANSMITTER_state_i0_i0_LC_14_23_1 .LUT_INIT=16'b1011101010001010;
    LogicCell40 \c0.UART_TRANSMITTER_state_i0_i0_LC_14_23_1  (
            .in0(N__47240),
            .in1(N__42778),
            .in2(N__42131),
            .in3(N__42011),
            .lcout(UART_TRANSMITTER_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50382),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5065_3_lut_4_lut_LC_14_23_2 .C_ON=1'b0;
    defparam \c0.i5065_3_lut_4_lut_LC_14_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5065_3_lut_4_lut_LC_14_23_2 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \c0.i5065_3_lut_4_lut_LC_14_23_2  (
            .in0(N__42553),
            .in1(N__42128),
            .in2(N__49363),
            .in3(N__42109),
            .lcout(\c0.n7428 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_i0_i12_LC_14_23_3 .C_ON=1'b0;
    defparam \c0.delay_counter_i0_i12_LC_14_23_3 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_i0_i12_LC_14_23_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.delay_counter_i0_i12_LC_14_23_3  (
            .in0(N__42448),
            .in1(N__42095),
            .in2(_gnd_net_),
            .in3(N__42081),
            .lcout(\c0.delay_counter_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50382),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_1005_LC_14_23_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_1005_LC_14_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_1005_LC_14_23_4 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_1005_LC_14_23_4  (
            .in0(N__42932),
            .in1(N__42554),
            .in2(N__42986),
            .in3(N__42048),
            .lcout(),
            .ltout(UART_TRANSMITTER_state_7_N_1749_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15721_4_lut_LC_14_23_5.C_ON=1'b0;
    defparam i15721_4_lut_LC_14_23_5.SEQ_MODE=4'b0000;
    defparam i15721_4_lut_LC_14_23_5.LUT_INIT=16'b0000000001010001;
    LogicCell40 i15721_4_lut_LC_14_23_5 (
            .in0(N__46724),
            .in1(N__49304),
            .in2(N__42014),
            .in3(N__47236),
            .lcout(n18032),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_1027_LC_14_23_7 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_1027_LC_14_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_1027_LC_14_23_7 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \c0.i2_4_lut_adj_1027_LC_14_23_7  (
            .in0(N__46723),
            .in1(N__42005),
            .in2(N__47142),
            .in3(N__41990),
            .lcout(n16485),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15304_4_lut_LC_14_24_1 .C_ON=1'b0;
    defparam \c0.i15304_4_lut_LC_14_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.i15304_4_lut_LC_14_24_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i15304_4_lut_LC_14_24_1  (
            .in0(N__42379),
            .in1(N__42354),
            .in2(N__41974),
            .in3(N__41931),
            .lcout(\c0.n17753 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_i0_i7_LC_14_24_2 .C_ON=1'b0;
    defparam \c0.delay_counter_i0_i7_LC_14_24_2 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_i0_i7_LC_14_24_2 .LUT_INIT=16'b1010101011000000;
    LogicCell40 \c0.delay_counter_i0_i7_LC_14_24_2  (
            .in0(N__42375),
            .in1(N__42568),
            .in2(N__42461),
            .in3(N__42449),
            .lcout(\c0.delay_counter_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50390),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_adj_1037_LC_14_24_3 .C_ON=1'b0;
    defparam \c0.i2_2_lut_adj_1037_LC_14_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_adj_1037_LC_14_24_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i2_2_lut_adj_1037_LC_14_24_3  (
            .in0(_gnd_net_),
            .in1(N__42374),
            .in2(_gnd_net_),
            .in3(N__42353),
            .lcout(),
            .ltout(\c0.n10_adj_2532_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_1040_LC_14_24_4 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_1040_LC_14_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_1040_LC_14_24_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i7_4_lut_adj_1040_LC_14_24_4  (
            .in0(N__42335),
            .in1(N__42296),
            .in2(N__42275),
            .in3(N__42272),
            .lcout(n17306),
            .ltout(n17306_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1041_LC_14_24_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1041_LC_14_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1041_LC_14_24_5 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \c0.i1_2_lut_adj_1041_LC_14_24_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42251),
            .in3(N__42241),
            .lcout(\c0.n6_adj_2534 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i4_LC_14_24_6 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i4_LC_14_24_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i4_LC_14_24_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.tx.r_Tx_Data_i4_LC_14_24_6  (
            .in0(N__48675),
            .in1(N__42205),
            .in2(_gnd_net_),
            .in3(N__42218),
            .lcout(r_Tx_Data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50390),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_adj_873_LC_14_25_0 .C_ON=1'b0;
    defparam \c0.i1_3_lut_adj_873_LC_14_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_adj_873_LC_14_25_0 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \c0.i1_3_lut_adj_873_LC_14_25_0  (
            .in0(N__49291),
            .in1(N__46672),
            .in2(_gnd_net_),
            .in3(N__43006),
            .lcout(),
            .ltout(\c0.n16_adj_2445_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_874_LC_14_25_1 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_874_LC_14_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_874_LC_14_25_1 .LUT_INIT=16'b0010001011110010;
    LogicCell40 \c0.i1_4_lut_adj_874_LC_14_25_1  (
            .in0(N__43079),
            .in1(N__42602),
            .in2(N__42191),
            .in3(N__42836),
            .lcout(),
            .ltout(\c0.n19_adj_2446_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_transmit_3509_LC_14_25_2 .C_ON=1'b0;
    defparam \c0.tx_transmit_3509_LC_14_25_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx_transmit_3509_LC_14_25_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \c0.tx_transmit_3509_LC_14_25_2  (
            .in0(N__47276),
            .in1(N__42874),
            .in2(N__42188),
            .in3(N__42183),
            .lcout(\c0.tx_transmit ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50396),
            .ce(),
            .sr(N__47144));
    defparam \c0.i11059_2_lut_LC_14_25_3 .C_ON=1'b0;
    defparam \c0.i11059_2_lut_LC_14_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.i11059_2_lut_LC_14_25_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \c0.i11059_2_lut_LC_14_25_3  (
            .in0(N__46671),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49290),
            .lcout(\c0.n2650 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1112_LC_14_25_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1112_LC_14_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1112_LC_14_25_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1112_LC_14_25_4  (
            .in0(N__43068),
            .in1(N__43050),
            .in2(_gnd_net_),
            .in3(N__43026),
            .lcout(\c0.n97 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11030_2_lut_LC_14_25_5 .C_ON=1'b0;
    defparam \c0.i11030_2_lut_LC_14_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.i11030_2_lut_LC_14_25_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i11030_2_lut_LC_14_25_5  (
            .in0(_gnd_net_),
            .in1(N__42950),
            .in2(_gnd_net_),
            .in3(N__42931),
            .lcout(n13415),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15888_2_lut_3_lut_LC_14_25_7 .C_ON=1'b0;
    defparam \c0.i15888_2_lut_3_lut_LC_14_25_7 .SEQ_MODE=4'b0000;
    defparam \c0.i15888_2_lut_3_lut_LC_14_25_7 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \c0.i15888_2_lut_3_lut_LC_14_25_7  (
            .in0(N__46670),
            .in1(N__49289),
            .in2(_gnd_net_),
            .in3(N__47275),
            .lcout(data_out_10__7__N_114),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i3_LC_14_26_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i3_LC_14_26_0 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i3_LC_14_26_0 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \c0.byte_transmit_counter__i3_LC_14_26_0  (
            .in0(N__48738),
            .in1(N__42837),
            .in2(N__42713),
            .in3(N__42744),
            .lcout(byte_transmit_counter_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50403),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i5_LC_14_26_1 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i5_LC_14_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i5_LC_14_26_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.tx.r_Tx_Data_i5_LC_14_26_1  (
            .in0(N__48661),
            .in1(N__42793),
            .in2(_gnd_net_),
            .in3(N__44339),
            .lcout(r_Tx_Data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50403),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.UART_TRANSMITTER_state_i0_i1_LC_14_26_2 .C_ON=1'b0;
    defparam \c0.UART_TRANSMITTER_state_i0_i1_LC_14_26_2 .SEQ_MODE=4'b1000;
    defparam \c0.UART_TRANSMITTER_state_i0_i1_LC_14_26_2 .LUT_INIT=16'b1101100111001000;
    LogicCell40 \c0.UART_TRANSMITTER_state_i0_i1_LC_14_26_2  (
            .in0(N__42779),
            .in1(N__46646),
            .in2(N__42764),
            .in3(N__47341),
            .lcout(UART_TRANSMITTER_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50403),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i6_LC_14_26_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i6_LC_14_26_3 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i6_LC_14_26_3 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \c0.byte_transmit_counter__i6_LC_14_26_3  (
            .in0(N__42745),
            .in1(N__42712),
            .in2(N__42635),
            .in3(N__42616),
            .lcout(byte_transmit_counter_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50403),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15292_2_lut_LC_14_26_4 .C_ON=1'b0;
    defparam \c0.i15292_2_lut_LC_14_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.i15292_2_lut_LC_14_26_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i15292_2_lut_LC_14_26_4  (
            .in0(_gnd_net_),
            .in1(N__46645),
            .in2(_gnd_net_),
            .in3(N__42601),
            .lcout(\c0.n17741 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i1_LC_14_26_5 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i1_LC_14_26_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i1_LC_14_26_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.tx.r_Tx_Data_i1_LC_14_26_5  (
            .in0(N__48660),
            .in1(N__43180),
            .in2(_gnd_net_),
            .in3(N__44318),
            .lcout(r_Tx_Data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50403),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_1_i1_3_lut_LC_14_26_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_1_i1_3_lut_LC_14_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_1_i1_3_lut_LC_14_26_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_1_i1_3_lut_LC_14_26_6  (
            .in0(N__47635),
            .in1(N__43810),
            .in2(_gnd_net_),
            .in3(N__48429),
            .lcout(\c0.n1_adj_2522 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15800_2_lut_LC_14_27_0 .C_ON=1'b0;
    defparam \c0.i15800_2_lut_LC_14_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.i15800_2_lut_LC_14_27_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \c0.i15800_2_lut_LC_14_27_0  (
            .in0(N__48417),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43106),
            .lcout(\c0.n18071 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_2_i8_3_lut_LC_14_27_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_2_i8_3_lut_LC_14_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_2_i8_3_lut_LC_14_27_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_2_i8_3_lut_LC_14_27_1  (
            .in0(N__43100),
            .in1(N__43333),
            .in2(_gnd_net_),
            .in3(N__48416),
            .lcout(),
            .ltout(\c0.n8_adj_2526_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15802_4_lut_LC_14_27_2 .C_ON=1'b0;
    defparam \c0.i15802_4_lut_LC_14_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.i15802_4_lut_LC_14_27_2 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \c0.i15802_4_lut_LC_14_27_2  (
            .in0(N__43166),
            .in1(N__48134),
            .in2(N__43160),
            .in3(N__47974),
            .lcout(\c0.n18072 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_858_LC_14_27_3 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_858_LC_14_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_858_LC_14_27_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_858_LC_14_27_3  (
            .in0(N__49792),
            .in1(N__48589),
            .in2(N__43145),
            .in3(N__43589),
            .lcout(\c0.data_out_7__2__N_574 ),
            .ltout(\c0.data_out_7__2__N_574_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_10__2__3515_LC_14_27_4 .C_ON=1'b0;
    defparam \c0.data_out_10__2__3515_LC_14_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_10__2__3515_LC_14_27_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_10__2__3515_LC_14_27_4  (
            .in0(N__43490),
            .in1(N__46310),
            .in2(N__43109),
            .in3(N__45834),
            .lcout(\c0.data_out_10_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50409),
            .ce(N__46008),
            .sr(_gnd_net_));
    defparam \c0.data_out_9__2__3523_LC_14_27_5 .C_ON=1'b0;
    defparam \c0.data_out_9__2__3523_LC_14_27_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_9__2__3523_LC_14_27_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.data_out_9__2__3523_LC_14_27_5  (
            .in0(N__43811),
            .in1(N__49637),
            .in2(_gnd_net_),
            .in3(N__44138),
            .lcout(\c0.data_out_9_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50409),
            .ce(N__46008),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_3_i8_3_lut_LC_14_28_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_3_i8_3_lut_LC_14_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_3_i8_3_lut_LC_14_28_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_3_i8_3_lut_LC_14_28_0  (
            .in0(N__43094),
            .in1(N__49566),
            .in2(_gnd_net_),
            .in3(N__48402),
            .lcout(\c0.n8_adj_2531 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15803_2_lut_LC_14_28_1 .C_ON=1'b0;
    defparam \c0.i15803_2_lut_LC_14_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.i15803_2_lut_LC_14_28_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \c0.i15803_2_lut_LC_14_28_1  (
            .in0(N__48403),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45800),
            .lcout(),
            .ltout(\c0.n18073_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15828_4_lut_LC_14_28_2 .C_ON=1'b0;
    defparam \c0.i15828_4_lut_LC_14_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.i15828_4_lut_LC_14_28_2 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \c0.i15828_4_lut_LC_14_28_2  (
            .in0(N__44453),
            .in1(N__48163),
            .in2(N__43358),
            .in3(N__47985),
            .lcout(\c0.n18014 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_8__3__3530_LC_14_28_3 .C_ON=1'b0;
    defparam \c0.data_out_8__3__3530_LC_14_28_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_8__3__3530_LC_14_28_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_out_8__3__3530_LC_14_28_3  (
            .in0(N__49567),
            .in1(N__46022),
            .in2(_gnd_net_),
            .in3(N__43355),
            .lcout(data_out_8_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50415),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1063_LC_14_28_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1063_LC_14_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1063_LC_14_28_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1063_LC_14_28_4  (
            .in0(N__43334),
            .in1(N__49565),
            .in2(_gnd_net_),
            .in3(N__43301),
            .lcout(\c0.n9091 ),
            .ltout(\c0.n9091_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1064_LC_14_28_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1064_LC_14_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1064_LC_14_28_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_1064_LC_14_28_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43280),
            .in3(N__43466),
            .lcout(),
            .ltout(\c0.n17566_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_1066_LC_14_28_6 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_1066_LC_14_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_1066_LC_14_28_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_1066_LC_14_28_6  (
            .in0(N__44512),
            .in1(N__48591),
            .in2(N__43277),
            .in3(N__43270),
            .lcout(\c0.n9195 ),
            .ltout(\c0.n9195_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1070_LC_14_28_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1070_LC_14_28_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1070_LC_14_28_7 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_1070_LC_14_28_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43235),
            .in3(N__43232),
            .lcout(\c0.n17608 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15806_4_lut_LC_14_29_0 .C_ON=1'b0;
    defparam \c0.i15806_4_lut_LC_14_29_0 .SEQ_MODE=4'b0000;
    defparam \c0.i15806_4_lut_LC_14_29_0 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \c0.i15806_4_lut_LC_14_29_0  (
            .in0(N__48155),
            .in1(N__43427),
            .in2(N__43190),
            .in3(N__47983),
            .lcout(\c0.n18015 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i8_3_lut_LC_14_29_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i8_3_lut_LC_14_29_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i8_3_lut_LC_14_29_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_0_i8_3_lut_LC_14_29_1  (
            .in0(N__43439),
            .in1(N__47833),
            .in2(_gnd_net_),
            .in3(N__48418),
            .lcout(\c0.n8_adj_2516 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1073_LC_14_29_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1073_LC_14_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1073_LC_14_29_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1073_LC_14_29_2  (
            .in0(_gnd_net_),
            .in1(N__49633),
            .in2(_gnd_net_),
            .in3(N__43528),
            .lcout(\c0.n17668 ),
            .ltout(\c0.n17668_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_3_lut_LC_14_29_3 .C_ON=1'b0;
    defparam \c0.i3_3_lut_LC_14_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_3_lut_LC_14_29_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i3_3_lut_LC_14_29_3  (
            .in0(N__43499),
            .in1(_gnd_net_),
            .in2(N__43493),
            .in3(N__43486),
            .lcout(),
            .ltout(\c0.n8_adj_2511_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_10__0__3517_LC_14_29_4 .C_ON=1'b0;
    defparam \c0.data_out_10__0__3517_LC_14_29_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_10__0__3517_LC_14_29_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_10__0__3517_LC_14_29_4  (
            .in0(N__46112),
            .in1(N__47533),
            .in2(N__43475),
            .in3(N__43472),
            .lcout(\c0.data_out_10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50420),
            .ce(N__46035),
            .sr(_gnd_net_));
    defparam \c0.data_out_9__0__3525_LC_14_29_5 .C_ON=1'b0;
    defparam \c0.data_out_9__0__3525_LC_14_29_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_9__0__3525_LC_14_29_5 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \c0.data_out_9__0__3525_LC_14_29_5  (
            .in0(N__47769),
            .in1(N__44419),
            .in2(_gnd_net_),
            .in3(N__43465),
            .lcout(\c0.data_out_9_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50420),
            .ce(N__46035),
            .sr(_gnd_net_));
    defparam \c0.i15843_2_lut_LC_14_29_6 .C_ON=1'b0;
    defparam \c0.i15843_2_lut_LC_14_29_6 .SEQ_MODE=4'b0000;
    defparam \c0.i15843_2_lut_LC_14_29_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \c0.i15843_2_lut_LC_14_29_6  (
            .in0(N__48419),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43433),
            .lcout(\c0.n18016 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1056_LC_14_30_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1056_LC_14_30_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1056_LC_14_30_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1056_LC_14_30_0  (
            .in0(N__49872),
            .in1(N__43584),
            .in2(N__44272),
            .in3(N__43655),
            .lcout(\c0.data_out_6__5__N_752 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1097_LC_14_30_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1097_LC_14_30_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1097_LC_14_30_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1097_LC_14_30_1  (
            .in0(_gnd_net_),
            .in1(N__47703),
            .in2(_gnd_net_),
            .in3(N__46447),
            .lcout(),
            .ltout(\c0.n4_adj_2543_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.mux_754_i1_4_lut_LC_14_30_2 .C_ON=1'b0;
    defparam \c0.mux_754_i1_4_lut_LC_14_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.mux_754_i1_4_lut_LC_14_30_2 .LUT_INIT=16'b1010101000111100;
    LogicCell40 \c0.mux_754_i1_4_lut_LC_14_30_2  (
            .in0(N__46255),
            .in1(N__43420),
            .in2(N__43361),
            .in3(N__49414),
            .lcout(),
            .ltout(\c0.n9656_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__5__3544_LC_14_30_3 .C_ON=1'b0;
    defparam \c0.data_out_6__5__3544_LC_14_30_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__5__3544_LC_14_30_3 .LUT_INIT=16'b1000101100000011;
    LogicCell40 \c0.data_out_6__5__3544_LC_14_30_3  (
            .in0(N__43889),
            .in1(N__46902),
            .in2(N__43868),
            .in3(N__47410),
            .lcout(\c0.data_out_6_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50425),
            .ce(N__46547),
            .sr(_gnd_net_));
    defparam \c0.mux_858_i1_4_lut_LC_14_30_4 .C_ON=1'b0;
    defparam \c0.mux_858_i1_4_lut_LC_14_30_4 .SEQ_MODE=4'b0000;
    defparam \c0.mux_858_i1_4_lut_LC_14_30_4 .LUT_INIT=16'b1100110010100101;
    LogicCell40 \c0.mux_858_i1_4_lut_LC_14_30_4  (
            .in0(N__43661),
            .in1(N__43825),
            .in2(N__49487),
            .in3(N__49415),
            .lcout(),
            .ltout(\c0.n2251_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__1__3548_LC_14_30_5 .C_ON=1'b0;
    defparam \c0.data_out_6__1__3548_LC_14_30_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__1__3548_LC_14_30_5 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \c0.data_out_6__1__3548_LC_14_30_5  (
            .in0(N__43865),
            .in1(N__46901),
            .in2(N__43841),
            .in3(N__47409),
            .lcout(\c0.data_out_6_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50425),
            .ce(N__46547),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_1065_LC_14_30_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_1065_LC_14_30_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_1065_LC_14_30_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_1065_LC_14_30_6  (
            .in0(_gnd_net_),
            .in1(N__44388),
            .in2(_gnd_net_),
            .in3(N__46275),
            .lcout(\c0.n17510 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_5__1__3556_LC_14_30_7 .C_ON=1'b0;
    defparam \c0.data_out_5__1__3556_LC_14_30_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_5__1__3556_LC_14_30_7 .LUT_INIT=16'b1100110011111010;
    LogicCell40 \c0.data_out_5__1__3556_LC_14_30_7  (
            .in0(N__49416),
            .in1(N__43838),
            .in2(N__43829),
            .in3(N__46903),
            .lcout(\c0.data_out_5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50425),
            .ce(N__46547),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_892_LC_14_31_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_892_LC_14_31_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_892_LC_14_31_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_892_LC_14_31_1  (
            .in0(N__43797),
            .in1(N__47768),
            .in2(N__43771),
            .in3(N__43947),
            .lcout(\c0.n8767 ),
            .ltout(\c0.n8767_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_836_LC_14_31_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_836_LC_14_31_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_836_LC_14_31_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \c0.i1_2_lut_adj_836_LC_14_31_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43721),
            .in3(N__49868),
            .lcout(\c0.n17457 ),
            .ltout(\c0.n17457_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_LC_14_31_3 .C_ON=1'b0;
    defparam \c0.i1_4_lut_LC_14_31_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_LC_14_31_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_4_lut_LC_14_31_3  (
            .in0(N__43718),
            .in1(N__43709),
            .in2(N__43682),
            .in3(N__43679),
            .lcout(\c0.n17415 ),
            .ltout(\c0.n17415_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_999_LC_14_31_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_999_LC_14_31_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_999_LC_14_31_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_999_LC_14_31_4  (
            .in0(N__43646),
            .in1(N__44264),
            .in2(N__43592),
            .in3(N__43580),
            .lcout(\c0.n17659 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__1__3540_LC_14_31_5 .C_ON=1'b0;
    defparam \c0.data_out_7__1__3540_LC_14_31_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__1__3540_LC_14_31_5 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \c0.data_out_7__1__3540_LC_14_31_5  (
            .in0(N__49163),
            .in1(N__46786),
            .in2(N__44219),
            .in3(N__47411),
            .lcout(\c0.data_out_7_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50428),
            .ce(N__44186),
            .sr(_gnd_net_));
    defparam \c0.data_out_3__0__3573_LC_14_32_1 .C_ON=1'b0;
    defparam \c0.data_out_3__0__3573_LC_14_32_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_3__0__3573_LC_14_32_1 .LUT_INIT=16'b1101110010001100;
    LogicCell40 \c0.data_out_3__0__3573_LC_14_32_1  (
            .in0(N__47110),
            .in1(N__44124),
            .in2(N__47449),
            .in3(N__47476),
            .lcout(data_out_6__2__N_804),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50431),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1068_LC_14_32_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1068_LC_14_32_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1068_LC_14_32_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_1068_LC_14_32_7  (
            .in0(N__46378),
            .in1(N__44080),
            .in2(_gnd_net_),
            .in3(N__49744),
            .lcout(\c0.n17654 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15781_4_lut_LC_15_23_7 .C_ON=1'b0;
    defparam \c0.i15781_4_lut_LC_15_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.i15781_4_lut_LC_15_23_7 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \c0.i15781_4_lut_LC_15_23_7  (
            .in0(N__45875),
            .in1(N__48148),
            .in2(N__43961),
            .in3(N__47970),
            .lcout(\c0.n18061 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15694_2_lut_LC_15_25_0 .C_ON=1'b0;
    defparam \c0.i15694_2_lut_LC_15_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.i15694_2_lut_LC_15_25_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i15694_2_lut_LC_15_25_0  (
            .in0(_gnd_net_),
            .in1(N__44050),
            .in2(_gnd_net_),
            .in3(N__48430),
            .lcout(\c0.n17943 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i2_3_lut_LC_15_25_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i2_3_lut_LC_15_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i2_3_lut_LC_15_25_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_7_i2_3_lut_LC_15_25_5  (
            .in0(N__48431),
            .in1(N__46440),
            .in2(_gnd_net_),
            .in3(N__44015),
            .lcout(\c0.n2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15746_2_lut_LC_15_25_6 .C_ON=1'b0;
    defparam \c0.i15746_2_lut_LC_15_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.i15746_2_lut_LC_15_25_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.i15746_2_lut_LC_15_25_6  (
            .in0(_gnd_net_),
            .in1(N__45758),
            .in2(_gnd_net_),
            .in3(N__48432),
            .lcout(\c0.n18060 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15784_2_lut_LC_15_26_0 .C_ON=1'b0;
    defparam \c0.i15784_2_lut_LC_15_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.i15784_2_lut_LC_15_26_0 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \c0.i15784_2_lut_LC_15_26_0  (
            .in0(N__43948),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48428),
            .lcout(\c0.n18091 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15791_4_lut_LC_15_26_1 .C_ON=1'b0;
    defparam \c0.i15791_4_lut_LC_15_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.i15791_4_lut_LC_15_26_1 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \c0.i15791_4_lut_LC_15_26_1  (
            .in0(N__46235),
            .in1(N__48151),
            .in2(N__45857),
            .in3(N__47968),
            .lcout(),
            .ltout(\c0.n18065_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11411_4_lut_LC_15_26_2 .C_ON=1'b0;
    defparam \c0.i11411_4_lut_LC_15_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.i11411_4_lut_LC_15_26_2 .LUT_INIT=16'b0101000001000100;
    LogicCell40 \c0.i11411_4_lut_LC_15_26_2  (
            .in0(N__48840),
            .in1(N__44279),
            .in2(N__44342),
            .in3(N__48736),
            .lcout(tx_data_5_N_keep),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_1029_LC_15_26_3 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_1029_LC_15_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_1029_LC_15_26_3 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \c0.i1_4_lut_adj_1029_LC_15_26_3  (
            .in0(N__48737),
            .in1(N__44225),
            .in2(N__44330),
            .in3(N__48839),
            .lcout(tx_data_1_N_keep),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i5_3_lut_LC_15_26_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i5_3_lut_LC_15_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i5_3_lut_LC_15_26_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_5_i5_3_lut_LC_15_26_4  (
            .in0(N__45596),
            .in1(N__46280),
            .in2(_gnd_net_),
            .in3(N__48427),
            .lcout(),
            .ltout(\c0.n5_adj_2481_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15955_LC_15_26_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15955_LC_15_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15955_LC_15_26_5 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter_1__bdd_4_lut_15955_LC_15_26_5  (
            .in0(N__44312),
            .in1(N__48149),
            .in2(N__44303),
            .in3(N__47967),
            .lcout(),
            .ltout(\c0.n18402_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18402_bdd_4_lut_LC_15_26_6 .C_ON=1'b0;
    defparam \c0.n18402_bdd_4_lut_LC_15_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.n18402_bdd_4_lut_LC_15_26_6 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n18402_bdd_4_lut_LC_15_26_6  (
            .in0(N__48150),
            .in1(N__44300),
            .in2(N__44294),
            .in3(N__44291),
            .lcout(\c0.n18405 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i59_3_lut_LC_15_27_0 .C_ON=1'b0;
    defparam \c0.i59_3_lut_LC_15_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.i59_3_lut_LC_15_27_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.i59_3_lut_LC_15_27_0  (
            .in0(N__46309),
            .in1(N__44395),
            .in2(_gnd_net_),
            .in3(N__48464),
            .lcout(),
            .ltout(\c0.n45_adj_2518_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i60_4_lut_LC_15_27_1 .C_ON=1'b0;
    defparam \c0.i60_4_lut_LC_15_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.i60_4_lut_LC_15_27_1 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \c0.i60_4_lut_LC_15_27_1  (
            .in0(N__48466),
            .in1(N__44273),
            .in2(N__44240),
            .in3(N__47972),
            .lcout(),
            .ltout(\c0.n46_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i58_4_lut_LC_15_27_2 .C_ON=1'b0;
    defparam \c0.i58_4_lut_LC_15_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.i58_4_lut_LC_15_27_2 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \c0.i58_4_lut_LC_15_27_2  (
            .in0(N__47973),
            .in1(N__44237),
            .in2(N__44228),
            .in3(N__48136),
            .lcout(\c0.n44_adj_2524 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_840_LC_15_27_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_840_LC_15_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_840_LC_15_27_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_840_LC_15_27_4  (
            .in0(_gnd_net_),
            .in1(N__47704),
            .in2(_gnd_net_),
            .in3(N__47636),
            .lcout(\c0.n8777 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15797_2_lut_LC_15_27_5 .C_ON=1'b0;
    defparam \c0.i15797_2_lut_LC_15_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.i15797_2_lut_LC_15_27_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \c0.i15797_2_lut_LC_15_27_5  (
            .in0(N__48465),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45542),
            .lcout(),
            .ltout(\c0.n18069_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15799_4_lut_LC_15_27_6 .C_ON=1'b0;
    defparam \c0.i15799_4_lut_LC_15_27_6 .SEQ_MODE=4'b0000;
    defparam \c0.i15799_4_lut_LC_15_27_6 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \c0.i15799_4_lut_LC_15_27_6  (
            .in0(N__47971),
            .in1(N__45533),
            .in2(N__45527),
            .in3(N__48135),
            .lcout(\c0.n18070 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0___i111_LC_15_27_7 .C_ON=1'b0;
    defparam \c0.data_in_0___i111_LC_15_27_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0___i111_LC_15_27_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0___i111_LC_15_27_7  (
            .in0(N__44944),
            .in1(N__44533),
            .in2(_gnd_net_),
            .in3(N__44561),
            .lcout(data_in_13_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50416),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_9__1__3524_LC_15_28_0 .C_ON=1'b0;
    defparam \c0.data_out_9__1__3524_LC_15_28_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_9__1__3524_LC_15_28_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_9__1__3524_LC_15_28_0  (
            .in0(N__49549),
            .in1(N__44522),
            .in2(N__47783),
            .in3(N__44513),
            .lcout(\c0.data_out_9_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50421),
            .ce(N__46015),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_1_i8_3_lut_LC_15_28_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_1_i8_3_lut_LC_15_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_1_i8_3_lut_LC_15_28_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_1_i8_3_lut_LC_15_28_1  (
            .in0(N__44495),
            .in1(N__44488),
            .in2(_gnd_net_),
            .in3(N__48467),
            .lcout(\c0.n8_adj_2519 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i8_3_lut_LC_15_28_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i8_3_lut_LC_15_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i8_3_lut_LC_15_28_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_4_i8_3_lut_LC_15_28_3  (
            .in0(N__44402),
            .in1(N__49616),
            .in2(_gnd_net_),
            .in3(N__48468),
            .lcout(\c0.n8_adj_2535 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_9__4__3521_LC_15_28_4 .C_ON=1'b0;
    defparam \c0.data_out_9__4__3521_LC_15_28_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_9__4__3521_LC_15_28_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_9__4__3521_LC_15_28_4  (
            .in0(N__45913),
            .in1(N__44435),
            .in2(N__44423),
            .in3(N__45838),
            .lcout(\c0.data_out_9_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50421),
            .ce(N__46015),
            .sr(_gnd_net_));
    defparam \c0.data_out_10__5__3512_LC_15_28_6 .C_ON=1'b0;
    defparam \c0.data_out_10__5__3512_LC_15_28_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_10__5__3512_LC_15_28_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_10__5__3512_LC_15_28_6  (
            .in0(N__47779),
            .in1(N__44396),
            .in2(N__44375),
            .in3(N__44354),
            .lcout(\c0.data_out_10_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50421),
            .ce(N__46015),
            .sr(_gnd_net_));
    defparam \c0.i15788_2_lut_LC_15_28_7 .C_ON=1'b0;
    defparam \c0.i15788_2_lut_LC_15_28_7 .SEQ_MODE=4'b0000;
    defparam \c0.i15788_2_lut_LC_15_28_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.i15788_2_lut_LC_15_28_7  (
            .in0(_gnd_net_),
            .in1(N__45863),
            .in2(_gnd_net_),
            .in3(N__48469),
            .lcout(\c0.n18064 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_3_lut_4_lut_LC_15_29_1 .C_ON=1'b0;
    defparam \c0.i3_3_lut_4_lut_LC_15_29_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_3_lut_4_lut_LC_15_29_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_3_lut_4_lut_LC_15_29_1  (
            .in0(N__45599),
            .in1(N__45845),
            .in2(N__45839),
            .in3(N__45657),
            .lcout(),
            .ltout(\c0.n8_adj_2528_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_10__1__3516_LC_15_29_2 .C_ON=1'b0;
    defparam \c0.data_out_10__1__3516_LC_15_29_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_10__1__3516_LC_15_29_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_10__1__3516_LC_15_29_2  (
            .in0(N__49476),
            .in1(N__49505),
            .in2(N__45803),
            .in3(N__46198),
            .lcout(\c0.data_out_10_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50426),
            .ce(N__46036),
            .sr(_gnd_net_));
    defparam \c0.data_out_10__7__3510_LC_15_29_3 .C_ON=1'b0;
    defparam \c0.data_out_10__7__3510_LC_15_29_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_10__7__3510_LC_15_29_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_out_10__7__3510_LC_15_29_3  (
            .in0(N__45557),
            .in1(N__45794),
            .in2(_gnd_net_),
            .in3(N__45778),
            .lcout(\c0.data_out_10_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50426),
            .ce(N__46036),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_863_LC_15_29_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_863_LC_15_29_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_863_LC_15_29_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_863_LC_15_29_4  (
            .in0(N__49783),
            .in1(N__45745),
            .in2(_gnd_net_),
            .in3(N__45721),
            .lcout(\c0.n17635 ),
            .ltout(\c0.n17635_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15674_3_lut_LC_15_29_5 .C_ON=1'b0;
    defparam \c0.i15674_3_lut_LC_15_29_5 .SEQ_MODE=4'b0000;
    defparam \c0.i15674_3_lut_LC_15_29_5 .LUT_INIT=16'b1100001100000000;
    LogicCell40 \c0.i15674_3_lut_LC_15_29_5  (
            .in0(_gnd_net_),
            .in1(N__45655),
            .in2(N__45680),
            .in3(N__49397),
            .lcout(\c0.n17922 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1032_LC_15_29_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1032_LC_15_29_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1032_LC_15_29_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1032_LC_15_29_6  (
            .in0(N__45656),
            .in1(N__45598),
            .in2(_gnd_net_),
            .in3(N__48208),
            .lcout(\c0.n17492 ),
            .ltout(\c0.n17492_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_10__3__3514_LC_15_29_7 .C_ON=1'b0;
    defparam \c0.data_out_10__3__3514_LC_15_29_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_10__3__3514_LC_15_29_7 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_10__3__3514_LC_15_29_7  (
            .in0(N__46286),
            .in1(N__45551),
            .in2(N__45545),
            .in3(N__46364),
            .lcout(\c0.data_out_10_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50426),
            .ce(N__46036),
            .sr(_gnd_net_));
    defparam \c0.data_out_9__6__3519_LC_15_30_0 .C_ON=1'b0;
    defparam \c0.data_out_9__6__3519_LC_15_30_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_9__6__3519_LC_15_30_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_9__6__3519_LC_15_30_0  (
            .in0(N__46183),
            .in1(N__46367),
            .in2(N__46328),
            .in3(N__49708),
            .lcout(\c0.data_out_9_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50429),
            .ce(N__46037),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i8_3_lut_LC_15_30_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i8_3_lut_LC_15_30_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i8_3_lut_LC_15_30_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_6_i8_3_lut_LC_15_30_1  (
            .in0(N__46316),
            .in1(N__46150),
            .in2(_gnd_net_),
            .in3(N__48458),
            .lcout(\c0.n8_adj_2539 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_997_LC_15_30_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_997_LC_15_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_997_LC_15_30_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_997_LC_15_30_2  (
            .in0(N__45912),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46302),
            .lcout(\c0.n17454 ),
            .ltout(\c0.n17454_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_9__5__3520_LC_15_30_3 .C_ON=1'b0;
    defparam \c0.data_out_9__5__3520_LC_15_30_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_9__5__3520_LC_15_30_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_9__5__3520_LC_15_30_3  (
            .in0(N__46279),
            .in1(N__46256),
            .in2(N__46244),
            .in3(N__49550),
            .lcout(\c0.data_out_9_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50429),
            .ce(N__46037),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i8_3_lut_LC_15_30_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i8_3_lut_LC_15_30_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i8_3_lut_LC_15_30_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_5_i8_3_lut_LC_15_30_4  (
            .in0(N__48459),
            .in1(N__46241),
            .in2(_gnd_net_),
            .in3(N__49707),
            .lcout(\c0.n8_adj_2537 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_949_LC_15_30_5 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_949_LC_15_30_5 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_949_LC_15_30_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_949_LC_15_30_5  (
            .in0(N__46223),
            .in1(N__46199),
            .in2(N__46184),
            .in3(N__46163),
            .lcout(),
            .ltout(\c0.n12_adj_2482_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_9__7__3518_LC_15_30_6 .C_ON=1'b0;
    defparam \c0.data_out_9__7__3518_LC_15_30_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_9__7__3518_LC_15_30_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_9__7__3518_LC_15_30_6  (
            .in0(N__46151),
            .in1(N__46105),
            .in2(N__46091),
            .in3(N__46088),
            .lcout(\c0.data_out_9_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50429),
            .ce(N__46037),
            .sr(_gnd_net_));
    defparam \c0.i10536_3_lut_LC_15_30_7 .C_ON=1'b0;
    defparam \c0.i10536_3_lut_LC_15_30_7 .SEQ_MODE=4'b0000;
    defparam \c0.i10536_3_lut_LC_15_30_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.i10536_3_lut_LC_15_30_7  (
            .in0(N__45920),
            .in1(N__45911),
            .in2(_gnd_net_),
            .in3(N__48457),
            .lcout(\c0.n8_adj_2538 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i1_3_lut_LC_15_31_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i1_3_lut_LC_15_31_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i1_3_lut_LC_15_31_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_6_i1_3_lut_LC_15_31_0  (
            .in0(N__46978),
            .in1(N__47770),
            .in2(_gnd_net_),
            .in3(N__48473),
            .lcout(\c0.n1_adj_2484 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_1124_LC_15_31_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_1124_LC_15_31_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_1124_LC_15_31_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_1124_LC_15_31_1  (
            .in0(N__47695),
            .in1(N__47640),
            .in2(_gnd_net_),
            .in3(N__47578),
            .lcout(\c0.n8926 ),
            .ltout(\c0.n8926_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_1109_LC_15_31_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_1109_LC_15_31_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_1109_LC_15_31_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i2_3_lut_adj_1109_LC_15_31_2  (
            .in0(_gnd_net_),
            .in1(N__47507),
            .in2(N__47501),
            .in3(N__46976),
            .lcout(\c0.n17438 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.mux_1207_i1_3_lut_LC_15_31_3 .C_ON=1'b0;
    defparam \c0.mux_1207_i1_3_lut_LC_15_31_3 .SEQ_MODE=4'b0000;
    defparam \c0.mux_1207_i1_3_lut_LC_15_31_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.mux_1207_i1_3_lut_LC_15_31_3  (
            .in0(N__49384),
            .in1(N__46800),
            .in2(_gnd_net_),
            .in3(N__47412),
            .lcout(n2720),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_1__6__3583_LC_15_31_4 .C_ON=1'b0;
    defparam \c0.data_out_1__6__3583_LC_15_31_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_1__6__3583_LC_15_31_4 .LUT_INIT=16'b1100111011000100;
    LogicCell40 \c0.data_out_1__6__3583_LC_15_31_4  (
            .in0(N__47413),
            .in1(N__46977),
            .in2(N__47134),
            .in3(N__46804),
            .lcout(data_out_1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50432),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_LC_15_31_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_LC_15_31_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_LC_15_31_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_LC_15_31_5  (
            .in0(N__46955),
            .in1(N__48502),
            .in2(_gnd_net_),
            .in3(N__46451),
            .lcout(\c0.data_out_6__3__N_781 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_3__6__3567_LC_15_31_6 .C_ON=1'b0;
    defparam \c0.data_out_3__6__3567_LC_15_31_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_3__6__3567_LC_15_31_6 .LUT_INIT=16'b0000110010101010;
    LogicCell40 \c0.data_out_3__6__3567_LC_15_31_6  (
            .in0(N__48503),
            .in1(N__49385),
            .in2(N__46881),
            .in3(N__46531),
            .lcout(data_out_3_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50432),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__4__I_567_2_lut_LC_15_31_7 .C_ON=1'b0;
    defparam \c0.data_out_6__4__I_567_2_lut_LC_15_31_7 .SEQ_MODE=4'b0000;
    defparam \c0.data_out_6__4__I_567_2_lut_LC_15_31_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.data_out_6__4__I_567_2_lut_LC_15_31_7  (
            .in0(_gnd_net_),
            .in1(N__48501),
            .in2(_gnd_net_),
            .in3(N__46450),
            .lcout(\c0.data_out_6__4__N_765 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15965_LC_16_27_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15965_LC_16_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15965_LC_16_27_0 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter_1__bdd_4_lut_15965_LC_16_27_0  (
            .in0(N__48533),
            .in1(N__48158),
            .in2(N__48182),
            .in3(N__47987),
            .lcout(),
            .ltout(\c0.n18414_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18414_bdd_4_lut_LC_16_27_1 .C_ON=1'b0;
    defparam \c0.n18414_bdd_4_lut_LC_16_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.n18414_bdd_4_lut_LC_16_27_1 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n18414_bdd_4_lut_LC_16_27_1  (
            .in0(N__48159),
            .in1(N__48860),
            .in2(N__48848),
            .in3(N__48479),
            .lcout(),
            .ltout(\c0.n18417_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11407_4_lut_LC_16_27_2 .C_ON=1'b0;
    defparam \c0.i11407_4_lut_LC_16_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.i11407_4_lut_LC_16_27_2 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \c0.i11407_4_lut_LC_16_27_2  (
            .in0(N__48838),
            .in1(N__47846),
            .in2(N__48764),
            .in3(N__48760),
            .lcout(),
            .ltout(tx_data_6_N_keep_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i6_LC_16_27_3 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i6_LC_16_27_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i6_LC_16_27_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \c0.tx.r_Tx_Data_i6_LC_16_27_3  (
            .in0(N__48682),
            .in1(_gnd_net_),
            .in2(N__48617),
            .in3(N__48607),
            .lcout(r_Tx_Data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50422),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15698_2_lut_LC_16_27_4 .C_ON=1'b0;
    defparam \c0.i15698_2_lut_LC_16_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.i15698_2_lut_LC_16_27_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i15698_2_lut_LC_16_27_4  (
            .in0(_gnd_net_),
            .in1(N__48593),
            .in2(_gnd_net_),
            .in3(N__48461),
            .lcout(\c0.n17949 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15720_2_lut_LC_16_27_5 .C_ON=1'b0;
    defparam \c0.i15720_2_lut_LC_16_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.i15720_2_lut_LC_16_27_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i15720_2_lut_LC_16_27_5  (
            .in0(N__48463),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48522),
            .lcout(\c0.n18090 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i5_3_lut_LC_16_27_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i5_3_lut_LC_16_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i5_3_lut_LC_16_27_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_6_i5_3_lut_LC_16_27_7  (
            .in0(N__48462),
            .in1(N__49663),
            .in2(_gnd_net_),
            .in3(N__48209),
            .lcout(\c0.n5_adj_2444 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15787_4_lut_LC_16_28_0 .C_ON=1'b0;
    defparam \c0.i15787_4_lut_LC_16_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.i15787_4_lut_LC_16_28_0 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \c0.i15787_4_lut_LC_16_28_0  (
            .in0(N__48173),
            .in1(N__48157),
            .in2(N__47999),
            .in3(N__47986),
            .lcout(\c0.n18063 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_888_LC_16_28_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_888_LC_16_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_888_LC_16_28_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_888_LC_16_28_3  (
            .in0(_gnd_net_),
            .in1(N__47840),
            .in2(_gnd_net_),
            .in3(N__47807),
            .lcout(\c0.n17638 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2271__i0_LC_16_29_0.C_ON=1'b1;
    defparam blink_counter_2271__i0_LC_16_29_0.SEQ_MODE=4'b1000;
    defparam blink_counter_2271__i0_LC_16_29_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2271__i0_LC_16_29_0 (
            .in0(_gnd_net_),
            .in1(N__48932),
            .in2(_gnd_net_),
            .in3(N__48926),
            .lcout(n26),
            .ltout(),
            .carryin(bfn_16_29_0_),
            .carryout(n16380),
            .clk(N__50430),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2271__i1_LC_16_29_1.C_ON=1'b1;
    defparam blink_counter_2271__i1_LC_16_29_1.SEQ_MODE=4'b1000;
    defparam blink_counter_2271__i1_LC_16_29_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2271__i1_LC_16_29_1 (
            .in0(_gnd_net_),
            .in1(N__48923),
            .in2(_gnd_net_),
            .in3(N__48917),
            .lcout(n25),
            .ltout(),
            .carryin(n16380),
            .carryout(n16381),
            .clk(N__50430),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2271__i2_LC_16_29_2.C_ON=1'b1;
    defparam blink_counter_2271__i2_LC_16_29_2.SEQ_MODE=4'b1000;
    defparam blink_counter_2271__i2_LC_16_29_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2271__i2_LC_16_29_2 (
            .in0(_gnd_net_),
            .in1(N__48914),
            .in2(_gnd_net_),
            .in3(N__48908),
            .lcout(n24),
            .ltout(),
            .carryin(n16381),
            .carryout(n16382),
            .clk(N__50430),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2271__i3_LC_16_29_3.C_ON=1'b1;
    defparam blink_counter_2271__i3_LC_16_29_3.SEQ_MODE=4'b1000;
    defparam blink_counter_2271__i3_LC_16_29_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2271__i3_LC_16_29_3 (
            .in0(_gnd_net_),
            .in1(N__48905),
            .in2(_gnd_net_),
            .in3(N__48899),
            .lcout(n23),
            .ltout(),
            .carryin(n16382),
            .carryout(n16383),
            .clk(N__50430),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2271__i4_LC_16_29_4.C_ON=1'b1;
    defparam blink_counter_2271__i4_LC_16_29_4.SEQ_MODE=4'b1000;
    defparam blink_counter_2271__i4_LC_16_29_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2271__i4_LC_16_29_4 (
            .in0(_gnd_net_),
            .in1(N__48896),
            .in2(_gnd_net_),
            .in3(N__48890),
            .lcout(n22_adj_2655),
            .ltout(),
            .carryin(n16383),
            .carryout(n16384),
            .clk(N__50430),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2271__i5_LC_16_29_5.C_ON=1'b1;
    defparam blink_counter_2271__i5_LC_16_29_5.SEQ_MODE=4'b1000;
    defparam blink_counter_2271__i5_LC_16_29_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2271__i5_LC_16_29_5 (
            .in0(_gnd_net_),
            .in1(N__48887),
            .in2(_gnd_net_),
            .in3(N__48881),
            .lcout(n21),
            .ltout(),
            .carryin(n16384),
            .carryout(n16385),
            .clk(N__50430),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2271__i6_LC_16_29_6.C_ON=1'b1;
    defparam blink_counter_2271__i6_LC_16_29_6.SEQ_MODE=4'b1000;
    defparam blink_counter_2271__i6_LC_16_29_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2271__i6_LC_16_29_6 (
            .in0(_gnd_net_),
            .in1(N__48878),
            .in2(_gnd_net_),
            .in3(N__48872),
            .lcout(n20),
            .ltout(),
            .carryin(n16385),
            .carryout(n16386),
            .clk(N__50430),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2271__i7_LC_16_29_7.C_ON=1'b1;
    defparam blink_counter_2271__i7_LC_16_29_7.SEQ_MODE=4'b1000;
    defparam blink_counter_2271__i7_LC_16_29_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2271__i7_LC_16_29_7 (
            .in0(_gnd_net_),
            .in1(N__48869),
            .in2(_gnd_net_),
            .in3(N__48863),
            .lcout(n19),
            .ltout(),
            .carryin(n16386),
            .carryout(n16387),
            .clk(N__50430),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2271__i8_LC_16_30_0.C_ON=1'b1;
    defparam blink_counter_2271__i8_LC_16_30_0.SEQ_MODE=4'b1000;
    defparam blink_counter_2271__i8_LC_16_30_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2271__i8_LC_16_30_0 (
            .in0(_gnd_net_),
            .in1(N__49010),
            .in2(_gnd_net_),
            .in3(N__49004),
            .lcout(n18),
            .ltout(),
            .carryin(bfn_16_30_0_),
            .carryout(n16388),
            .clk(N__50433),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2271__i9_LC_16_30_1.C_ON=1'b1;
    defparam blink_counter_2271__i9_LC_16_30_1.SEQ_MODE=4'b1000;
    defparam blink_counter_2271__i9_LC_16_30_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2271__i9_LC_16_30_1 (
            .in0(_gnd_net_),
            .in1(N__49001),
            .in2(_gnd_net_),
            .in3(N__48995),
            .lcout(n17),
            .ltout(),
            .carryin(n16388),
            .carryout(n16389),
            .clk(N__50433),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2271__i10_LC_16_30_2.C_ON=1'b1;
    defparam blink_counter_2271__i10_LC_16_30_2.SEQ_MODE=4'b1000;
    defparam blink_counter_2271__i10_LC_16_30_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2271__i10_LC_16_30_2 (
            .in0(_gnd_net_),
            .in1(N__48992),
            .in2(_gnd_net_),
            .in3(N__48986),
            .lcout(n16),
            .ltout(),
            .carryin(n16389),
            .carryout(n16390),
            .clk(N__50433),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2271__i11_LC_16_30_3.C_ON=1'b1;
    defparam blink_counter_2271__i11_LC_16_30_3.SEQ_MODE=4'b1000;
    defparam blink_counter_2271__i11_LC_16_30_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2271__i11_LC_16_30_3 (
            .in0(_gnd_net_),
            .in1(N__48983),
            .in2(_gnd_net_),
            .in3(N__48977),
            .lcout(n15),
            .ltout(),
            .carryin(n16390),
            .carryout(n16391),
            .clk(N__50433),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2271__i12_LC_16_30_4.C_ON=1'b1;
    defparam blink_counter_2271__i12_LC_16_30_4.SEQ_MODE=4'b1000;
    defparam blink_counter_2271__i12_LC_16_30_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2271__i12_LC_16_30_4 (
            .in0(_gnd_net_),
            .in1(N__48974),
            .in2(_gnd_net_),
            .in3(N__48968),
            .lcout(n14),
            .ltout(),
            .carryin(n16391),
            .carryout(n16392),
            .clk(N__50433),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2271__i13_LC_16_30_5.C_ON=1'b1;
    defparam blink_counter_2271__i13_LC_16_30_5.SEQ_MODE=4'b1000;
    defparam blink_counter_2271__i13_LC_16_30_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2271__i13_LC_16_30_5 (
            .in0(_gnd_net_),
            .in1(N__48965),
            .in2(_gnd_net_),
            .in3(N__48959),
            .lcout(n13),
            .ltout(),
            .carryin(n16392),
            .carryout(n16393),
            .clk(N__50433),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2271__i14_LC_16_30_6.C_ON=1'b1;
    defparam blink_counter_2271__i14_LC_16_30_6.SEQ_MODE=4'b1000;
    defparam blink_counter_2271__i14_LC_16_30_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2271__i14_LC_16_30_6 (
            .in0(_gnd_net_),
            .in1(N__48956),
            .in2(_gnd_net_),
            .in3(N__48950),
            .lcout(n12),
            .ltout(),
            .carryin(n16393),
            .carryout(n16394),
            .clk(N__50433),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2271__i15_LC_16_30_7.C_ON=1'b1;
    defparam blink_counter_2271__i15_LC_16_30_7.SEQ_MODE=4'b1000;
    defparam blink_counter_2271__i15_LC_16_30_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2271__i15_LC_16_30_7 (
            .in0(_gnd_net_),
            .in1(N__48947),
            .in2(_gnd_net_),
            .in3(N__48941),
            .lcout(n11),
            .ltout(),
            .carryin(n16394),
            .carryout(n16395),
            .clk(N__50433),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2271__i16_LC_16_31_0.C_ON=1'b1;
    defparam blink_counter_2271__i16_LC_16_31_0.SEQ_MODE=4'b1000;
    defparam blink_counter_2271__i16_LC_16_31_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2271__i16_LC_16_31_0 (
            .in0(_gnd_net_),
            .in1(N__48938),
            .in2(_gnd_net_),
            .in3(N__49151),
            .lcout(n10),
            .ltout(),
            .carryin(bfn_16_31_0_),
            .carryout(n16396),
            .clk(N__50434),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2271__i17_LC_16_31_1.C_ON=1'b1;
    defparam blink_counter_2271__i17_LC_16_31_1.SEQ_MODE=4'b1000;
    defparam blink_counter_2271__i17_LC_16_31_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2271__i17_LC_16_31_1 (
            .in0(_gnd_net_),
            .in1(N__49148),
            .in2(_gnd_net_),
            .in3(N__49142),
            .lcout(n9),
            .ltout(),
            .carryin(n16396),
            .carryout(n16397),
            .clk(N__50434),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2271__i18_LC_16_31_2.C_ON=1'b1;
    defparam blink_counter_2271__i18_LC_16_31_2.SEQ_MODE=4'b1000;
    defparam blink_counter_2271__i18_LC_16_31_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2271__i18_LC_16_31_2 (
            .in0(_gnd_net_),
            .in1(N__49139),
            .in2(_gnd_net_),
            .in3(N__49133),
            .lcout(n8_adj_2617),
            .ltout(),
            .carryin(n16397),
            .carryout(n16398),
            .clk(N__50434),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2271__i19_LC_16_31_3.C_ON=1'b1;
    defparam blink_counter_2271__i19_LC_16_31_3.SEQ_MODE=4'b1000;
    defparam blink_counter_2271__i19_LC_16_31_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2271__i19_LC_16_31_3 (
            .in0(_gnd_net_),
            .in1(N__49130),
            .in2(_gnd_net_),
            .in3(N__49124),
            .lcout(n7),
            .ltout(),
            .carryin(n16398),
            .carryout(n16399),
            .clk(N__50434),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2271__i20_LC_16_31_4.C_ON=1'b1;
    defparam blink_counter_2271__i20_LC_16_31_4.SEQ_MODE=4'b1000;
    defparam blink_counter_2271__i20_LC_16_31_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2271__i20_LC_16_31_4 (
            .in0(_gnd_net_),
            .in1(N__49121),
            .in2(_gnd_net_),
            .in3(N__49115),
            .lcout(n6),
            .ltout(),
            .carryin(n16399),
            .carryout(n16400),
            .clk(N__50434),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2271__i21_LC_16_31_5.C_ON=1'b1;
    defparam blink_counter_2271__i21_LC_16_31_5.SEQ_MODE=4'b1000;
    defparam blink_counter_2271__i21_LC_16_31_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2271__i21_LC_16_31_5 (
            .in0(_gnd_net_),
            .in1(N__49102),
            .in2(_gnd_net_),
            .in3(N__49091),
            .lcout(blink_counter_21),
            .ltout(),
            .carryin(n16400),
            .carryout(n16401),
            .clk(N__50434),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2271__i22_LC_16_31_6.C_ON=1'b1;
    defparam blink_counter_2271__i22_LC_16_31_6.SEQ_MODE=4'b1000;
    defparam blink_counter_2271__i22_LC_16_31_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2271__i22_LC_16_31_6 (
            .in0(_gnd_net_),
            .in1(N__49078),
            .in2(_gnd_net_),
            .in3(N__49067),
            .lcout(blink_counter_22),
            .ltout(),
            .carryin(n16401),
            .carryout(n16402),
            .clk(N__50434),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2271__i23_LC_16_31_7.C_ON=1'b1;
    defparam blink_counter_2271__i23_LC_16_31_7.SEQ_MODE=4'b1000;
    defparam blink_counter_2271__i23_LC_16_31_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2271__i23_LC_16_31_7 (
            .in0(_gnd_net_),
            .in1(N__49057),
            .in2(_gnd_net_),
            .in3(N__49046),
            .lcout(blink_counter_23),
            .ltout(),
            .carryin(n16402),
            .carryout(n16403),
            .clk(N__50434),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2271__i24_LC_16_32_0.C_ON=1'b1;
    defparam blink_counter_2271__i24_LC_16_32_0.SEQ_MODE=4'b1000;
    defparam blink_counter_2271__i24_LC_16_32_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2271__i24_LC_16_32_0 (
            .in0(_gnd_net_),
            .in1(N__49024),
            .in2(_gnd_net_),
            .in3(N__49013),
            .lcout(blink_counter_24),
            .ltout(),
            .carryin(bfn_16_32_0_),
            .carryout(n16404),
            .clk(N__50435),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2271__i25_LC_16_32_1.C_ON=1'b0;
    defparam blink_counter_2271__i25_LC_16_32_1.SEQ_MODE=4'b1000;
    defparam blink_counter_2271__i25_LC_16_32_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2271__i25_LC_16_32_1 (
            .in0(_gnd_net_),
            .in1(N__50446),
            .in2(_gnd_net_),
            .in3(N__50462),
            .lcout(blink_counter_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50435),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15672_4_lut_LC_16_32_3 .C_ON=1'b0;
    defparam \c0.i15672_4_lut_LC_16_32_3 .SEQ_MODE=4'b0000;
    defparam \c0.i15672_4_lut_LC_16_32_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i15672_4_lut_LC_16_32_3  (
            .in0(N__49873),
            .in1(N__49807),
            .in2(N__49793),
            .in3(N__49748),
            .lcout(\c0.n17976 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1054_LC_17_29_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1054_LC_17_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_1054_LC_17_29_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_1054_LC_17_29_2  (
            .in0(N__49610),
            .in1(N__49721),
            .in2(N__49709),
            .in3(N__49667),
            .lcout(\c0.n8922 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_929_LC_17_29_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_929_LC_17_29_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_929_LC_17_29_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_929_LC_17_29_5  (
            .in0(_gnd_net_),
            .in1(N__49611),
            .in2(_gnd_net_),
            .in3(N__49574),
            .lcout(\c0.n17620 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15663_4_lut_LC_18_29_0 .C_ON=1'b0;
    defparam \c0.i15663_4_lut_LC_18_29_0 .SEQ_MODE=4'b0000;
    defparam \c0.i15663_4_lut_LC_18_29_0 .LUT_INIT=16'b0110100100000000;
    LogicCell40 \c0.i15663_4_lut_LC_18_29_0  (
            .in0(N__49526),
            .in1(N__49504),
            .in2(N__49486),
            .in3(N__49436),
            .lcout(\c0.n17918 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // TinyFPGA_B
