// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 12 2017 08:25:46

// File Generated:     Sep 12 2019 19:45:28

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "TinyFPGA_B" view "INTERFACE"

module TinyFPGA_B (
    USBPU,
    PIN_9,
    PIN_8,
    PIN_7,
    PIN_6,
    PIN_5,
    PIN_4,
    PIN_3,
    PIN_24,
    PIN_23,
    PIN_22,
    PIN_21,
    PIN_20,
    PIN_2,
    PIN_19,
    PIN_18,
    PIN_17,
    PIN_16,
    PIN_15,
    PIN_14,
    PIN_13,
    PIN_12,
    PIN_11,
    PIN_10,
    PIN_1,
    LED,
    CLK);

    output USBPU;
    input PIN_9;
    input PIN_8;
    input PIN_7;
    input PIN_6;
    input PIN_5;
    input PIN_4;
    inout PIN_3;
    input PIN_24;
    input PIN_23;
    input PIN_22;
    input PIN_21;
    input PIN_20;
    inout PIN_2;
    input PIN_19;
    input PIN_18;
    input PIN_17;
    input PIN_16;
    input PIN_15;
    input PIN_14;
    input PIN_13;
    input PIN_12;
    input PIN_11;
    input PIN_10;
    inout PIN_1;
    output LED;
    input CLK;

    wire N__50887;
    wire N__50886;
    wire N__50885;
    wire N__50878;
    wire N__50877;
    wire N__50876;
    wire N__50869;
    wire N__50868;
    wire N__50867;
    wire N__50860;
    wire N__50859;
    wire N__50858;
    wire N__50851;
    wire N__50850;
    wire N__50849;
    wire N__50842;
    wire N__50841;
    wire N__50840;
    wire N__50823;
    wire N__50820;
    wire N__50819;
    wire N__50818;
    wire N__50817;
    wire N__50816;
    wire N__50813;
    wire N__50808;
    wire N__50805;
    wire N__50802;
    wire N__50799;
    wire N__50796;
    wire N__50793;
    wire N__50790;
    wire N__50781;
    wire N__50780;
    wire N__50777;
    wire N__50774;
    wire N__50773;
    wire N__50770;
    wire N__50767;
    wire N__50764;
    wire N__50763;
    wire N__50762;
    wire N__50755;
    wire N__50750;
    wire N__50745;
    wire N__50744;
    wire N__50743;
    wire N__50742;
    wire N__50741;
    wire N__50740;
    wire N__50737;
    wire N__50734;
    wire N__50733;
    wire N__50730;
    wire N__50727;
    wire N__50724;
    wire N__50723;
    wire N__50722;
    wire N__50721;
    wire N__50720;
    wire N__50719;
    wire N__50718;
    wire N__50717;
    wire N__50710;
    wire N__50707;
    wire N__50700;
    wire N__50699;
    wire N__50698;
    wire N__50695;
    wire N__50692;
    wire N__50689;
    wire N__50688;
    wire N__50685;
    wire N__50684;
    wire N__50681;
    wire N__50678;
    wire N__50677;
    wire N__50676;
    wire N__50673;
    wire N__50670;
    wire N__50667;
    wire N__50664;
    wire N__50657;
    wire N__50654;
    wire N__50649;
    wire N__50646;
    wire N__50643;
    wire N__50638;
    wire N__50631;
    wire N__50622;
    wire N__50617;
    wire N__50612;
    wire N__50607;
    wire N__50604;
    wire N__50601;
    wire N__50596;
    wire N__50589;
    wire N__50588;
    wire N__50587;
    wire N__50584;
    wire N__50583;
    wire N__50580;
    wire N__50577;
    wire N__50576;
    wire N__50575;
    wire N__50574;
    wire N__50571;
    wire N__50568;
    wire N__50567;
    wire N__50566;
    wire N__50563;
    wire N__50560;
    wire N__50557;
    wire N__50556;
    wire N__50555;
    wire N__50554;
    wire N__50553;
    wire N__50552;
    wire N__50549;
    wire N__50548;
    wire N__50547;
    wire N__50546;
    wire N__50543;
    wire N__50542;
    wire N__50541;
    wire N__50538;
    wire N__50537;
    wire N__50534;
    wire N__50533;
    wire N__50530;
    wire N__50529;
    wire N__50526;
    wire N__50521;
    wire N__50518;
    wire N__50511;
    wire N__50506;
    wire N__50505;
    wire N__50502;
    wire N__50499;
    wire N__50496;
    wire N__50493;
    wire N__50492;
    wire N__50491;
    wire N__50484;
    wire N__50481;
    wire N__50478;
    wire N__50475;
    wire N__50472;
    wire N__50471;
    wire N__50470;
    wire N__50467;
    wire N__50464;
    wire N__50457;
    wire N__50452;
    wire N__50449;
    wire N__50446;
    wire N__50443;
    wire N__50436;
    wire N__50433;
    wire N__50430;
    wire N__50427;
    wire N__50424;
    wire N__50419;
    wire N__50418;
    wire N__50415;
    wire N__50412;
    wire N__50411;
    wire N__50408;
    wire N__50405;
    wire N__50398;
    wire N__50391;
    wire N__50390;
    wire N__50387;
    wire N__50384;
    wire N__50377;
    wire N__50372;
    wire N__50369;
    wire N__50366;
    wire N__50357;
    wire N__50354;
    wire N__50337;
    wire N__50334;
    wire N__50333;
    wire N__50330;
    wire N__50329;
    wire N__50328;
    wire N__50325;
    wire N__50324;
    wire N__50323;
    wire N__50322;
    wire N__50321;
    wire N__50320;
    wire N__50319;
    wire N__50318;
    wire N__50317;
    wire N__50316;
    wire N__50315;
    wire N__50314;
    wire N__50311;
    wire N__50306;
    wire N__50301;
    wire N__50296;
    wire N__50293;
    wire N__50292;
    wire N__50291;
    wire N__50290;
    wire N__50287;
    wire N__50284;
    wire N__50281;
    wire N__50278;
    wire N__50277;
    wire N__50276;
    wire N__50275;
    wire N__50272;
    wire N__50271;
    wire N__50270;
    wire N__50267;
    wire N__50266;
    wire N__50263;
    wire N__50262;
    wire N__50261;
    wire N__50260;
    wire N__50259;
    wire N__50254;
    wire N__50249;
    wire N__50248;
    wire N__50245;
    wire N__50244;
    wire N__50241;
    wire N__50238;
    wire N__50237;
    wire N__50236;
    wire N__50233;
    wire N__50230;
    wire N__50227;
    wire N__50222;
    wire N__50215;
    wire N__50212;
    wire N__50207;
    wire N__50206;
    wire N__50205;
    wire N__50204;
    wire N__50201;
    wire N__50198;
    wire N__50195;
    wire N__50192;
    wire N__50187;
    wire N__50184;
    wire N__50179;
    wire N__50176;
    wire N__50173;
    wire N__50170;
    wire N__50165;
    wire N__50162;
    wire N__50159;
    wire N__50158;
    wire N__50157;
    wire N__50156;
    wire N__50155;
    wire N__50154;
    wire N__50153;
    wire N__50152;
    wire N__50151;
    wire N__50150;
    wire N__50147;
    wire N__50138;
    wire N__50137;
    wire N__50136;
    wire N__50135;
    wire N__50130;
    wire N__50125;
    wire N__50122;
    wire N__50119;
    wire N__50116;
    wire N__50111;
    wire N__50108;
    wire N__50105;
    wire N__50100;
    wire N__50097;
    wire N__50088;
    wire N__50081;
    wire N__50076;
    wire N__50073;
    wire N__50066;
    wire N__50061;
    wire N__50054;
    wire N__50047;
    wire N__50044;
    wire N__50033;
    wire N__50028;
    wire N__50007;
    wire N__50004;
    wire N__50003;
    wire N__50000;
    wire N__49997;
    wire N__49994;
    wire N__49989;
    wire N__49988;
    wire N__49985;
    wire N__49984;
    wire N__49981;
    wire N__49980;
    wire N__49979;
    wire N__49978;
    wire N__49977;
    wire N__49974;
    wire N__49971;
    wire N__49970;
    wire N__49967;
    wire N__49964;
    wire N__49963;
    wire N__49962;
    wire N__49959;
    wire N__49956;
    wire N__49953;
    wire N__49950;
    wire N__49947;
    wire N__49944;
    wire N__49939;
    wire N__49936;
    wire N__49935;
    wire N__49934;
    wire N__49931;
    wire N__49930;
    wire N__49929;
    wire N__49924;
    wire N__49921;
    wire N__49916;
    wire N__49913;
    wire N__49910;
    wire N__49907;
    wire N__49902;
    wire N__49897;
    wire N__49894;
    wire N__49889;
    wire N__49886;
    wire N__49881;
    wire N__49866;
    wire N__49865;
    wire N__49862;
    wire N__49859;
    wire N__49854;
    wire N__49851;
    wire N__49850;
    wire N__49849;
    wire N__49848;
    wire N__49847;
    wire N__49846;
    wire N__49845;
    wire N__49844;
    wire N__49843;
    wire N__49842;
    wire N__49841;
    wire N__49840;
    wire N__49839;
    wire N__49838;
    wire N__49837;
    wire N__49836;
    wire N__49835;
    wire N__49834;
    wire N__49833;
    wire N__49832;
    wire N__49831;
    wire N__49830;
    wire N__49829;
    wire N__49828;
    wire N__49827;
    wire N__49826;
    wire N__49825;
    wire N__49824;
    wire N__49823;
    wire N__49822;
    wire N__49821;
    wire N__49820;
    wire N__49819;
    wire N__49818;
    wire N__49817;
    wire N__49816;
    wire N__49815;
    wire N__49814;
    wire N__49813;
    wire N__49812;
    wire N__49811;
    wire N__49810;
    wire N__49809;
    wire N__49808;
    wire N__49807;
    wire N__49806;
    wire N__49805;
    wire N__49804;
    wire N__49803;
    wire N__49802;
    wire N__49801;
    wire N__49800;
    wire N__49799;
    wire N__49798;
    wire N__49797;
    wire N__49796;
    wire N__49795;
    wire N__49794;
    wire N__49793;
    wire N__49792;
    wire N__49791;
    wire N__49790;
    wire N__49789;
    wire N__49788;
    wire N__49787;
    wire N__49786;
    wire N__49785;
    wire N__49784;
    wire N__49783;
    wire N__49782;
    wire N__49781;
    wire N__49780;
    wire N__49779;
    wire N__49778;
    wire N__49777;
    wire N__49776;
    wire N__49775;
    wire N__49774;
    wire N__49773;
    wire N__49772;
    wire N__49771;
    wire N__49770;
    wire N__49769;
    wire N__49768;
    wire N__49767;
    wire N__49766;
    wire N__49765;
    wire N__49764;
    wire N__49763;
    wire N__49762;
    wire N__49761;
    wire N__49760;
    wire N__49759;
    wire N__49758;
    wire N__49757;
    wire N__49756;
    wire N__49755;
    wire N__49754;
    wire N__49753;
    wire N__49752;
    wire N__49751;
    wire N__49750;
    wire N__49749;
    wire N__49748;
    wire N__49747;
    wire N__49746;
    wire N__49745;
    wire N__49744;
    wire N__49743;
    wire N__49742;
    wire N__49741;
    wire N__49740;
    wire N__49739;
    wire N__49738;
    wire N__49737;
    wire N__49736;
    wire N__49735;
    wire N__49734;
    wire N__49733;
    wire N__49732;
    wire N__49731;
    wire N__49730;
    wire N__49729;
    wire N__49728;
    wire N__49727;
    wire N__49726;
    wire N__49725;
    wire N__49724;
    wire N__49723;
    wire N__49722;
    wire N__49721;
    wire N__49720;
    wire N__49719;
    wire N__49718;
    wire N__49717;
    wire N__49716;
    wire N__49715;
    wire N__49714;
    wire N__49713;
    wire N__49712;
    wire N__49711;
    wire N__49710;
    wire N__49709;
    wire N__49708;
    wire N__49707;
    wire N__49706;
    wire N__49705;
    wire N__49704;
    wire N__49703;
    wire N__49702;
    wire N__49701;
    wire N__49700;
    wire N__49699;
    wire N__49698;
    wire N__49697;
    wire N__49696;
    wire N__49695;
    wire N__49694;
    wire N__49693;
    wire N__49692;
    wire N__49691;
    wire N__49690;
    wire N__49689;
    wire N__49688;
    wire N__49687;
    wire N__49686;
    wire N__49685;
    wire N__49684;
    wire N__49683;
    wire N__49682;
    wire N__49681;
    wire N__49680;
    wire N__49679;
    wire N__49678;
    wire N__49677;
    wire N__49676;
    wire N__49675;
    wire N__49674;
    wire N__49673;
    wire N__49672;
    wire N__49671;
    wire N__49670;
    wire N__49669;
    wire N__49668;
    wire N__49667;
    wire N__49666;
    wire N__49665;
    wire N__49664;
    wire N__49663;
    wire N__49662;
    wire N__49661;
    wire N__49660;
    wire N__49659;
    wire N__49658;
    wire N__49657;
    wire N__49656;
    wire N__49655;
    wire N__49654;
    wire N__49653;
    wire N__49652;
    wire N__49651;
    wire N__49650;
    wire N__49649;
    wire N__49648;
    wire N__49647;
    wire N__49646;
    wire N__49645;
    wire N__49644;
    wire N__49643;
    wire N__49642;
    wire N__49641;
    wire N__49640;
    wire N__49639;
    wire N__49638;
    wire N__49637;
    wire N__49636;
    wire N__49635;
    wire N__49634;
    wire N__49633;
    wire N__49632;
    wire N__49631;
    wire N__49630;
    wire N__49629;
    wire N__49628;
    wire N__49627;
    wire N__49176;
    wire N__49173;
    wire N__49170;
    wire N__49169;
    wire N__49168;
    wire N__49165;
    wire N__49162;
    wire N__49161;
    wire N__49158;
    wire N__49155;
    wire N__49152;
    wire N__49151;
    wire N__49148;
    wire N__49147;
    wire N__49144;
    wire N__49141;
    wire N__49138;
    wire N__49135;
    wire N__49132;
    wire N__49129;
    wire N__49122;
    wire N__49113;
    wire N__49112;
    wire N__49111;
    wire N__49110;
    wire N__49109;
    wire N__49106;
    wire N__49103;
    wire N__49100;
    wire N__49099;
    wire N__49094;
    wire N__49091;
    wire N__49088;
    wire N__49085;
    wire N__49084;
    wire N__49081;
    wire N__49078;
    wire N__49075;
    wire N__49072;
    wire N__49069;
    wire N__49066;
    wire N__49065;
    wire N__49060;
    wire N__49051;
    wire N__49048;
    wire N__49041;
    wire N__49040;
    wire N__49037;
    wire N__49034;
    wire N__49033;
    wire N__49030;
    wire N__49025;
    wire N__49022;
    wire N__49019;
    wire N__49014;
    wire N__49013;
    wire N__49010;
    wire N__49007;
    wire N__49006;
    wire N__49005;
    wire N__49000;
    wire N__48997;
    wire N__48994;
    wire N__48991;
    wire N__48988;
    wire N__48981;
    wire N__48978;
    wire N__48975;
    wire N__48972;
    wire N__48971;
    wire N__48968;
    wire N__48965;
    wire N__48964;
    wire N__48963;
    wire N__48958;
    wire N__48953;
    wire N__48948;
    wire N__48945;
    wire N__48942;
    wire N__48939;
    wire N__48936;
    wire N__48933;
    wire N__48930;
    wire N__48927;
    wire N__48926;
    wire N__48925;
    wire N__48922;
    wire N__48919;
    wire N__48916;
    wire N__48913;
    wire N__48908;
    wire N__48903;
    wire N__48900;
    wire N__48897;
    wire N__48896;
    wire N__48893;
    wire N__48890;
    wire N__48885;
    wire N__48884;
    wire N__48883;
    wire N__48880;
    wire N__48877;
    wire N__48874;
    wire N__48871;
    wire N__48868;
    wire N__48865;
    wire N__48864;
    wire N__48861;
    wire N__48858;
    wire N__48855;
    wire N__48852;
    wire N__48849;
    wire N__48844;
    wire N__48841;
    wire N__48834;
    wire N__48831;
    wire N__48828;
    wire N__48827;
    wire N__48826;
    wire N__48825;
    wire N__48822;
    wire N__48819;
    wire N__48816;
    wire N__48815;
    wire N__48812;
    wire N__48805;
    wire N__48802;
    wire N__48795;
    wire N__48792;
    wire N__48791;
    wire N__48788;
    wire N__48785;
    wire N__48782;
    wire N__48779;
    wire N__48774;
    wire N__48771;
    wire N__48770;
    wire N__48767;
    wire N__48764;
    wire N__48759;
    wire N__48756;
    wire N__48753;
    wire N__48750;
    wire N__48747;
    wire N__48746;
    wire N__48745;
    wire N__48742;
    wire N__48737;
    wire N__48732;
    wire N__48729;
    wire N__48728;
    wire N__48725;
    wire N__48722;
    wire N__48719;
    wire N__48718;
    wire N__48717;
    wire N__48714;
    wire N__48713;
    wire N__48710;
    wire N__48707;
    wire N__48704;
    wire N__48701;
    wire N__48698;
    wire N__48687;
    wire N__48684;
    wire N__48683;
    wire N__48680;
    wire N__48677;
    wire N__48674;
    wire N__48673;
    wire N__48668;
    wire N__48665;
    wire N__48660;
    wire N__48659;
    wire N__48656;
    wire N__48653;
    wire N__48652;
    wire N__48647;
    wire N__48644;
    wire N__48641;
    wire N__48638;
    wire N__48635;
    wire N__48632;
    wire N__48629;
    wire N__48626;
    wire N__48621;
    wire N__48620;
    wire N__48617;
    wire N__48616;
    wire N__48615;
    wire N__48614;
    wire N__48611;
    wire N__48608;
    wire N__48603;
    wire N__48598;
    wire N__48591;
    wire N__48588;
    wire N__48585;
    wire N__48582;
    wire N__48579;
    wire N__48576;
    wire N__48573;
    wire N__48572;
    wire N__48571;
    wire N__48570;
    wire N__48567;
    wire N__48566;
    wire N__48561;
    wire N__48558;
    wire N__48555;
    wire N__48552;
    wire N__48549;
    wire N__48546;
    wire N__48543;
    wire N__48534;
    wire N__48533;
    wire N__48532;
    wire N__48529;
    wire N__48526;
    wire N__48523;
    wire N__48518;
    wire N__48513;
    wire N__48510;
    wire N__48507;
    wire N__48504;
    wire N__48501;
    wire N__48500;
    wire N__48497;
    wire N__48494;
    wire N__48489;
    wire N__48486;
    wire N__48483;
    wire N__48482;
    wire N__48477;
    wire N__48474;
    wire N__48473;
    wire N__48472;
    wire N__48469;
    wire N__48466;
    wire N__48465;
    wire N__48462;
    wire N__48457;
    wire N__48454;
    wire N__48447;
    wire N__48446;
    wire N__48443;
    wire N__48440;
    wire N__48437;
    wire N__48434;
    wire N__48431;
    wire N__48426;
    wire N__48425;
    wire N__48422;
    wire N__48421;
    wire N__48420;
    wire N__48419;
    wire N__48418;
    wire N__48417;
    wire N__48416;
    wire N__48413;
    wire N__48412;
    wire N__48411;
    wire N__48410;
    wire N__48409;
    wire N__48406;
    wire N__48405;
    wire N__48404;
    wire N__48401;
    wire N__48396;
    wire N__48393;
    wire N__48392;
    wire N__48389;
    wire N__48388;
    wire N__48385;
    wire N__48384;
    wire N__48383;
    wire N__48382;
    wire N__48381;
    wire N__48380;
    wire N__48379;
    wire N__48376;
    wire N__48373;
    wire N__48372;
    wire N__48371;
    wire N__48368;
    wire N__48365;
    wire N__48362;
    wire N__48359;
    wire N__48356;
    wire N__48353;
    wire N__48348;
    wire N__48343;
    wire N__48340;
    wire N__48337;
    wire N__48334;
    wire N__48331;
    wire N__48328;
    wire N__48325;
    wire N__48322;
    wire N__48319;
    wire N__48316;
    wire N__48315;
    wire N__48314;
    wire N__48313;
    wire N__48310;
    wire N__48307;
    wire N__48304;
    wire N__48303;
    wire N__48302;
    wire N__48299;
    wire N__48298;
    wire N__48295;
    wire N__48292;
    wire N__48285;
    wire N__48282;
    wire N__48279;
    wire N__48278;
    wire N__48277;
    wire N__48276;
    wire N__48273;
    wire N__48264;
    wire N__48259;
    wire N__48254;
    wire N__48247;
    wire N__48244;
    wire N__48241;
    wire N__48236;
    wire N__48233;
    wire N__48230;
    wire N__48225;
    wire N__48220;
    wire N__48217;
    wire N__48212;
    wire N__48205;
    wire N__48198;
    wire N__48187;
    wire N__48168;
    wire N__48167;
    wire N__48166;
    wire N__48165;
    wire N__48164;
    wire N__48161;
    wire N__48158;
    wire N__48157;
    wire N__48156;
    wire N__48155;
    wire N__48154;
    wire N__48153;
    wire N__48152;
    wire N__48151;
    wire N__48150;
    wire N__48145;
    wire N__48144;
    wire N__48141;
    wire N__48138;
    wire N__48135;
    wire N__48134;
    wire N__48133;
    wire N__48132;
    wire N__48131;
    wire N__48130;
    wire N__48129;
    wire N__48128;
    wire N__48127;
    wire N__48124;
    wire N__48123;
    wire N__48122;
    wire N__48121;
    wire N__48118;
    wire N__48115;
    wire N__48114;
    wire N__48113;
    wire N__48112;
    wire N__48111;
    wire N__48110;
    wire N__48101;
    wire N__48100;
    wire N__48099;
    wire N__48096;
    wire N__48093;
    wire N__48090;
    wire N__48089;
    wire N__48088;
    wire N__48085;
    wire N__48082;
    wire N__48079;
    wire N__48076;
    wire N__48073;
    wire N__48066;
    wire N__48059;
    wire N__48050;
    wire N__48047;
    wire N__48042;
    wire N__48039;
    wire N__48036;
    wire N__48033;
    wire N__48032;
    wire N__48029;
    wire N__48026;
    wire N__48023;
    wire N__48022;
    wire N__48021;
    wire N__48020;
    wire N__48017;
    wire N__48014;
    wire N__48011;
    wire N__48008;
    wire N__48003;
    wire N__47996;
    wire N__47993;
    wire N__47990;
    wire N__47987;
    wire N__47978;
    wire N__47971;
    wire N__47968;
    wire N__47965;
    wire N__47962;
    wire N__47959;
    wire N__47956;
    wire N__47953;
    wire N__47948;
    wire N__47941;
    wire N__47938;
    wire N__47935;
    wire N__47924;
    wire N__47901;
    wire N__47898;
    wire N__47895;
    wire N__47894;
    wire N__47891;
    wire N__47888;
    wire N__47885;
    wire N__47882;
    wire N__47877;
    wire N__47876;
    wire N__47875;
    wire N__47874;
    wire N__47873;
    wire N__47866;
    wire N__47861;
    wire N__47858;
    wire N__47853;
    wire N__47850;
    wire N__47847;
    wire N__47846;
    wire N__47843;
    wire N__47842;
    wire N__47841;
    wire N__47840;
    wire N__47839;
    wire N__47838;
    wire N__47835;
    wire N__47834;
    wire N__47833;
    wire N__47832;
    wire N__47831;
    wire N__47830;
    wire N__47829;
    wire N__47828;
    wire N__47827;
    wire N__47826;
    wire N__47825;
    wire N__47822;
    wire N__47821;
    wire N__47820;
    wire N__47819;
    wire N__47818;
    wire N__47817;
    wire N__47814;
    wire N__47813;
    wire N__47812;
    wire N__47811;
    wire N__47806;
    wire N__47805;
    wire N__47804;
    wire N__47803;
    wire N__47802;
    wire N__47797;
    wire N__47796;
    wire N__47795;
    wire N__47794;
    wire N__47793;
    wire N__47792;
    wire N__47791;
    wire N__47788;
    wire N__47787;
    wire N__47782;
    wire N__47777;
    wire N__47772;
    wire N__47769;
    wire N__47764;
    wire N__47761;
    wire N__47758;
    wire N__47755;
    wire N__47752;
    wire N__47749;
    wire N__47744;
    wire N__47741;
    wire N__47740;
    wire N__47733;
    wire N__47730;
    wire N__47723;
    wire N__47720;
    wire N__47717;
    wire N__47714;
    wire N__47709;
    wire N__47704;
    wire N__47701;
    wire N__47700;
    wire N__47697;
    wire N__47694;
    wire N__47689;
    wire N__47686;
    wire N__47681;
    wire N__47678;
    wire N__47677;
    wire N__47676;
    wire N__47675;
    wire N__47674;
    wire N__47673;
    wire N__47672;
    wire N__47671;
    wire N__47670;
    wire N__47669;
    wire N__47662;
    wire N__47657;
    wire N__47654;
    wire N__47653;
    wire N__47650;
    wire N__47637;
    wire N__47630;
    wire N__47627;
    wire N__47622;
    wire N__47613;
    wire N__47608;
    wire N__47599;
    wire N__47596;
    wire N__47591;
    wire N__47586;
    wire N__47583;
    wire N__47580;
    wire N__47575;
    wire N__47566;
    wire N__47547;
    wire N__47546;
    wire N__47543;
    wire N__47540;
    wire N__47537;
    wire N__47536;
    wire N__47533;
    wire N__47530;
    wire N__47527;
    wire N__47524;
    wire N__47517;
    wire N__47514;
    wire N__47513;
    wire N__47510;
    wire N__47509;
    wire N__47508;
    wire N__47507;
    wire N__47504;
    wire N__47501;
    wire N__47498;
    wire N__47497;
    wire N__47496;
    wire N__47495;
    wire N__47494;
    wire N__47489;
    wire N__47488;
    wire N__47487;
    wire N__47486;
    wire N__47485;
    wire N__47484;
    wire N__47483;
    wire N__47482;
    wire N__47481;
    wire N__47478;
    wire N__47473;
    wire N__47470;
    wire N__47465;
    wire N__47462;
    wire N__47459;
    wire N__47458;
    wire N__47455;
    wire N__47454;
    wire N__47451;
    wire N__47448;
    wire N__47445;
    wire N__47442;
    wire N__47439;
    wire N__47438;
    wire N__47435;
    wire N__47432;
    wire N__47431;
    wire N__47428;
    wire N__47423;
    wire N__47416;
    wire N__47413;
    wire N__47410;
    wire N__47407;
    wire N__47404;
    wire N__47395;
    wire N__47392;
    wire N__47387;
    wire N__47384;
    wire N__47379;
    wire N__47376;
    wire N__47365;
    wire N__47352;
    wire N__47349;
    wire N__47346;
    wire N__47343;
    wire N__47340;
    wire N__47337;
    wire N__47334;
    wire N__47331;
    wire N__47328;
    wire N__47325;
    wire N__47322;
    wire N__47321;
    wire N__47320;
    wire N__47317;
    wire N__47314;
    wire N__47313;
    wire N__47310;
    wire N__47307;
    wire N__47304;
    wire N__47301;
    wire N__47300;
    wire N__47297;
    wire N__47294;
    wire N__47289;
    wire N__47286;
    wire N__47277;
    wire N__47274;
    wire N__47271;
    wire N__47268;
    wire N__47265;
    wire N__47264;
    wire N__47263;
    wire N__47260;
    wire N__47257;
    wire N__47256;
    wire N__47253;
    wire N__47250;
    wire N__47247;
    wire N__47244;
    wire N__47241;
    wire N__47234;
    wire N__47231;
    wire N__47230;
    wire N__47227;
    wire N__47224;
    wire N__47221;
    wire N__47218;
    wire N__47211;
    wire N__47208;
    wire N__47205;
    wire N__47202;
    wire N__47199;
    wire N__47196;
    wire N__47195;
    wire N__47194;
    wire N__47191;
    wire N__47188;
    wire N__47185;
    wire N__47182;
    wire N__47179;
    wire N__47176;
    wire N__47173;
    wire N__47168;
    wire N__47163;
    wire N__47162;
    wire N__47157;
    wire N__47156;
    wire N__47153;
    wire N__47150;
    wire N__47147;
    wire N__47144;
    wire N__47141;
    wire N__47138;
    wire N__47133;
    wire N__47132;
    wire N__47131;
    wire N__47128;
    wire N__47125;
    wire N__47124;
    wire N__47121;
    wire N__47120;
    wire N__47119;
    wire N__47116;
    wire N__47113;
    wire N__47110;
    wire N__47107;
    wire N__47106;
    wire N__47103;
    wire N__47100;
    wire N__47097;
    wire N__47092;
    wire N__47089;
    wire N__47086;
    wire N__47085;
    wire N__47082;
    wire N__47075;
    wire N__47070;
    wire N__47067;
    wire N__47058;
    wire N__47055;
    wire N__47052;
    wire N__47049;
    wire N__47048;
    wire N__47045;
    wire N__47042;
    wire N__47039;
    wire N__47038;
    wire N__47035;
    wire N__47032;
    wire N__47029;
    wire N__47026;
    wire N__47019;
    wire N__47016;
    wire N__47015;
    wire N__47014;
    wire N__47013;
    wire N__47010;
    wire N__47007;
    wire N__47004;
    wire N__47001;
    wire N__46998;
    wire N__46997;
    wire N__46994;
    wire N__46991;
    wire N__46986;
    wire N__46983;
    wire N__46980;
    wire N__46977;
    wire N__46972;
    wire N__46965;
    wire N__46962;
    wire N__46959;
    wire N__46958;
    wire N__46955;
    wire N__46952;
    wire N__46947;
    wire N__46944;
    wire N__46943;
    wire N__46938;
    wire N__46935;
    wire N__46934;
    wire N__46933;
    wire N__46930;
    wire N__46927;
    wire N__46924;
    wire N__46923;
    wire N__46922;
    wire N__46919;
    wire N__46918;
    wire N__46915;
    wire N__46912;
    wire N__46909;
    wire N__46906;
    wire N__46905;
    wire N__46902;
    wire N__46899;
    wire N__46898;
    wire N__46895;
    wire N__46890;
    wire N__46887;
    wire N__46884;
    wire N__46881;
    wire N__46878;
    wire N__46875;
    wire N__46870;
    wire N__46867;
    wire N__46864;
    wire N__46859;
    wire N__46856;
    wire N__46853;
    wire N__46850;
    wire N__46847;
    wire N__46842;
    wire N__46833;
    wire N__46832;
    wire N__46829;
    wire N__46826;
    wire N__46825;
    wire N__46824;
    wire N__46821;
    wire N__46818;
    wire N__46817;
    wire N__46814;
    wire N__46811;
    wire N__46806;
    wire N__46803;
    wire N__46798;
    wire N__46795;
    wire N__46788;
    wire N__46785;
    wire N__46784;
    wire N__46781;
    wire N__46778;
    wire N__46773;
    wire N__46770;
    wire N__46767;
    wire N__46766;
    wire N__46763;
    wire N__46760;
    wire N__46759;
    wire N__46754;
    wire N__46751;
    wire N__46750;
    wire N__46747;
    wire N__46744;
    wire N__46741;
    wire N__46734;
    wire N__46731;
    wire N__46728;
    wire N__46727;
    wire N__46726;
    wire N__46723;
    wire N__46720;
    wire N__46717;
    wire N__46714;
    wire N__46711;
    wire N__46704;
    wire N__46703;
    wire N__46700;
    wire N__46697;
    wire N__46696;
    wire N__46695;
    wire N__46690;
    wire N__46687;
    wire N__46684;
    wire N__46681;
    wire N__46678;
    wire N__46675;
    wire N__46670;
    wire N__46667;
    wire N__46662;
    wire N__46659;
    wire N__46658;
    wire N__46655;
    wire N__46652;
    wire N__46647;
    wire N__46646;
    wire N__46643;
    wire N__46640;
    wire N__46637;
    wire N__46634;
    wire N__46631;
    wire N__46628;
    wire N__46627;
    wire N__46626;
    wire N__46623;
    wire N__46620;
    wire N__46617;
    wire N__46614;
    wire N__46611;
    wire N__46606;
    wire N__46599;
    wire N__46596;
    wire N__46593;
    wire N__46590;
    wire N__46589;
    wire N__46586;
    wire N__46583;
    wire N__46578;
    wire N__46575;
    wire N__46574;
    wire N__46571;
    wire N__46568;
    wire N__46565;
    wire N__46562;
    wire N__46559;
    wire N__46554;
    wire N__46551;
    wire N__46548;
    wire N__46547;
    wire N__46546;
    wire N__46543;
    wire N__46540;
    wire N__46537;
    wire N__46530;
    wire N__46529;
    wire N__46526;
    wire N__46523;
    wire N__46518;
    wire N__46517;
    wire N__46512;
    wire N__46509;
    wire N__46508;
    wire N__46507;
    wire N__46506;
    wire N__46503;
    wire N__46500;
    wire N__46497;
    wire N__46494;
    wire N__46491;
    wire N__46488;
    wire N__46483;
    wire N__46480;
    wire N__46477;
    wire N__46476;
    wire N__46473;
    wire N__46470;
    wire N__46467;
    wire N__46464;
    wire N__46461;
    wire N__46456;
    wire N__46449;
    wire N__46446;
    wire N__46443;
    wire N__46440;
    wire N__46437;
    wire N__46434;
    wire N__46431;
    wire N__46428;
    wire N__46425;
    wire N__46422;
    wire N__46419;
    wire N__46416;
    wire N__46415;
    wire N__46414;
    wire N__46413;
    wire N__46410;
    wire N__46407;
    wire N__46404;
    wire N__46403;
    wire N__46402;
    wire N__46401;
    wire N__46400;
    wire N__46397;
    wire N__46392;
    wire N__46389;
    wire N__46386;
    wire N__46383;
    wire N__46380;
    wire N__46379;
    wire N__46376;
    wire N__46375;
    wire N__46372;
    wire N__46369;
    wire N__46360;
    wire N__46357;
    wire N__46354;
    wire N__46351;
    wire N__46346;
    wire N__46343;
    wire N__46332;
    wire N__46329;
    wire N__46326;
    wire N__46323;
    wire N__46322;
    wire N__46321;
    wire N__46316;
    wire N__46315;
    wire N__46314;
    wire N__46313;
    wire N__46310;
    wire N__46307;
    wire N__46300;
    wire N__46299;
    wire N__46298;
    wire N__46297;
    wire N__46296;
    wire N__46295;
    wire N__46294;
    wire N__46293;
    wire N__46292;
    wire N__46291;
    wire N__46290;
    wire N__46289;
    wire N__46288;
    wire N__46285;
    wire N__46280;
    wire N__46277;
    wire N__46274;
    wire N__46267;
    wire N__46262;
    wire N__46259;
    wire N__46256;
    wire N__46255;
    wire N__46254;
    wire N__46253;
    wire N__46252;
    wire N__46251;
    wire N__46250;
    wire N__46247;
    wire N__46244;
    wire N__46241;
    wire N__46234;
    wire N__46227;
    wire N__46222;
    wire N__46219;
    wire N__46216;
    wire N__46211;
    wire N__46206;
    wire N__46201;
    wire N__46196;
    wire N__46191;
    wire N__46176;
    wire N__46173;
    wire N__46170;
    wire N__46167;
    wire N__46164;
    wire N__46161;
    wire N__46158;
    wire N__46155;
    wire N__46154;
    wire N__46153;
    wire N__46150;
    wire N__46147;
    wire N__46144;
    wire N__46137;
    wire N__46134;
    wire N__46131;
    wire N__46128;
    wire N__46125;
    wire N__46124;
    wire N__46123;
    wire N__46122;
    wire N__46121;
    wire N__46120;
    wire N__46119;
    wire N__46112;
    wire N__46111;
    wire N__46106;
    wire N__46101;
    wire N__46098;
    wire N__46095;
    wire N__46086;
    wire N__46085;
    wire N__46084;
    wire N__46081;
    wire N__46078;
    wire N__46075;
    wire N__46070;
    wire N__46067;
    wire N__46062;
    wire N__46059;
    wire N__46056;
    wire N__46055;
    wire N__46052;
    wire N__46051;
    wire N__46048;
    wire N__46045;
    wire N__46042;
    wire N__46035;
    wire N__46032;
    wire N__46029;
    wire N__46026;
    wire N__46023;
    wire N__46022;
    wire N__46021;
    wire N__46018;
    wire N__46015;
    wire N__46012;
    wire N__46005;
    wire N__46002;
    wire N__45999;
    wire N__45996;
    wire N__45993;
    wire N__45990;
    wire N__45987;
    wire N__45986;
    wire N__45985;
    wire N__45982;
    wire N__45979;
    wire N__45976;
    wire N__45973;
    wire N__45966;
    wire N__45965;
    wire N__45964;
    wire N__45963;
    wire N__45962;
    wire N__45961;
    wire N__45960;
    wire N__45959;
    wire N__45958;
    wire N__45955;
    wire N__45952;
    wire N__45949;
    wire N__45946;
    wire N__45945;
    wire N__45942;
    wire N__45941;
    wire N__45940;
    wire N__45937;
    wire N__45934;
    wire N__45931;
    wire N__45928;
    wire N__45927;
    wire N__45926;
    wire N__45925;
    wire N__45924;
    wire N__45915;
    wire N__45912;
    wire N__45909;
    wire N__45904;
    wire N__45895;
    wire N__45894;
    wire N__45891;
    wire N__45884;
    wire N__45881;
    wire N__45872;
    wire N__45869;
    wire N__45866;
    wire N__45859;
    wire N__45852;
    wire N__45849;
    wire N__45846;
    wire N__45843;
    wire N__45840;
    wire N__45839;
    wire N__45838;
    wire N__45837;
    wire N__45836;
    wire N__45833;
    wire N__45830;
    wire N__45827;
    wire N__45824;
    wire N__45821;
    wire N__45818;
    wire N__45813;
    wire N__45810;
    wire N__45807;
    wire N__45802;
    wire N__45797;
    wire N__45792;
    wire N__45789;
    wire N__45786;
    wire N__45785;
    wire N__45784;
    wire N__45781;
    wire N__45778;
    wire N__45775;
    wire N__45768;
    wire N__45765;
    wire N__45762;
    wire N__45759;
    wire N__45756;
    wire N__45753;
    wire N__45750;
    wire N__45747;
    wire N__45744;
    wire N__45743;
    wire N__45740;
    wire N__45737;
    wire N__45734;
    wire N__45733;
    wire N__45732;
    wire N__45729;
    wire N__45728;
    wire N__45727;
    wire N__45724;
    wire N__45719;
    wire N__45716;
    wire N__45711;
    wire N__45708;
    wire N__45705;
    wire N__45696;
    wire N__45693;
    wire N__45690;
    wire N__45687;
    wire N__45684;
    wire N__45681;
    wire N__45678;
    wire N__45675;
    wire N__45672;
    wire N__45671;
    wire N__45670;
    wire N__45667;
    wire N__45662;
    wire N__45657;
    wire N__45656;
    wire N__45653;
    wire N__45650;
    wire N__45647;
    wire N__45646;
    wire N__45643;
    wire N__45640;
    wire N__45637;
    wire N__45634;
    wire N__45631;
    wire N__45626;
    wire N__45621;
    wire N__45620;
    wire N__45617;
    wire N__45616;
    wire N__45615;
    wire N__45614;
    wire N__45611;
    wire N__45608;
    wire N__45605;
    wire N__45600;
    wire N__45591;
    wire N__45590;
    wire N__45587;
    wire N__45584;
    wire N__45579;
    wire N__45576;
    wire N__45573;
    wire N__45570;
    wire N__45569;
    wire N__45568;
    wire N__45565;
    wire N__45562;
    wire N__45559;
    wire N__45552;
    wire N__45549;
    wire N__45546;
    wire N__45543;
    wire N__45542;
    wire N__45541;
    wire N__45538;
    wire N__45535;
    wire N__45532;
    wire N__45529;
    wire N__45522;
    wire N__45519;
    wire N__45516;
    wire N__45513;
    wire N__45510;
    wire N__45509;
    wire N__45506;
    wire N__45503;
    wire N__45500;
    wire N__45495;
    wire N__45494;
    wire N__45491;
    wire N__45488;
    wire N__45485;
    wire N__45482;
    wire N__45479;
    wire N__45476;
    wire N__45473;
    wire N__45468;
    wire N__45465;
    wire N__45464;
    wire N__45463;
    wire N__45460;
    wire N__45457;
    wire N__45454;
    wire N__45451;
    wire N__45448;
    wire N__45441;
    wire N__45438;
    wire N__45435;
    wire N__45434;
    wire N__45433;
    wire N__45430;
    wire N__45425;
    wire N__45420;
    wire N__45417;
    wire N__45414;
    wire N__45413;
    wire N__45410;
    wire N__45407;
    wire N__45406;
    wire N__45405;
    wire N__45402;
    wire N__45399;
    wire N__45398;
    wire N__45393;
    wire N__45388;
    wire N__45385;
    wire N__45378;
    wire N__45375;
    wire N__45372;
    wire N__45369;
    wire N__45366;
    wire N__45363;
    wire N__45360;
    wire N__45357;
    wire N__45354;
    wire N__45351;
    wire N__45348;
    wire N__45345;
    wire N__45342;
    wire N__45339;
    wire N__45336;
    wire N__45333;
    wire N__45330;
    wire N__45327;
    wire N__45324;
    wire N__45323;
    wire N__45318;
    wire N__45315;
    wire N__45312;
    wire N__45309;
    wire N__45308;
    wire N__45305;
    wire N__45302;
    wire N__45299;
    wire N__45294;
    wire N__45293;
    wire N__45290;
    wire N__45287;
    wire N__45284;
    wire N__45281;
    wire N__45278;
    wire N__45275;
    wire N__45272;
    wire N__45267;
    wire N__45264;
    wire N__45263;
    wire N__45262;
    wire N__45261;
    wire N__45260;
    wire N__45259;
    wire N__45258;
    wire N__45255;
    wire N__45252;
    wire N__45247;
    wire N__45244;
    wire N__45241;
    wire N__45238;
    wire N__45235;
    wire N__45230;
    wire N__45227;
    wire N__45224;
    wire N__45221;
    wire N__45220;
    wire N__45219;
    wire N__45218;
    wire N__45217;
    wire N__45216;
    wire N__45211;
    wire N__45208;
    wire N__45203;
    wire N__45200;
    wire N__45191;
    wire N__45188;
    wire N__45177;
    wire N__45176;
    wire N__45175;
    wire N__45172;
    wire N__45169;
    wire N__45166;
    wire N__45163;
    wire N__45160;
    wire N__45157;
    wire N__45156;
    wire N__45153;
    wire N__45150;
    wire N__45147;
    wire N__45144;
    wire N__45135;
    wire N__45134;
    wire N__45133;
    wire N__45132;
    wire N__45131;
    wire N__45130;
    wire N__45127;
    wire N__45124;
    wire N__45121;
    wire N__45120;
    wire N__45113;
    wire N__45110;
    wire N__45107;
    wire N__45104;
    wire N__45101;
    wire N__45098;
    wire N__45097;
    wire N__45094;
    wire N__45089;
    wire N__45086;
    wire N__45083;
    wire N__45080;
    wire N__45077;
    wire N__45074;
    wire N__45071;
    wire N__45068;
    wire N__45065;
    wire N__45054;
    wire N__45051;
    wire N__45050;
    wire N__45047;
    wire N__45044;
    wire N__45041;
    wire N__45036;
    wire N__45033;
    wire N__45032;
    wire N__45031;
    wire N__45030;
    wire N__45029;
    wire N__45028;
    wire N__45025;
    wire N__45022;
    wire N__45021;
    wire N__45020;
    wire N__45019;
    wire N__45018;
    wire N__45017;
    wire N__45014;
    wire N__45011;
    wire N__45008;
    wire N__45005;
    wire N__45002;
    wire N__44999;
    wire N__44996;
    wire N__44993;
    wire N__44992;
    wire N__44991;
    wire N__44990;
    wire N__44987;
    wire N__44986;
    wire N__44983;
    wire N__44982;
    wire N__44979;
    wire N__44978;
    wire N__44977;
    wire N__44976;
    wire N__44975;
    wire N__44972;
    wire N__44967;
    wire N__44964;
    wire N__44955;
    wire N__44952;
    wire N__44949;
    wire N__44946;
    wire N__44945;
    wire N__44942;
    wire N__44939;
    wire N__44936;
    wire N__44933;
    wire N__44932;
    wire N__44931;
    wire N__44928;
    wire N__44925;
    wire N__44922;
    wire N__44919;
    wire N__44916;
    wire N__44915;
    wire N__44912;
    wire N__44907;
    wire N__44898;
    wire N__44895;
    wire N__44892;
    wire N__44889;
    wire N__44884;
    wire N__44881;
    wire N__44878;
    wire N__44871;
    wire N__44866;
    wire N__44863;
    wire N__44862;
    wire N__44859;
    wire N__44854;
    wire N__44851;
    wire N__44840;
    wire N__44833;
    wire N__44830;
    wire N__44817;
    wire N__44814;
    wire N__44813;
    wire N__44812;
    wire N__44811;
    wire N__44808;
    wire N__44805;
    wire N__44802;
    wire N__44801;
    wire N__44800;
    wire N__44799;
    wire N__44798;
    wire N__44795;
    wire N__44792;
    wire N__44787;
    wire N__44784;
    wire N__44781;
    wire N__44778;
    wire N__44777;
    wire N__44776;
    wire N__44773;
    wire N__44772;
    wire N__44769;
    wire N__44768;
    wire N__44757;
    wire N__44754;
    wire N__44751;
    wire N__44748;
    wire N__44745;
    wire N__44742;
    wire N__44739;
    wire N__44738;
    wire N__44737;
    wire N__44730;
    wire N__44725;
    wire N__44724;
    wire N__44719;
    wire N__44718;
    wire N__44715;
    wire N__44714;
    wire N__44711;
    wire N__44706;
    wire N__44703;
    wire N__44702;
    wire N__44699;
    wire N__44696;
    wire N__44693;
    wire N__44690;
    wire N__44687;
    wire N__44682;
    wire N__44679;
    wire N__44678;
    wire N__44677;
    wire N__44676;
    wire N__44675;
    wire N__44674;
    wire N__44673;
    wire N__44668;
    wire N__44663;
    wire N__44656;
    wire N__44653;
    wire N__44650;
    wire N__44647;
    wire N__44644;
    wire N__44641;
    wire N__44638;
    wire N__44619;
    wire N__44618;
    wire N__44617;
    wire N__44616;
    wire N__44615;
    wire N__44612;
    wire N__44611;
    wire N__44610;
    wire N__44607;
    wire N__44606;
    wire N__44605;
    wire N__44604;
    wire N__44603;
    wire N__44602;
    wire N__44601;
    wire N__44600;
    wire N__44599;
    wire N__44596;
    wire N__44593;
    wire N__44590;
    wire N__44587;
    wire N__44584;
    wire N__44583;
    wire N__44580;
    wire N__44577;
    wire N__44574;
    wire N__44573;
    wire N__44570;
    wire N__44567;
    wire N__44566;
    wire N__44565;
    wire N__44564;
    wire N__44561;
    wire N__44558;
    wire N__44555;
    wire N__44552;
    wire N__44549;
    wire N__44546;
    wire N__44543;
    wire N__44542;
    wire N__44539;
    wire N__44536;
    wire N__44533;
    wire N__44530;
    wire N__44523;
    wire N__44520;
    wire N__44517;
    wire N__44514;
    wire N__44513;
    wire N__44512;
    wire N__44511;
    wire N__44510;
    wire N__44507;
    wire N__44504;
    wire N__44501;
    wire N__44498;
    wire N__44493;
    wire N__44486;
    wire N__44483;
    wire N__44480;
    wire N__44473;
    wire N__44470;
    wire N__44467;
    wire N__44460;
    wire N__44457;
    wire N__44454;
    wire N__44451;
    wire N__44448;
    wire N__44445;
    wire N__44442;
    wire N__44437;
    wire N__44430;
    wire N__44425;
    wire N__44424;
    wire N__44415;
    wire N__44414;
    wire N__44407;
    wire N__44400;
    wire N__44395;
    wire N__44392;
    wire N__44389;
    wire N__44386;
    wire N__44373;
    wire N__44372;
    wire N__44371;
    wire N__44366;
    wire N__44363;
    wire N__44360;
    wire N__44357;
    wire N__44354;
    wire N__44349;
    wire N__44346;
    wire N__44343;
    wire N__44340;
    wire N__44337;
    wire N__44334;
    wire N__44333;
    wire N__44328;
    wire N__44325;
    wire N__44322;
    wire N__44319;
    wire N__44316;
    wire N__44313;
    wire N__44310;
    wire N__44307;
    wire N__44304;
    wire N__44301;
    wire N__44298;
    wire N__44295;
    wire N__44292;
    wire N__44289;
    wire N__44288;
    wire N__44287;
    wire N__44286;
    wire N__44285;
    wire N__44282;
    wire N__44279;
    wire N__44274;
    wire N__44271;
    wire N__44268;
    wire N__44265;
    wire N__44262;
    wire N__44259;
    wire N__44256;
    wire N__44253;
    wire N__44250;
    wire N__44245;
    wire N__44238;
    wire N__44235;
    wire N__44232;
    wire N__44229;
    wire N__44226;
    wire N__44223;
    wire N__44220;
    wire N__44217;
    wire N__44214;
    wire N__44213;
    wire N__44212;
    wire N__44209;
    wire N__44208;
    wire N__44205;
    wire N__44204;
    wire N__44203;
    wire N__44200;
    wire N__44197;
    wire N__44194;
    wire N__44193;
    wire N__44192;
    wire N__44191;
    wire N__44188;
    wire N__44181;
    wire N__44180;
    wire N__44179;
    wire N__44178;
    wire N__44173;
    wire N__44170;
    wire N__44167;
    wire N__44164;
    wire N__44161;
    wire N__44158;
    wire N__44155;
    wire N__44152;
    wire N__44149;
    wire N__44146;
    wire N__44139;
    wire N__44134;
    wire N__44121;
    wire N__44118;
    wire N__44115;
    wire N__44112;
    wire N__44109;
    wire N__44106;
    wire N__44105;
    wire N__44104;
    wire N__44103;
    wire N__44100;
    wire N__44099;
    wire N__44098;
    wire N__44097;
    wire N__44094;
    wire N__44091;
    wire N__44088;
    wire N__44085;
    wire N__44082;
    wire N__44079;
    wire N__44076;
    wire N__44075;
    wire N__44072;
    wire N__44069;
    wire N__44066;
    wire N__44063;
    wire N__44060;
    wire N__44055;
    wire N__44052;
    wire N__44049;
    wire N__44044;
    wire N__44039;
    wire N__44036;
    wire N__44033;
    wire N__44022;
    wire N__44019;
    wire N__44016;
    wire N__44015;
    wire N__44014;
    wire N__44011;
    wire N__44008;
    wire N__44005;
    wire N__44004;
    wire N__44003;
    wire N__44000;
    wire N__43999;
    wire N__43998;
    wire N__43993;
    wire N__43990;
    wire N__43987;
    wire N__43986;
    wire N__43985;
    wire N__43982;
    wire N__43977;
    wire N__43974;
    wire N__43965;
    wire N__43956;
    wire N__43953;
    wire N__43952;
    wire N__43951;
    wire N__43950;
    wire N__43947;
    wire N__43942;
    wire N__43939;
    wire N__43938;
    wire N__43937;
    wire N__43936;
    wire N__43933;
    wire N__43930;
    wire N__43927;
    wire N__43924;
    wire N__43919;
    wire N__43908;
    wire N__43905;
    wire N__43902;
    wire N__43899;
    wire N__43896;
    wire N__43893;
    wire N__43890;
    wire N__43887;
    wire N__43884;
    wire N__43881;
    wire N__43880;
    wire N__43877;
    wire N__43874;
    wire N__43871;
    wire N__43868;
    wire N__43863;
    wire N__43862;
    wire N__43859;
    wire N__43856;
    wire N__43851;
    wire N__43848;
    wire N__43845;
    wire N__43844;
    wire N__43843;
    wire N__43842;
    wire N__43841;
    wire N__43840;
    wire N__43837;
    wire N__43836;
    wire N__43831;
    wire N__43828;
    wire N__43825;
    wire N__43822;
    wire N__43819;
    wire N__43816;
    wire N__43815;
    wire N__43814;
    wire N__43813;
    wire N__43810;
    wire N__43807;
    wire N__43804;
    wire N__43801;
    wire N__43796;
    wire N__43793;
    wire N__43788;
    wire N__43785;
    wire N__43778;
    wire N__43775;
    wire N__43764;
    wire N__43761;
    wire N__43758;
    wire N__43757;
    wire N__43754;
    wire N__43751;
    wire N__43748;
    wire N__43743;
    wire N__43740;
    wire N__43737;
    wire N__43736;
    wire N__43733;
    wire N__43730;
    wire N__43727;
    wire N__43724;
    wire N__43719;
    wire N__43718;
    wire N__43717;
    wire N__43716;
    wire N__43715;
    wire N__43712;
    wire N__43709;
    wire N__43706;
    wire N__43703;
    wire N__43700;
    wire N__43697;
    wire N__43694;
    wire N__43693;
    wire N__43690;
    wire N__43687;
    wire N__43684;
    wire N__43681;
    wire N__43678;
    wire N__43675;
    wire N__43668;
    wire N__43665;
    wire N__43662;
    wire N__43657;
    wire N__43650;
    wire N__43647;
    wire N__43646;
    wire N__43643;
    wire N__43640;
    wire N__43637;
    wire N__43634;
    wire N__43629;
    wire N__43626;
    wire N__43625;
    wire N__43624;
    wire N__43621;
    wire N__43616;
    wire N__43613;
    wire N__43608;
    wire N__43605;
    wire N__43602;
    wire N__43601;
    wire N__43598;
    wire N__43595;
    wire N__43592;
    wire N__43587;
    wire N__43584;
    wire N__43581;
    wire N__43578;
    wire N__43575;
    wire N__43574;
    wire N__43571;
    wire N__43568;
    wire N__43563;
    wire N__43560;
    wire N__43557;
    wire N__43554;
    wire N__43551;
    wire N__43550;
    wire N__43549;
    wire N__43546;
    wire N__43543;
    wire N__43540;
    wire N__43533;
    wire N__43530;
    wire N__43529;
    wire N__43526;
    wire N__43523;
    wire N__43518;
    wire N__43515;
    wire N__43512;
    wire N__43511;
    wire N__43508;
    wire N__43505;
    wire N__43502;
    wire N__43497;
    wire N__43494;
    wire N__43491;
    wire N__43488;
    wire N__43485;
    wire N__43482;
    wire N__43479;
    wire N__43476;
    wire N__43473;
    wire N__43470;
    wire N__43469;
    wire N__43466;
    wire N__43465;
    wire N__43462;
    wire N__43459;
    wire N__43456;
    wire N__43453;
    wire N__43450;
    wire N__43447;
    wire N__43444;
    wire N__43441;
    wire N__43438;
    wire N__43431;
    wire N__43428;
    wire N__43425;
    wire N__43422;
    wire N__43419;
    wire N__43416;
    wire N__43415;
    wire N__43410;
    wire N__43407;
    wire N__43406;
    wire N__43403;
    wire N__43400;
    wire N__43399;
    wire N__43398;
    wire N__43395;
    wire N__43392;
    wire N__43387;
    wire N__43386;
    wire N__43383;
    wire N__43378;
    wire N__43375;
    wire N__43372;
    wire N__43369;
    wire N__43362;
    wire N__43361;
    wire N__43360;
    wire N__43359;
    wire N__43358;
    wire N__43353;
    wire N__43350;
    wire N__43345;
    wire N__43342;
    wire N__43337;
    wire N__43334;
    wire N__43331;
    wire N__43326;
    wire N__43323;
    wire N__43320;
    wire N__43317;
    wire N__43314;
    wire N__43313;
    wire N__43310;
    wire N__43309;
    wire N__43308;
    wire N__43305;
    wire N__43302;
    wire N__43297;
    wire N__43290;
    wire N__43287;
    wire N__43284;
    wire N__43281;
    wire N__43280;
    wire N__43277;
    wire N__43274;
    wire N__43271;
    wire N__43266;
    wire N__43265;
    wire N__43264;
    wire N__43261;
    wire N__43256;
    wire N__43253;
    wire N__43250;
    wire N__43245;
    wire N__43242;
    wire N__43239;
    wire N__43236;
    wire N__43233;
    wire N__43230;
    wire N__43229;
    wire N__43226;
    wire N__43225;
    wire N__43222;
    wire N__43219;
    wire N__43216;
    wire N__43211;
    wire N__43206;
    wire N__43203;
    wire N__43200;
    wire N__43197;
    wire N__43194;
    wire N__43191;
    wire N__43190;
    wire N__43187;
    wire N__43184;
    wire N__43183;
    wire N__43180;
    wire N__43177;
    wire N__43174;
    wire N__43171;
    wire N__43164;
    wire N__43161;
    wire N__43158;
    wire N__43157;
    wire N__43154;
    wire N__43151;
    wire N__43150;
    wire N__43147;
    wire N__43144;
    wire N__43141;
    wire N__43138;
    wire N__43131;
    wire N__43128;
    wire N__43125;
    wire N__43122;
    wire N__43119;
    wire N__43118;
    wire N__43115;
    wire N__43114;
    wire N__43111;
    wire N__43108;
    wire N__43105;
    wire N__43100;
    wire N__43097;
    wire N__43094;
    wire N__43089;
    wire N__43086;
    wire N__43083;
    wire N__43080;
    wire N__43077;
    wire N__43076;
    wire N__43075;
    wire N__43072;
    wire N__43069;
    wire N__43066;
    wire N__43059;
    wire N__43056;
    wire N__43053;
    wire N__43050;
    wire N__43047;
    wire N__43044;
    wire N__43043;
    wire N__43042;
    wire N__43041;
    wire N__43040;
    wire N__43039;
    wire N__43038;
    wire N__43035;
    wire N__43030;
    wire N__43027;
    wire N__43022;
    wire N__43019;
    wire N__43008;
    wire N__43005;
    wire N__43002;
    wire N__42999;
    wire N__42996;
    wire N__42993;
    wire N__42990;
    wire N__42989;
    wire N__42986;
    wire N__42985;
    wire N__42982;
    wire N__42979;
    wire N__42976;
    wire N__42973;
    wire N__42966;
    wire N__42963;
    wire N__42962;
    wire N__42961;
    wire N__42958;
    wire N__42955;
    wire N__42952;
    wire N__42945;
    wire N__42942;
    wire N__42939;
    wire N__42936;
    wire N__42935;
    wire N__42934;
    wire N__42931;
    wire N__42928;
    wire N__42925;
    wire N__42918;
    wire N__42915;
    wire N__42912;
    wire N__42909;
    wire N__42906;
    wire N__42905;
    wire N__42902;
    wire N__42899;
    wire N__42894;
    wire N__42891;
    wire N__42888;
    wire N__42887;
    wire N__42884;
    wire N__42881;
    wire N__42876;
    wire N__42875;
    wire N__42874;
    wire N__42871;
    wire N__42868;
    wire N__42865;
    wire N__42862;
    wire N__42855;
    wire N__42852;
    wire N__42849;
    wire N__42846;
    wire N__42845;
    wire N__42844;
    wire N__42843;
    wire N__42842;
    wire N__42841;
    wire N__42838;
    wire N__42835;
    wire N__42832;
    wire N__42825;
    wire N__42816;
    wire N__42813;
    wire N__42810;
    wire N__42807;
    wire N__42806;
    wire N__42803;
    wire N__42800;
    wire N__42797;
    wire N__42794;
    wire N__42793;
    wire N__42790;
    wire N__42787;
    wire N__42784;
    wire N__42781;
    wire N__42778;
    wire N__42775;
    wire N__42768;
    wire N__42765;
    wire N__42762;
    wire N__42761;
    wire N__42758;
    wire N__42755;
    wire N__42752;
    wire N__42747;
    wire N__42744;
    wire N__42741;
    wire N__42738;
    wire N__42735;
    wire N__42734;
    wire N__42731;
    wire N__42728;
    wire N__42723;
    wire N__42720;
    wire N__42717;
    wire N__42716;
    wire N__42713;
    wire N__42710;
    wire N__42707;
    wire N__42702;
    wire N__42699;
    wire N__42698;
    wire N__42695;
    wire N__42692;
    wire N__42687;
    wire N__42684;
    wire N__42681;
    wire N__42678;
    wire N__42675;
    wire N__42672;
    wire N__42671;
    wire N__42670;
    wire N__42667;
    wire N__42662;
    wire N__42657;
    wire N__42656;
    wire N__42655;
    wire N__42650;
    wire N__42647;
    wire N__42642;
    wire N__42641;
    wire N__42640;
    wire N__42637;
    wire N__42636;
    wire N__42633;
    wire N__42630;
    wire N__42627;
    wire N__42626;
    wire N__42625;
    wire N__42624;
    wire N__42621;
    wire N__42618;
    wire N__42615;
    wire N__42612;
    wire N__42607;
    wire N__42602;
    wire N__42591;
    wire N__42588;
    wire N__42585;
    wire N__42584;
    wire N__42583;
    wire N__42580;
    wire N__42579;
    wire N__42578;
    wire N__42575;
    wire N__42572;
    wire N__42569;
    wire N__42564;
    wire N__42555;
    wire N__42554;
    wire N__42551;
    wire N__42550;
    wire N__42547;
    wire N__42546;
    wire N__42543;
    wire N__42540;
    wire N__42537;
    wire N__42534;
    wire N__42531;
    wire N__42522;
    wire N__42519;
    wire N__42518;
    wire N__42515;
    wire N__42512;
    wire N__42509;
    wire N__42506;
    wire N__42503;
    wire N__42500;
    wire N__42497;
    wire N__42492;
    wire N__42489;
    wire N__42486;
    wire N__42483;
    wire N__42480;
    wire N__42477;
    wire N__42474;
    wire N__42471;
    wire N__42468;
    wire N__42465;
    wire N__42462;
    wire N__42461;
    wire N__42460;
    wire N__42457;
    wire N__42456;
    wire N__42453;
    wire N__42452;
    wire N__42449;
    wire N__42448;
    wire N__42447;
    wire N__42446;
    wire N__42443;
    wire N__42438;
    wire N__42435;
    wire N__42432;
    wire N__42429;
    wire N__42426;
    wire N__42423;
    wire N__42418;
    wire N__42415;
    wire N__42412;
    wire N__42405;
    wire N__42402;
    wire N__42399;
    wire N__42396;
    wire N__42393;
    wire N__42390;
    wire N__42387;
    wire N__42382;
    wire N__42377;
    wire N__42374;
    wire N__42369;
    wire N__42368;
    wire N__42367;
    wire N__42366;
    wire N__42365;
    wire N__42358;
    wire N__42355;
    wire N__42352;
    wire N__42351;
    wire N__42350;
    wire N__42345;
    wire N__42342;
    wire N__42339;
    wire N__42336;
    wire N__42327;
    wire N__42324;
    wire N__42323;
    wire N__42320;
    wire N__42317;
    wire N__42312;
    wire N__42309;
    wire N__42306;
    wire N__42303;
    wire N__42300;
    wire N__42297;
    wire N__42294;
    wire N__42293;
    wire N__42290;
    wire N__42287;
    wire N__42284;
    wire N__42281;
    wire N__42276;
    wire N__42273;
    wire N__42270;
    wire N__42267;
    wire N__42264;
    wire N__42261;
    wire N__42258;
    wire N__42255;
    wire N__42252;
    wire N__42249;
    wire N__42246;
    wire N__42243;
    wire N__42240;
    wire N__42237;
    wire N__42234;
    wire N__42231;
    wire N__42228;
    wire N__42225;
    wire N__42222;
    wire N__42219;
    wire N__42216;
    wire N__42213;
    wire N__42210;
    wire N__42207;
    wire N__42204;
    wire N__42201;
    wire N__42198;
    wire N__42195;
    wire N__42192;
    wire N__42189;
    wire N__42186;
    wire N__42183;
    wire N__42180;
    wire N__42177;
    wire N__42176;
    wire N__42171;
    wire N__42168;
    wire N__42167;
    wire N__42164;
    wire N__42161;
    wire N__42158;
    wire N__42155;
    wire N__42150;
    wire N__42147;
    wire N__42144;
    wire N__42143;
    wire N__42140;
    wire N__42137;
    wire N__42136;
    wire N__42133;
    wire N__42130;
    wire N__42129;
    wire N__42126;
    wire N__42123;
    wire N__42120;
    wire N__42117;
    wire N__42108;
    wire N__42105;
    wire N__42102;
    wire N__42099;
    wire N__42096;
    wire N__42095;
    wire N__42094;
    wire N__42093;
    wire N__42090;
    wire N__42087;
    wire N__42086;
    wire N__42085;
    wire N__42084;
    wire N__42081;
    wire N__42078;
    wire N__42075;
    wire N__42072;
    wire N__42069;
    wire N__42066;
    wire N__42063;
    wire N__42060;
    wire N__42057;
    wire N__42054;
    wire N__42053;
    wire N__42050;
    wire N__42047;
    wire N__42044;
    wire N__42041;
    wire N__42040;
    wire N__42035;
    wire N__42032;
    wire N__42029;
    wire N__42024;
    wire N__42019;
    wire N__42016;
    wire N__42015;
    wire N__42014;
    wire N__42011;
    wire N__42006;
    wire N__42003;
    wire N__42000;
    wire N__41997;
    wire N__41994;
    wire N__41991;
    wire N__41976;
    wire N__41973;
    wire N__41972;
    wire N__41969;
    wire N__41968;
    wire N__41967;
    wire N__41964;
    wire N__41961;
    wire N__41958;
    wire N__41957;
    wire N__41956;
    wire N__41953;
    wire N__41950;
    wire N__41947;
    wire N__41946;
    wire N__41943;
    wire N__41938;
    wire N__41935;
    wire N__41932;
    wire N__41929;
    wire N__41926;
    wire N__41919;
    wire N__41916;
    wire N__41907;
    wire N__41906;
    wire N__41905;
    wire N__41904;
    wire N__41903;
    wire N__41892;
    wire N__41891;
    wire N__41890;
    wire N__41889;
    wire N__41888;
    wire N__41887;
    wire N__41886;
    wire N__41885;
    wire N__41884;
    wire N__41883;
    wire N__41882;
    wire N__41881;
    wire N__41880;
    wire N__41879;
    wire N__41878;
    wire N__41877;
    wire N__41876;
    wire N__41875;
    wire N__41874;
    wire N__41873;
    wire N__41872;
    wire N__41871;
    wire N__41870;
    wire N__41869;
    wire N__41868;
    wire N__41867;
    wire N__41866;
    wire N__41865;
    wire N__41864;
    wire N__41863;
    wire N__41862;
    wire N__41861;
    wire N__41860;
    wire N__41859;
    wire N__41858;
    wire N__41855;
    wire N__41854;
    wire N__41853;
    wire N__41852;
    wire N__41851;
    wire N__41850;
    wire N__41849;
    wire N__41848;
    wire N__41847;
    wire N__41846;
    wire N__41845;
    wire N__41844;
    wire N__41843;
    wire N__41842;
    wire N__41841;
    wire N__41840;
    wire N__41839;
    wire N__41838;
    wire N__41837;
    wire N__41836;
    wire N__41825;
    wire N__41814;
    wire N__41801;
    wire N__41794;
    wire N__41779;
    wire N__41766;
    wire N__41765;
    wire N__41760;
    wire N__41757;
    wire N__41742;
    wire N__41741;
    wire N__41730;
    wire N__41715;
    wire N__41704;
    wire N__41701;
    wire N__41700;
    wire N__41697;
    wire N__41694;
    wire N__41689;
    wire N__41686;
    wire N__41683;
    wire N__41676;
    wire N__41675;
    wire N__41674;
    wire N__41673;
    wire N__41672;
    wire N__41671;
    wire N__41670;
    wire N__41669;
    wire N__41668;
    wire N__41665;
    wire N__41662;
    wire N__41657;
    wire N__41654;
    wire N__41649;
    wire N__41636;
    wire N__41633;
    wire N__41630;
    wire N__41613;
    wire N__41610;
    wire N__41607;
    wire N__41606;
    wire N__41605;
    wire N__41602;
    wire N__41599;
    wire N__41596;
    wire N__41593;
    wire N__41592;
    wire N__41589;
    wire N__41586;
    wire N__41583;
    wire N__41580;
    wire N__41577;
    wire N__41570;
    wire N__41567;
    wire N__41564;
    wire N__41559;
    wire N__41556;
    wire N__41553;
    wire N__41552;
    wire N__41549;
    wire N__41546;
    wire N__41545;
    wire N__41542;
    wire N__41539;
    wire N__41536;
    wire N__41529;
    wire N__41526;
    wire N__41525;
    wire N__41524;
    wire N__41519;
    wire N__41516;
    wire N__41511;
    wire N__41508;
    wire N__41505;
    wire N__41502;
    wire N__41499;
    wire N__41498;
    wire N__41495;
    wire N__41494;
    wire N__41493;
    wire N__41492;
    wire N__41491;
    wire N__41482;
    wire N__41479;
    wire N__41478;
    wire N__41475;
    wire N__41474;
    wire N__41473;
    wire N__41472;
    wire N__41469;
    wire N__41458;
    wire N__41457;
    wire N__41454;
    wire N__41449;
    wire N__41446;
    wire N__41445;
    wire N__41442;
    wire N__41437;
    wire N__41434;
    wire N__41427;
    wire N__41424;
    wire N__41423;
    wire N__41422;
    wire N__41421;
    wire N__41420;
    wire N__41419;
    wire N__41418;
    wire N__41417;
    wire N__41414;
    wire N__41411;
    wire N__41408;
    wire N__41407;
    wire N__41404;
    wire N__41401;
    wire N__41400;
    wire N__41397;
    wire N__41396;
    wire N__41393;
    wire N__41390;
    wire N__41389;
    wire N__41386;
    wire N__41383;
    wire N__41374;
    wire N__41363;
    wire N__41362;
    wire N__41359;
    wire N__41354;
    wire N__41349;
    wire N__41346;
    wire N__41337;
    wire N__41336;
    wire N__41335;
    wire N__41334;
    wire N__41333;
    wire N__41332;
    wire N__41323;
    wire N__41322;
    wire N__41321;
    wire N__41320;
    wire N__41319;
    wire N__41318;
    wire N__41315;
    wire N__41312;
    wire N__41309;
    wire N__41298;
    wire N__41297;
    wire N__41296;
    wire N__41293;
    wire N__41290;
    wire N__41285;
    wire N__41282;
    wire N__41279;
    wire N__41268;
    wire N__41265;
    wire N__41264;
    wire N__41263;
    wire N__41260;
    wire N__41257;
    wire N__41254;
    wire N__41251;
    wire N__41248;
    wire N__41245;
    wire N__41242;
    wire N__41235;
    wire N__41232;
    wire N__41229;
    wire N__41228;
    wire N__41227;
    wire N__41224;
    wire N__41221;
    wire N__41218;
    wire N__41215;
    wire N__41208;
    wire N__41205;
    wire N__41202;
    wire N__41199;
    wire N__41196;
    wire N__41193;
    wire N__41192;
    wire N__41189;
    wire N__41188;
    wire N__41185;
    wire N__41182;
    wire N__41179;
    wire N__41176;
    wire N__41169;
    wire N__41166;
    wire N__41163;
    wire N__41160;
    wire N__41157;
    wire N__41156;
    wire N__41153;
    wire N__41150;
    wire N__41149;
    wire N__41146;
    wire N__41145;
    wire N__41144;
    wire N__41141;
    wire N__41138;
    wire N__41135;
    wire N__41132;
    wire N__41129;
    wire N__41126;
    wire N__41123;
    wire N__41118;
    wire N__41109;
    wire N__41108;
    wire N__41107;
    wire N__41106;
    wire N__41105;
    wire N__41102;
    wire N__41099;
    wire N__41098;
    wire N__41093;
    wire N__41090;
    wire N__41087;
    wire N__41084;
    wire N__41081;
    wire N__41078;
    wire N__41075;
    wire N__41072;
    wire N__41065;
    wire N__41060;
    wire N__41055;
    wire N__41052;
    wire N__41049;
    wire N__41046;
    wire N__41043;
    wire N__41040;
    wire N__41037;
    wire N__41034;
    wire N__41033;
    wire N__41032;
    wire N__41031;
    wire N__41030;
    wire N__41027;
    wire N__41024;
    wire N__41021;
    wire N__41018;
    wire N__41015;
    wire N__41012;
    wire N__41009;
    wire N__41006;
    wire N__41003;
    wire N__41000;
    wire N__40989;
    wire N__40988;
    wire N__40985;
    wire N__40984;
    wire N__40979;
    wire N__40978;
    wire N__40975;
    wire N__40972;
    wire N__40969;
    wire N__40966;
    wire N__40963;
    wire N__40960;
    wire N__40953;
    wire N__40952;
    wire N__40947;
    wire N__40944;
    wire N__40941;
    wire N__40938;
    wire N__40935;
    wire N__40934;
    wire N__40933;
    wire N__40930;
    wire N__40929;
    wire N__40926;
    wire N__40925;
    wire N__40922;
    wire N__40919;
    wire N__40914;
    wire N__40911;
    wire N__40908;
    wire N__40903;
    wire N__40896;
    wire N__40893;
    wire N__40892;
    wire N__40891;
    wire N__40888;
    wire N__40885;
    wire N__40882;
    wire N__40879;
    wire N__40876;
    wire N__40873;
    wire N__40868;
    wire N__40865;
    wire N__40864;
    wire N__40863;
    wire N__40858;
    wire N__40855;
    wire N__40852;
    wire N__40849;
    wire N__40842;
    wire N__40839;
    wire N__40836;
    wire N__40833;
    wire N__40830;
    wire N__40827;
    wire N__40824;
    wire N__40821;
    wire N__40820;
    wire N__40815;
    wire N__40814;
    wire N__40811;
    wire N__40808;
    wire N__40807;
    wire N__40802;
    wire N__40799;
    wire N__40798;
    wire N__40797;
    wire N__40796;
    wire N__40795;
    wire N__40794;
    wire N__40793;
    wire N__40792;
    wire N__40789;
    wire N__40786;
    wire N__40773;
    wire N__40770;
    wire N__40761;
    wire N__40760;
    wire N__40759;
    wire N__40756;
    wire N__40753;
    wire N__40750;
    wire N__40747;
    wire N__40744;
    wire N__40741;
    wire N__40738;
    wire N__40731;
    wire N__40728;
    wire N__40725;
    wire N__40722;
    wire N__40719;
    wire N__40718;
    wire N__40715;
    wire N__40712;
    wire N__40711;
    wire N__40706;
    wire N__40703;
    wire N__40702;
    wire N__40699;
    wire N__40694;
    wire N__40689;
    wire N__40686;
    wire N__40683;
    wire N__40680;
    wire N__40677;
    wire N__40674;
    wire N__40673;
    wire N__40672;
    wire N__40669;
    wire N__40664;
    wire N__40663;
    wire N__40660;
    wire N__40657;
    wire N__40654;
    wire N__40651;
    wire N__40648;
    wire N__40645;
    wire N__40642;
    wire N__40639;
    wire N__40632;
    wire N__40629;
    wire N__40626;
    wire N__40625;
    wire N__40624;
    wire N__40623;
    wire N__40620;
    wire N__40619;
    wire N__40618;
    wire N__40615;
    wire N__40614;
    wire N__40611;
    wire N__40610;
    wire N__40607;
    wire N__40606;
    wire N__40601;
    wire N__40600;
    wire N__40599;
    wire N__40598;
    wire N__40595;
    wire N__40592;
    wire N__40587;
    wire N__40584;
    wire N__40579;
    wire N__40578;
    wire N__40577;
    wire N__40574;
    wire N__40571;
    wire N__40568;
    wire N__40567;
    wire N__40564;
    wire N__40561;
    wire N__40558;
    wire N__40553;
    wire N__40550;
    wire N__40545;
    wire N__40538;
    wire N__40535;
    wire N__40528;
    wire N__40525;
    wire N__40518;
    wire N__40509;
    wire N__40506;
    wire N__40505;
    wire N__40504;
    wire N__40503;
    wire N__40502;
    wire N__40501;
    wire N__40500;
    wire N__40499;
    wire N__40496;
    wire N__40493;
    wire N__40490;
    wire N__40487;
    wire N__40484;
    wire N__40481;
    wire N__40478;
    wire N__40475;
    wire N__40472;
    wire N__40467;
    wire N__40464;
    wire N__40461;
    wire N__40458;
    wire N__40455;
    wire N__40450;
    wire N__40445;
    wire N__40434;
    wire N__40433;
    wire N__40432;
    wire N__40431;
    wire N__40430;
    wire N__40429;
    wire N__40428;
    wire N__40427;
    wire N__40426;
    wire N__40425;
    wire N__40424;
    wire N__40423;
    wire N__40422;
    wire N__40421;
    wire N__40420;
    wire N__40419;
    wire N__40418;
    wire N__40415;
    wire N__40412;
    wire N__40411;
    wire N__40410;
    wire N__40409;
    wire N__40408;
    wire N__40407;
    wire N__40406;
    wire N__40403;
    wire N__40400;
    wire N__40397;
    wire N__40390;
    wire N__40387;
    wire N__40382;
    wire N__40379;
    wire N__40374;
    wire N__40367;
    wire N__40358;
    wire N__40349;
    wire N__40346;
    wire N__40341;
    wire N__40338;
    wire N__40317;
    wire N__40316;
    wire N__40315;
    wire N__40314;
    wire N__40313;
    wire N__40310;
    wire N__40305;
    wire N__40300;
    wire N__40293;
    wire N__40290;
    wire N__40287;
    wire N__40286;
    wire N__40283;
    wire N__40280;
    wire N__40277;
    wire N__40274;
    wire N__40273;
    wire N__40272;
    wire N__40267;
    wire N__40264;
    wire N__40261;
    wire N__40258;
    wire N__40255;
    wire N__40248;
    wire N__40247;
    wire N__40246;
    wire N__40245;
    wire N__40244;
    wire N__40243;
    wire N__40240;
    wire N__40239;
    wire N__40236;
    wire N__40235;
    wire N__40234;
    wire N__40227;
    wire N__40224;
    wire N__40221;
    wire N__40220;
    wire N__40219;
    wire N__40216;
    wire N__40213;
    wire N__40208;
    wire N__40203;
    wire N__40200;
    wire N__40199;
    wire N__40198;
    wire N__40197;
    wire N__40194;
    wire N__40193;
    wire N__40192;
    wire N__40189;
    wire N__40186;
    wire N__40181;
    wire N__40176;
    wire N__40171;
    wire N__40168;
    wire N__40161;
    wire N__40146;
    wire N__40145;
    wire N__40144;
    wire N__40143;
    wire N__40142;
    wire N__40141;
    wire N__40140;
    wire N__40137;
    wire N__40134;
    wire N__40129;
    wire N__40126;
    wire N__40121;
    wire N__40118;
    wire N__40107;
    wire N__40104;
    wire N__40103;
    wire N__40100;
    wire N__40097;
    wire N__40094;
    wire N__40093;
    wire N__40090;
    wire N__40089;
    wire N__40086;
    wire N__40083;
    wire N__40080;
    wire N__40079;
    wire N__40076;
    wire N__40071;
    wire N__40068;
    wire N__40063;
    wire N__40060;
    wire N__40057;
    wire N__40050;
    wire N__40049;
    wire N__40046;
    wire N__40043;
    wire N__40040;
    wire N__40037;
    wire N__40034;
    wire N__40031;
    wire N__40026;
    wire N__40023;
    wire N__40022;
    wire N__40021;
    wire N__40020;
    wire N__40019;
    wire N__40016;
    wire N__40011;
    wire N__40006;
    wire N__39999;
    wire N__39998;
    wire N__39995;
    wire N__39994;
    wire N__39993;
    wire N__39990;
    wire N__39987;
    wire N__39984;
    wire N__39983;
    wire N__39980;
    wire N__39977;
    wire N__39972;
    wire N__39969;
    wire N__39966;
    wire N__39957;
    wire N__39954;
    wire N__39951;
    wire N__39948;
    wire N__39947;
    wire N__39946;
    wire N__39945;
    wire N__39944;
    wire N__39943;
    wire N__39940;
    wire N__39937;
    wire N__39936;
    wire N__39935;
    wire N__39934;
    wire N__39929;
    wire N__39924;
    wire N__39921;
    wire N__39918;
    wire N__39915;
    wire N__39910;
    wire N__39905;
    wire N__39902;
    wire N__39899;
    wire N__39896;
    wire N__39893;
    wire N__39890;
    wire N__39879;
    wire N__39878;
    wire N__39877;
    wire N__39876;
    wire N__39875;
    wire N__39874;
    wire N__39871;
    wire N__39866;
    wire N__39863;
    wire N__39860;
    wire N__39857;
    wire N__39846;
    wire N__39845;
    wire N__39844;
    wire N__39841;
    wire N__39838;
    wire N__39837;
    wire N__39836;
    wire N__39835;
    wire N__39832;
    wire N__39831;
    wire N__39828;
    wire N__39827;
    wire N__39826;
    wire N__39825;
    wire N__39824;
    wire N__39821;
    wire N__39818;
    wire N__39815;
    wire N__39812;
    wire N__39807;
    wire N__39804;
    wire N__39795;
    wire N__39792;
    wire N__39789;
    wire N__39782;
    wire N__39779;
    wire N__39776;
    wire N__39773;
    wire N__39768;
    wire N__39759;
    wire N__39758;
    wire N__39755;
    wire N__39754;
    wire N__39753;
    wire N__39750;
    wire N__39747;
    wire N__39742;
    wire N__39739;
    wire N__39734;
    wire N__39729;
    wire N__39726;
    wire N__39725;
    wire N__39724;
    wire N__39719;
    wire N__39716;
    wire N__39711;
    wire N__39708;
    wire N__39705;
    wire N__39702;
    wire N__39701;
    wire N__39698;
    wire N__39697;
    wire N__39694;
    wire N__39693;
    wire N__39690;
    wire N__39687;
    wire N__39684;
    wire N__39683;
    wire N__39680;
    wire N__39679;
    wire N__39678;
    wire N__39675;
    wire N__39672;
    wire N__39669;
    wire N__39666;
    wire N__39663;
    wire N__39660;
    wire N__39657;
    wire N__39652;
    wire N__39649;
    wire N__39646;
    wire N__39643;
    wire N__39640;
    wire N__39637;
    wire N__39624;
    wire N__39623;
    wire N__39622;
    wire N__39619;
    wire N__39616;
    wire N__39613;
    wire N__39612;
    wire N__39609;
    wire N__39606;
    wire N__39603;
    wire N__39600;
    wire N__39593;
    wire N__39588;
    wire N__39585;
    wire N__39582;
    wire N__39579;
    wire N__39576;
    wire N__39573;
    wire N__39572;
    wire N__39569;
    wire N__39566;
    wire N__39563;
    wire N__39560;
    wire N__39555;
    wire N__39554;
    wire N__39553;
    wire N__39552;
    wire N__39549;
    wire N__39546;
    wire N__39545;
    wire N__39542;
    wire N__39541;
    wire N__39538;
    wire N__39535;
    wire N__39530;
    wire N__39527;
    wire N__39524;
    wire N__39523;
    wire N__39520;
    wire N__39519;
    wire N__39516;
    wire N__39511;
    wire N__39508;
    wire N__39505;
    wire N__39502;
    wire N__39499;
    wire N__39492;
    wire N__39489;
    wire N__39480;
    wire N__39479;
    wire N__39478;
    wire N__39477;
    wire N__39476;
    wire N__39473;
    wire N__39470;
    wire N__39469;
    wire N__39466;
    wire N__39463;
    wire N__39462;
    wire N__39459;
    wire N__39456;
    wire N__39453;
    wire N__39450;
    wire N__39447;
    wire N__39446;
    wire N__39443;
    wire N__39440;
    wire N__39433;
    wire N__39430;
    wire N__39427;
    wire N__39424;
    wire N__39421;
    wire N__39418;
    wire N__39415;
    wire N__39410;
    wire N__39407;
    wire N__39396;
    wire N__39395;
    wire N__39394;
    wire N__39391;
    wire N__39390;
    wire N__39389;
    wire N__39388;
    wire N__39387;
    wire N__39386;
    wire N__39385;
    wire N__39382;
    wire N__39379;
    wire N__39376;
    wire N__39373;
    wire N__39372;
    wire N__39371;
    wire N__39370;
    wire N__39363;
    wire N__39362;
    wire N__39361;
    wire N__39360;
    wire N__39359;
    wire N__39354;
    wire N__39351;
    wire N__39348;
    wire N__39343;
    wire N__39336;
    wire N__39333;
    wire N__39330;
    wire N__39327;
    wire N__39324;
    wire N__39321;
    wire N__39318;
    wire N__39311;
    wire N__39306;
    wire N__39303;
    wire N__39288;
    wire N__39285;
    wire N__39282;
    wire N__39281;
    wire N__39278;
    wire N__39275;
    wire N__39272;
    wire N__39267;
    wire N__39264;
    wire N__39263;
    wire N__39260;
    wire N__39259;
    wire N__39258;
    wire N__39255;
    wire N__39252;
    wire N__39249;
    wire N__39246;
    wire N__39243;
    wire N__39238;
    wire N__39235;
    wire N__39232;
    wire N__39229;
    wire N__39222;
    wire N__39221;
    wire N__39220;
    wire N__39219;
    wire N__39218;
    wire N__39217;
    wire N__39216;
    wire N__39215;
    wire N__39214;
    wire N__39213;
    wire N__39212;
    wire N__39211;
    wire N__39210;
    wire N__39209;
    wire N__39208;
    wire N__39207;
    wire N__39206;
    wire N__39205;
    wire N__39204;
    wire N__39201;
    wire N__39200;
    wire N__39195;
    wire N__39194;
    wire N__39191;
    wire N__39190;
    wire N__39187;
    wire N__39186;
    wire N__39185;
    wire N__39184;
    wire N__39179;
    wire N__39174;
    wire N__39163;
    wire N__39160;
    wire N__39157;
    wire N__39154;
    wire N__39149;
    wire N__39146;
    wire N__39143;
    wire N__39142;
    wire N__39139;
    wire N__39136;
    wire N__39133;
    wire N__39132;
    wire N__39131;
    wire N__39130;
    wire N__39129;
    wire N__39126;
    wire N__39119;
    wire N__39116;
    wire N__39103;
    wire N__39096;
    wire N__39095;
    wire N__39094;
    wire N__39093;
    wire N__39090;
    wire N__39087;
    wire N__39082;
    wire N__39079;
    wire N__39072;
    wire N__39067;
    wire N__39060;
    wire N__39059;
    wire N__39056;
    wire N__39051;
    wire N__39044;
    wire N__39037;
    wire N__39034;
    wire N__39031;
    wire N__39030;
    wire N__39025;
    wire N__39022;
    wire N__39017;
    wire N__39016;
    wire N__39013;
    wire N__39010;
    wire N__39007;
    wire N__39004;
    wire N__39001;
    wire N__38998;
    wire N__38985;
    wire N__38982;
    wire N__38979;
    wire N__38978;
    wire N__38977;
    wire N__38974;
    wire N__38971;
    wire N__38968;
    wire N__38967;
    wire N__38964;
    wire N__38961;
    wire N__38958;
    wire N__38955;
    wire N__38950;
    wire N__38947;
    wire N__38940;
    wire N__38939;
    wire N__38936;
    wire N__38933;
    wire N__38932;
    wire N__38929;
    wire N__38926;
    wire N__38923;
    wire N__38922;
    wire N__38919;
    wire N__38914;
    wire N__38911;
    wire N__38906;
    wire N__38901;
    wire N__38900;
    wire N__38899;
    wire N__38896;
    wire N__38893;
    wire N__38892;
    wire N__38889;
    wire N__38886;
    wire N__38885;
    wire N__38882;
    wire N__38879;
    wire N__38876;
    wire N__38873;
    wire N__38870;
    wire N__38867;
    wire N__38864;
    wire N__38853;
    wire N__38850;
    wire N__38849;
    wire N__38846;
    wire N__38843;
    wire N__38840;
    wire N__38835;
    wire N__38832;
    wire N__38829;
    wire N__38828;
    wire N__38827;
    wire N__38824;
    wire N__38823;
    wire N__38822;
    wire N__38819;
    wire N__38816;
    wire N__38813;
    wire N__38808;
    wire N__38803;
    wire N__38796;
    wire N__38793;
    wire N__38790;
    wire N__38789;
    wire N__38786;
    wire N__38783;
    wire N__38778;
    wire N__38775;
    wire N__38772;
    wire N__38771;
    wire N__38766;
    wire N__38763;
    wire N__38760;
    wire N__38757;
    wire N__38756;
    wire N__38753;
    wire N__38750;
    wire N__38745;
    wire N__38744;
    wire N__38741;
    wire N__38738;
    wire N__38733;
    wire N__38730;
    wire N__38727;
    wire N__38726;
    wire N__38721;
    wire N__38718;
    wire N__38715;
    wire N__38712;
    wire N__38711;
    wire N__38708;
    wire N__38703;
    wire N__38700;
    wire N__38697;
    wire N__38694;
    wire N__38691;
    wire N__38690;
    wire N__38687;
    wire N__38684;
    wire N__38681;
    wire N__38676;
    wire N__38675;
    wire N__38672;
    wire N__38669;
    wire N__38664;
    wire N__38663;
    wire N__38662;
    wire N__38661;
    wire N__38660;
    wire N__38657;
    wire N__38654;
    wire N__38653;
    wire N__38652;
    wire N__38649;
    wire N__38648;
    wire N__38647;
    wire N__38646;
    wire N__38643;
    wire N__38640;
    wire N__38639;
    wire N__38638;
    wire N__38637;
    wire N__38636;
    wire N__38635;
    wire N__38632;
    wire N__38625;
    wire N__38622;
    wire N__38615;
    wire N__38608;
    wire N__38605;
    wire N__38598;
    wire N__38595;
    wire N__38580;
    wire N__38579;
    wire N__38578;
    wire N__38571;
    wire N__38570;
    wire N__38569;
    wire N__38568;
    wire N__38567;
    wire N__38566;
    wire N__38565;
    wire N__38564;
    wire N__38563;
    wire N__38562;
    wire N__38561;
    wire N__38560;
    wire N__38559;
    wire N__38558;
    wire N__38555;
    wire N__38552;
    wire N__38543;
    wire N__38534;
    wire N__38527;
    wire N__38524;
    wire N__38511;
    wire N__38508;
    wire N__38505;
    wire N__38504;
    wire N__38501;
    wire N__38498;
    wire N__38493;
    wire N__38492;
    wire N__38489;
    wire N__38486;
    wire N__38481;
    wire N__38478;
    wire N__38475;
    wire N__38472;
    wire N__38469;
    wire N__38466;
    wire N__38463;
    wire N__38460;
    wire N__38457;
    wire N__38454;
    wire N__38453;
    wire N__38450;
    wire N__38447;
    wire N__38442;
    wire N__38439;
    wire N__38438;
    wire N__38435;
    wire N__38432;
    wire N__38427;
    wire N__38424;
    wire N__38421;
    wire N__38418;
    wire N__38415;
    wire N__38414;
    wire N__38411;
    wire N__38408;
    wire N__38405;
    wire N__38402;
    wire N__38397;
    wire N__38394;
    wire N__38393;
    wire N__38390;
    wire N__38387;
    wire N__38384;
    wire N__38381;
    wire N__38376;
    wire N__38373;
    wire N__38370;
    wire N__38369;
    wire N__38366;
    wire N__38361;
    wire N__38358;
    wire N__38355;
    wire N__38352;
    wire N__38349;
    wire N__38346;
    wire N__38343;
    wire N__38342;
    wire N__38341;
    wire N__38340;
    wire N__38337;
    wire N__38332;
    wire N__38329;
    wire N__38322;
    wire N__38319;
    wire N__38316;
    wire N__38313;
    wire N__38310;
    wire N__38307;
    wire N__38304;
    wire N__38301;
    wire N__38298;
    wire N__38295;
    wire N__38292;
    wire N__38289;
    wire N__38286;
    wire N__38283;
    wire N__38280;
    wire N__38277;
    wire N__38274;
    wire N__38271;
    wire N__38268;
    wire N__38265;
    wire N__38264;
    wire N__38261;
    wire N__38258;
    wire N__38253;
    wire N__38250;
    wire N__38249;
    wire N__38246;
    wire N__38243;
    wire N__38240;
    wire N__38235;
    wire N__38232;
    wire N__38229;
    wire N__38226;
    wire N__38223;
    wire N__38220;
    wire N__38217;
    wire N__38214;
    wire N__38211;
    wire N__38208;
    wire N__38205;
    wire N__38202;
    wire N__38199;
    wire N__38196;
    wire N__38193;
    wire N__38190;
    wire N__38187;
    wire N__38184;
    wire N__38181;
    wire N__38178;
    wire N__38175;
    wire N__38172;
    wire N__38169;
    wire N__38166;
    wire N__38163;
    wire N__38160;
    wire N__38157;
    wire N__38154;
    wire N__38153;
    wire N__38150;
    wire N__38147;
    wire N__38144;
    wire N__38141;
    wire N__38136;
    wire N__38135;
    wire N__38132;
    wire N__38127;
    wire N__38124;
    wire N__38121;
    wire N__38120;
    wire N__38117;
    wire N__38114;
    wire N__38111;
    wire N__38108;
    wire N__38103;
    wire N__38100;
    wire N__38099;
    wire N__38096;
    wire N__38093;
    wire N__38090;
    wire N__38087;
    wire N__38082;
    wire N__38079;
    wire N__38076;
    wire N__38073;
    wire N__38070;
    wire N__38069;
    wire N__38066;
    wire N__38065;
    wire N__38062;
    wire N__38059;
    wire N__38056;
    wire N__38053;
    wire N__38050;
    wire N__38043;
    wire N__38040;
    wire N__38037;
    wire N__38034;
    wire N__38031;
    wire N__38028;
    wire N__38025;
    wire N__38022;
    wire N__38019;
    wire N__38018;
    wire N__38015;
    wire N__38012;
    wire N__38009;
    wire N__38006;
    wire N__38001;
    wire N__37998;
    wire N__37995;
    wire N__37994;
    wire N__37991;
    wire N__37988;
    wire N__37983;
    wire N__37980;
    wire N__37977;
    wire N__37974;
    wire N__37973;
    wire N__37970;
    wire N__37967;
    wire N__37962;
    wire N__37961;
    wire N__37956;
    wire N__37953;
    wire N__37950;
    wire N__37949;
    wire N__37948;
    wire N__37947;
    wire N__37938;
    wire N__37935;
    wire N__37934;
    wire N__37933;
    wire N__37930;
    wire N__37925;
    wire N__37920;
    wire N__37919;
    wire N__37918;
    wire N__37917;
    wire N__37908;
    wire N__37907;
    wire N__37904;
    wire N__37903;
    wire N__37902;
    wire N__37899;
    wire N__37896;
    wire N__37891;
    wire N__37888;
    wire N__37885;
    wire N__37882;
    wire N__37875;
    wire N__37872;
    wire N__37869;
    wire N__37868;
    wire N__37865;
    wire N__37862;
    wire N__37857;
    wire N__37854;
    wire N__37853;
    wire N__37852;
    wire N__37851;
    wire N__37848;
    wire N__37841;
    wire N__37836;
    wire N__37833;
    wire N__37830;
    wire N__37829;
    wire N__37826;
    wire N__37823;
    wire N__37818;
    wire N__37815;
    wire N__37812;
    wire N__37809;
    wire N__37808;
    wire N__37805;
    wire N__37802;
    wire N__37797;
    wire N__37794;
    wire N__37793;
    wire N__37790;
    wire N__37787;
    wire N__37784;
    wire N__37781;
    wire N__37778;
    wire N__37773;
    wire N__37770;
    wire N__37767;
    wire N__37766;
    wire N__37765;
    wire N__37758;
    wire N__37755;
    wire N__37752;
    wire N__37749;
    wire N__37746;
    wire N__37745;
    wire N__37742;
    wire N__37741;
    wire N__37740;
    wire N__37737;
    wire N__37736;
    wire N__37735;
    wire N__37734;
    wire N__37733;
    wire N__37732;
    wire N__37731;
    wire N__37730;
    wire N__37729;
    wire N__37728;
    wire N__37721;
    wire N__37718;
    wire N__37715;
    wire N__37710;
    wire N__37707;
    wire N__37704;
    wire N__37701;
    wire N__37696;
    wire N__37693;
    wire N__37692;
    wire N__37691;
    wire N__37690;
    wire N__37687;
    wire N__37682;
    wire N__37671;
    wire N__37668;
    wire N__37661;
    wire N__37658;
    wire N__37649;
    wire N__37644;
    wire N__37641;
    wire N__37638;
    wire N__37637;
    wire N__37636;
    wire N__37633;
    wire N__37630;
    wire N__37627;
    wire N__37624;
    wire N__37623;
    wire N__37622;
    wire N__37619;
    wire N__37616;
    wire N__37613;
    wire N__37610;
    wire N__37607;
    wire N__37600;
    wire N__37593;
    wire N__37590;
    wire N__37587;
    wire N__37584;
    wire N__37583;
    wire N__37582;
    wire N__37581;
    wire N__37580;
    wire N__37577;
    wire N__37574;
    wire N__37569;
    wire N__37568;
    wire N__37565;
    wire N__37562;
    wire N__37559;
    wire N__37556;
    wire N__37553;
    wire N__37550;
    wire N__37547;
    wire N__37542;
    wire N__37539;
    wire N__37536;
    wire N__37533;
    wire N__37524;
    wire N__37523;
    wire N__37520;
    wire N__37517;
    wire N__37514;
    wire N__37511;
    wire N__37508;
    wire N__37503;
    wire N__37502;
    wire N__37499;
    wire N__37496;
    wire N__37491;
    wire N__37488;
    wire N__37487;
    wire N__37484;
    wire N__37481;
    wire N__37478;
    wire N__37473;
    wire N__37472;
    wire N__37471;
    wire N__37468;
    wire N__37465;
    wire N__37464;
    wire N__37461;
    wire N__37458;
    wire N__37455;
    wire N__37452;
    wire N__37443;
    wire N__37440;
    wire N__37439;
    wire N__37438;
    wire N__37435;
    wire N__37430;
    wire N__37427;
    wire N__37422;
    wire N__37419;
    wire N__37418;
    wire N__37417;
    wire N__37414;
    wire N__37411;
    wire N__37408;
    wire N__37401;
    wire N__37398;
    wire N__37397;
    wire N__37396;
    wire N__37393;
    wire N__37390;
    wire N__37389;
    wire N__37386;
    wire N__37381;
    wire N__37380;
    wire N__37379;
    wire N__37378;
    wire N__37377;
    wire N__37376;
    wire N__37373;
    wire N__37370;
    wire N__37367;
    wire N__37364;
    wire N__37357;
    wire N__37354;
    wire N__37341;
    wire N__37338;
    wire N__37335;
    wire N__37334;
    wire N__37331;
    wire N__37328;
    wire N__37327;
    wire N__37324;
    wire N__37321;
    wire N__37318;
    wire N__37315;
    wire N__37308;
    wire N__37305;
    wire N__37302;
    wire N__37299;
    wire N__37296;
    wire N__37295;
    wire N__37292;
    wire N__37289;
    wire N__37286;
    wire N__37285;
    wire N__37282;
    wire N__37279;
    wire N__37276;
    wire N__37269;
    wire N__37266;
    wire N__37263;
    wire N__37260;
    wire N__37257;
    wire N__37254;
    wire N__37253;
    wire N__37252;
    wire N__37249;
    wire N__37246;
    wire N__37245;
    wire N__37242;
    wire N__37239;
    wire N__37238;
    wire N__37235;
    wire N__37232;
    wire N__37229;
    wire N__37226;
    wire N__37223;
    wire N__37220;
    wire N__37215;
    wire N__37212;
    wire N__37203;
    wire N__37200;
    wire N__37197;
    wire N__37194;
    wire N__37191;
    wire N__37188;
    wire N__37187;
    wire N__37186;
    wire N__37185;
    wire N__37182;
    wire N__37179;
    wire N__37176;
    wire N__37175;
    wire N__37174;
    wire N__37171;
    wire N__37168;
    wire N__37163;
    wire N__37160;
    wire N__37157;
    wire N__37156;
    wire N__37155;
    wire N__37152;
    wire N__37143;
    wire N__37140;
    wire N__37137;
    wire N__37132;
    wire N__37129;
    wire N__37126;
    wire N__37123;
    wire N__37120;
    wire N__37113;
    wire N__37112;
    wire N__37109;
    wire N__37106;
    wire N__37105;
    wire N__37102;
    wire N__37099;
    wire N__37096;
    wire N__37089;
    wire N__37088;
    wire N__37085;
    wire N__37082;
    wire N__37081;
    wire N__37080;
    wire N__37079;
    wire N__37078;
    wire N__37077;
    wire N__37074;
    wire N__37071;
    wire N__37062;
    wire N__37059;
    wire N__37050;
    wire N__37047;
    wire N__37046;
    wire N__37045;
    wire N__37044;
    wire N__37043;
    wire N__37040;
    wire N__37037;
    wire N__37034;
    wire N__37029;
    wire N__37026;
    wire N__37017;
    wire N__37014;
    wire N__37011;
    wire N__37010;
    wire N__37007;
    wire N__37004;
    wire N__36999;
    wire N__36996;
    wire N__36993;
    wire N__36992;
    wire N__36989;
    wire N__36986;
    wire N__36983;
    wire N__36978;
    wire N__36975;
    wire N__36972;
    wire N__36969;
    wire N__36966;
    wire N__36963;
    wire N__36960;
    wire N__36957;
    wire N__36954;
    wire N__36953;
    wire N__36950;
    wire N__36949;
    wire N__36948;
    wire N__36947;
    wire N__36944;
    wire N__36941;
    wire N__36938;
    wire N__36935;
    wire N__36932;
    wire N__36921;
    wire N__36918;
    wire N__36917;
    wire N__36914;
    wire N__36911;
    wire N__36906;
    wire N__36903;
    wire N__36902;
    wire N__36899;
    wire N__36898;
    wire N__36895;
    wire N__36892;
    wire N__36889;
    wire N__36882;
    wire N__36881;
    wire N__36878;
    wire N__36877;
    wire N__36876;
    wire N__36873;
    wire N__36870;
    wire N__36867;
    wire N__36864;
    wire N__36863;
    wire N__36862;
    wire N__36861;
    wire N__36858;
    wire N__36853;
    wire N__36850;
    wire N__36847;
    wire N__36844;
    wire N__36841;
    wire N__36840;
    wire N__36835;
    wire N__36830;
    wire N__36827;
    wire N__36824;
    wire N__36821;
    wire N__36818;
    wire N__36815;
    wire N__36804;
    wire N__36803;
    wire N__36802;
    wire N__36801;
    wire N__36800;
    wire N__36799;
    wire N__36798;
    wire N__36795;
    wire N__36790;
    wire N__36787;
    wire N__36782;
    wire N__36779;
    wire N__36778;
    wire N__36775;
    wire N__36770;
    wire N__36765;
    wire N__36762;
    wire N__36757;
    wire N__36754;
    wire N__36751;
    wire N__36748;
    wire N__36745;
    wire N__36738;
    wire N__36735;
    wire N__36732;
    wire N__36729;
    wire N__36726;
    wire N__36723;
    wire N__36720;
    wire N__36719;
    wire N__36718;
    wire N__36711;
    wire N__36710;
    wire N__36707;
    wire N__36704;
    wire N__36699;
    wire N__36696;
    wire N__36693;
    wire N__36690;
    wire N__36689;
    wire N__36688;
    wire N__36687;
    wire N__36684;
    wire N__36681;
    wire N__36680;
    wire N__36679;
    wire N__36676;
    wire N__36675;
    wire N__36670;
    wire N__36665;
    wire N__36662;
    wire N__36659;
    wire N__36656;
    wire N__36655;
    wire N__36652;
    wire N__36649;
    wire N__36646;
    wire N__36641;
    wire N__36638;
    wire N__36635;
    wire N__36632;
    wire N__36627;
    wire N__36618;
    wire N__36615;
    wire N__36612;
    wire N__36609;
    wire N__36606;
    wire N__36603;
    wire N__36600;
    wire N__36597;
    wire N__36594;
    wire N__36591;
    wire N__36588;
    wire N__36585;
    wire N__36582;
    wire N__36579;
    wire N__36576;
    wire N__36573;
    wire N__36570;
    wire N__36567;
    wire N__36564;
    wire N__36561;
    wire N__36558;
    wire N__36555;
    wire N__36552;
    wire N__36551;
    wire N__36548;
    wire N__36545;
    wire N__36542;
    wire N__36539;
    wire N__36536;
    wire N__36533;
    wire N__36528;
    wire N__36525;
    wire N__36522;
    wire N__36519;
    wire N__36516;
    wire N__36513;
    wire N__36510;
    wire N__36507;
    wire N__36504;
    wire N__36501;
    wire N__36498;
    wire N__36495;
    wire N__36492;
    wire N__36489;
    wire N__36486;
    wire N__36483;
    wire N__36480;
    wire N__36477;
    wire N__36474;
    wire N__36471;
    wire N__36468;
    wire N__36465;
    wire N__36462;
    wire N__36459;
    wire N__36456;
    wire N__36453;
    wire N__36450;
    wire N__36447;
    wire N__36444;
    wire N__36441;
    wire N__36438;
    wire N__36435;
    wire N__36432;
    wire N__36429;
    wire N__36426;
    wire N__36425;
    wire N__36422;
    wire N__36417;
    wire N__36414;
    wire N__36411;
    wire N__36410;
    wire N__36407;
    wire N__36404;
    wire N__36401;
    wire N__36398;
    wire N__36393;
    wire N__36392;
    wire N__36389;
    wire N__36386;
    wire N__36383;
    wire N__36378;
    wire N__36375;
    wire N__36372;
    wire N__36371;
    wire N__36370;
    wire N__36367;
    wire N__36362;
    wire N__36357;
    wire N__36354;
    wire N__36351;
    wire N__36348;
    wire N__36345;
    wire N__36342;
    wire N__36339;
    wire N__36338;
    wire N__36335;
    wire N__36332;
    wire N__36329;
    wire N__36326;
    wire N__36321;
    wire N__36318;
    wire N__36315;
    wire N__36314;
    wire N__36311;
    wire N__36308;
    wire N__36305;
    wire N__36302;
    wire N__36297;
    wire N__36294;
    wire N__36293;
    wire N__36290;
    wire N__36287;
    wire N__36284;
    wire N__36279;
    wire N__36276;
    wire N__36275;
    wire N__36272;
    wire N__36269;
    wire N__36266;
    wire N__36263;
    wire N__36258;
    wire N__36257;
    wire N__36254;
    wire N__36251;
    wire N__36246;
    wire N__36245;
    wire N__36242;
    wire N__36239;
    wire N__36236;
    wire N__36233;
    wire N__36230;
    wire N__36227;
    wire N__36226;
    wire N__36223;
    wire N__36220;
    wire N__36217;
    wire N__36210;
    wire N__36207;
    wire N__36204;
    wire N__36203;
    wire N__36200;
    wire N__36197;
    wire N__36194;
    wire N__36191;
    wire N__36190;
    wire N__36187;
    wire N__36184;
    wire N__36181;
    wire N__36174;
    wire N__36171;
    wire N__36170;
    wire N__36167;
    wire N__36164;
    wire N__36161;
    wire N__36158;
    wire N__36155;
    wire N__36154;
    wire N__36151;
    wire N__36148;
    wire N__36145;
    wire N__36138;
    wire N__36135;
    wire N__36132;
    wire N__36129;
    wire N__36126;
    wire N__36123;
    wire N__36120;
    wire N__36119;
    wire N__36118;
    wire N__36115;
    wire N__36110;
    wire N__36109;
    wire N__36104;
    wire N__36101;
    wire N__36096;
    wire N__36093;
    wire N__36092;
    wire N__36091;
    wire N__36090;
    wire N__36087;
    wire N__36086;
    wire N__36083;
    wire N__36078;
    wire N__36073;
    wire N__36072;
    wire N__36071;
    wire N__36070;
    wire N__36069;
    wire N__36066;
    wire N__36063;
    wire N__36062;
    wire N__36061;
    wire N__36058;
    wire N__36055;
    wire N__36050;
    wire N__36047;
    wire N__36044;
    wire N__36041;
    wire N__36036;
    wire N__36031;
    wire N__36028;
    wire N__36015;
    wire N__36012;
    wire N__36009;
    wire N__36006;
    wire N__36005;
    wire N__36002;
    wire N__35999;
    wire N__35994;
    wire N__35991;
    wire N__35988;
    wire N__35985;
    wire N__35982;
    wire N__35979;
    wire N__35976;
    wire N__35973;
    wire N__35970;
    wire N__35967;
    wire N__35964;
    wire N__35961;
    wire N__35958;
    wire N__35957;
    wire N__35954;
    wire N__35951;
    wire N__35950;
    wire N__35947;
    wire N__35942;
    wire N__35941;
    wire N__35940;
    wire N__35937;
    wire N__35934;
    wire N__35929;
    wire N__35926;
    wire N__35923;
    wire N__35920;
    wire N__35917;
    wire N__35914;
    wire N__35911;
    wire N__35904;
    wire N__35903;
    wire N__35902;
    wire N__35899;
    wire N__35896;
    wire N__35893;
    wire N__35892;
    wire N__35891;
    wire N__35888;
    wire N__35883;
    wire N__35878;
    wire N__35871;
    wire N__35868;
    wire N__35865;
    wire N__35862;
    wire N__35859;
    wire N__35858;
    wire N__35855;
    wire N__35852;
    wire N__35849;
    wire N__35844;
    wire N__35841;
    wire N__35838;
    wire N__35835;
    wire N__35832;
    wire N__35829;
    wire N__35828;
    wire N__35825;
    wire N__35822;
    wire N__35821;
    wire N__35820;
    wire N__35819;
    wire N__35818;
    wire N__35817;
    wire N__35814;
    wire N__35811;
    wire N__35806;
    wire N__35799;
    wire N__35790;
    wire N__35787;
    wire N__35786;
    wire N__35783;
    wire N__35780;
    wire N__35775;
    wire N__35772;
    wire N__35769;
    wire N__35766;
    wire N__35765;
    wire N__35762;
    wire N__35759;
    wire N__35758;
    wire N__35757;
    wire N__35754;
    wire N__35751;
    wire N__35750;
    wire N__35747;
    wire N__35746;
    wire N__35745;
    wire N__35744;
    wire N__35743;
    wire N__35740;
    wire N__35737;
    wire N__35734;
    wire N__35729;
    wire N__35726;
    wire N__35725;
    wire N__35724;
    wire N__35723;
    wire N__35720;
    wire N__35719;
    wire N__35716;
    wire N__35713;
    wire N__35712;
    wire N__35711;
    wire N__35708;
    wire N__35705;
    wire N__35704;
    wire N__35703;
    wire N__35702;
    wire N__35699;
    wire N__35696;
    wire N__35693;
    wire N__35690;
    wire N__35683;
    wire N__35682;
    wire N__35679;
    wire N__35676;
    wire N__35673;
    wire N__35668;
    wire N__35663;
    wire N__35660;
    wire N__35655;
    wire N__35644;
    wire N__35641;
    wire N__35622;
    wire N__35619;
    wire N__35616;
    wire N__35613;
    wire N__35610;
    wire N__35607;
    wire N__35606;
    wire N__35605;
    wire N__35602;
    wire N__35599;
    wire N__35596;
    wire N__35595;
    wire N__35590;
    wire N__35587;
    wire N__35584;
    wire N__35583;
    wire N__35582;
    wire N__35579;
    wire N__35574;
    wire N__35569;
    wire N__35566;
    wire N__35563;
    wire N__35560;
    wire N__35553;
    wire N__35552;
    wire N__35551;
    wire N__35550;
    wire N__35549;
    wire N__35546;
    wire N__35541;
    wire N__35536;
    wire N__35535;
    wire N__35534;
    wire N__35533;
    wire N__35532;
    wire N__35529;
    wire N__35526;
    wire N__35523;
    wire N__35518;
    wire N__35515;
    wire N__35512;
    wire N__35499;
    wire N__35496;
    wire N__35493;
    wire N__35492;
    wire N__35489;
    wire N__35486;
    wire N__35483;
    wire N__35480;
    wire N__35477;
    wire N__35474;
    wire N__35471;
    wire N__35468;
    wire N__35463;
    wire N__35462;
    wire N__35457;
    wire N__35454;
    wire N__35453;
    wire N__35448;
    wire N__35445;
    wire N__35442;
    wire N__35439;
    wire N__35438;
    wire N__35433;
    wire N__35430;
    wire N__35427;
    wire N__35424;
    wire N__35421;
    wire N__35420;
    wire N__35415;
    wire N__35412;
    wire N__35409;
    wire N__35406;
    wire N__35405;
    wire N__35402;
    wire N__35401;
    wire N__35398;
    wire N__35395;
    wire N__35390;
    wire N__35385;
    wire N__35384;
    wire N__35381;
    wire N__35378;
    wire N__35377;
    wire N__35374;
    wire N__35371;
    wire N__35370;
    wire N__35367;
    wire N__35364;
    wire N__35361;
    wire N__35358;
    wire N__35353;
    wire N__35346;
    wire N__35345;
    wire N__35342;
    wire N__35339;
    wire N__35336;
    wire N__35333;
    wire N__35330;
    wire N__35325;
    wire N__35324;
    wire N__35321;
    wire N__35318;
    wire N__35317;
    wire N__35314;
    wire N__35311;
    wire N__35308;
    wire N__35303;
    wire N__35298;
    wire N__35297;
    wire N__35294;
    wire N__35293;
    wire N__35292;
    wire N__35289;
    wire N__35288;
    wire N__35287;
    wire N__35284;
    wire N__35281;
    wire N__35278;
    wire N__35277;
    wire N__35276;
    wire N__35269;
    wire N__35264;
    wire N__35261;
    wire N__35258;
    wire N__35255;
    wire N__35250;
    wire N__35241;
    wire N__35238;
    wire N__35237;
    wire N__35234;
    wire N__35233;
    wire N__35230;
    wire N__35227;
    wire N__35224;
    wire N__35221;
    wire N__35214;
    wire N__35211;
    wire N__35210;
    wire N__35207;
    wire N__35204;
    wire N__35201;
    wire N__35200;
    wire N__35197;
    wire N__35194;
    wire N__35191;
    wire N__35188;
    wire N__35185;
    wire N__35178;
    wire N__35175;
    wire N__35172;
    wire N__35169;
    wire N__35166;
    wire N__35163;
    wire N__35160;
    wire N__35157;
    wire N__35154;
    wire N__35151;
    wire N__35148;
    wire N__35145;
    wire N__35142;
    wire N__35139;
    wire N__35136;
    wire N__35133;
    wire N__35130;
    wire N__35127;
    wire N__35124;
    wire N__35121;
    wire N__35120;
    wire N__35119;
    wire N__35116;
    wire N__35113;
    wire N__35110;
    wire N__35105;
    wire N__35102;
    wire N__35099;
    wire N__35094;
    wire N__35093;
    wire N__35092;
    wire N__35089;
    wire N__35084;
    wire N__35081;
    wire N__35078;
    wire N__35075;
    wire N__35074;
    wire N__35071;
    wire N__35068;
    wire N__35065;
    wire N__35062;
    wire N__35055;
    wire N__35052;
    wire N__35051;
    wire N__35050;
    wire N__35047;
    wire N__35044;
    wire N__35041;
    wire N__35034;
    wire N__35031;
    wire N__35030;
    wire N__35027;
    wire N__35026;
    wire N__35023;
    wire N__35020;
    wire N__35017;
    wire N__35010;
    wire N__35009;
    wire N__35006;
    wire N__35003;
    wire N__35000;
    wire N__34999;
    wire N__34996;
    wire N__34993;
    wire N__34990;
    wire N__34987;
    wire N__34980;
    wire N__34977;
    wire N__34974;
    wire N__34973;
    wire N__34970;
    wire N__34967;
    wire N__34962;
    wire N__34959;
    wire N__34958;
    wire N__34955;
    wire N__34952;
    wire N__34947;
    wire N__34944;
    wire N__34941;
    wire N__34938;
    wire N__34935;
    wire N__34934;
    wire N__34933;
    wire N__34930;
    wire N__34927;
    wire N__34924;
    wire N__34923;
    wire N__34920;
    wire N__34917;
    wire N__34914;
    wire N__34911;
    wire N__34908;
    wire N__34903;
    wire N__34896;
    wire N__34895;
    wire N__34894;
    wire N__34891;
    wire N__34890;
    wire N__34887;
    wire N__34884;
    wire N__34881;
    wire N__34878;
    wire N__34869;
    wire N__34866;
    wire N__34865;
    wire N__34862;
    wire N__34859;
    wire N__34856;
    wire N__34855;
    wire N__34854;
    wire N__34851;
    wire N__34848;
    wire N__34845;
    wire N__34842;
    wire N__34833;
    wire N__34832;
    wire N__34829;
    wire N__34826;
    wire N__34821;
    wire N__34820;
    wire N__34817;
    wire N__34814;
    wire N__34809;
    wire N__34806;
    wire N__34803;
    wire N__34800;
    wire N__34799;
    wire N__34798;
    wire N__34797;
    wire N__34796;
    wire N__34793;
    wire N__34790;
    wire N__34785;
    wire N__34782;
    wire N__34773;
    wire N__34772;
    wire N__34771;
    wire N__34768;
    wire N__34767;
    wire N__34766;
    wire N__34765;
    wire N__34764;
    wire N__34763;
    wire N__34760;
    wire N__34757;
    wire N__34754;
    wire N__34751;
    wire N__34744;
    wire N__34741;
    wire N__34728;
    wire N__34725;
    wire N__34724;
    wire N__34721;
    wire N__34718;
    wire N__34715;
    wire N__34714;
    wire N__34711;
    wire N__34710;
    wire N__34707;
    wire N__34704;
    wire N__34701;
    wire N__34698;
    wire N__34695;
    wire N__34692;
    wire N__34687;
    wire N__34680;
    wire N__34677;
    wire N__34674;
    wire N__34673;
    wire N__34670;
    wire N__34667;
    wire N__34664;
    wire N__34659;
    wire N__34656;
    wire N__34655;
    wire N__34652;
    wire N__34649;
    wire N__34646;
    wire N__34641;
    wire N__34638;
    wire N__34635;
    wire N__34632;
    wire N__34629;
    wire N__34628;
    wire N__34625;
    wire N__34622;
    wire N__34619;
    wire N__34614;
    wire N__34613;
    wire N__34610;
    wire N__34609;
    wire N__34608;
    wire N__34607;
    wire N__34604;
    wire N__34601;
    wire N__34596;
    wire N__34593;
    wire N__34590;
    wire N__34581;
    wire N__34578;
    wire N__34575;
    wire N__34574;
    wire N__34571;
    wire N__34568;
    wire N__34563;
    wire N__34562;
    wire N__34557;
    wire N__34554;
    wire N__34551;
    wire N__34550;
    wire N__34547;
    wire N__34544;
    wire N__34541;
    wire N__34536;
    wire N__34533;
    wire N__34530;
    wire N__34529;
    wire N__34528;
    wire N__34523;
    wire N__34522;
    wire N__34521;
    wire N__34518;
    wire N__34515;
    wire N__34512;
    wire N__34509;
    wire N__34506;
    wire N__34503;
    wire N__34500;
    wire N__34491;
    wire N__34488;
    wire N__34485;
    wire N__34484;
    wire N__34481;
    wire N__34478;
    wire N__34477;
    wire N__34476;
    wire N__34471;
    wire N__34468;
    wire N__34465;
    wire N__34462;
    wire N__34459;
    wire N__34456;
    wire N__34453;
    wire N__34446;
    wire N__34443;
    wire N__34442;
    wire N__34441;
    wire N__34438;
    wire N__34437;
    wire N__34434;
    wire N__34431;
    wire N__34428;
    wire N__34425;
    wire N__34416;
    wire N__34413;
    wire N__34410;
    wire N__34409;
    wire N__34404;
    wire N__34401;
    wire N__34398;
    wire N__34397;
    wire N__34396;
    wire N__34395;
    wire N__34392;
    wire N__34387;
    wire N__34384;
    wire N__34379;
    wire N__34376;
    wire N__34373;
    wire N__34368;
    wire N__34365;
    wire N__34364;
    wire N__34361;
    wire N__34358;
    wire N__34355;
    wire N__34350;
    wire N__34347;
    wire N__34344;
    wire N__34343;
    wire N__34340;
    wire N__34337;
    wire N__34334;
    wire N__34329;
    wire N__34326;
    wire N__34325;
    wire N__34322;
    wire N__34319;
    wire N__34318;
    wire N__34315;
    wire N__34314;
    wire N__34309;
    wire N__34306;
    wire N__34303;
    wire N__34300;
    wire N__34297;
    wire N__34294;
    wire N__34291;
    wire N__34288;
    wire N__34281;
    wire N__34278;
    wire N__34275;
    wire N__34272;
    wire N__34269;
    wire N__34266;
    wire N__34263;
    wire N__34260;
    wire N__34257;
    wire N__34254;
    wire N__34253;
    wire N__34250;
    wire N__34247;
    wire N__34244;
    wire N__34239;
    wire N__34238;
    wire N__34233;
    wire N__34230;
    wire N__34227;
    wire N__34226;
    wire N__34223;
    wire N__34220;
    wire N__34215;
    wire N__34214;
    wire N__34211;
    wire N__34208;
    wire N__34203;
    wire N__34200;
    wire N__34199;
    wire N__34196;
    wire N__34193;
    wire N__34190;
    wire N__34185;
    wire N__34184;
    wire N__34183;
    wire N__34176;
    wire N__34173;
    wire N__34172;
    wire N__34169;
    wire N__34166;
    wire N__34161;
    wire N__34160;
    wire N__34157;
    wire N__34154;
    wire N__34153;
    wire N__34150;
    wire N__34147;
    wire N__34144;
    wire N__34141;
    wire N__34138;
    wire N__34131;
    wire N__34128;
    wire N__34125;
    wire N__34122;
    wire N__34119;
    wire N__34116;
    wire N__34113;
    wire N__34112;
    wire N__34111;
    wire N__34110;
    wire N__34109;
    wire N__34108;
    wire N__34107;
    wire N__34106;
    wire N__34099;
    wire N__34088;
    wire N__34083;
    wire N__34080;
    wire N__34077;
    wire N__34074;
    wire N__34071;
    wire N__34068;
    wire N__34067;
    wire N__34064;
    wire N__34061;
    wire N__34058;
    wire N__34055;
    wire N__34050;
    wire N__34047;
    wire N__34044;
    wire N__34043;
    wire N__34038;
    wire N__34035;
    wire N__34032;
    wire N__34029;
    wire N__34026;
    wire N__34023;
    wire N__34020;
    wire N__34017;
    wire N__34014;
    wire N__34011;
    wire N__34008;
    wire N__34007;
    wire N__34002;
    wire N__33999;
    wire N__33996;
    wire N__33993;
    wire N__33990;
    wire N__33987;
    wire N__33984;
    wire N__33983;
    wire N__33980;
    wire N__33977;
    wire N__33974;
    wire N__33971;
    wire N__33966;
    wire N__33963;
    wire N__33960;
    wire N__33957;
    wire N__33954;
    wire N__33951;
    wire N__33948;
    wire N__33945;
    wire N__33944;
    wire N__33941;
    wire N__33938;
    wire N__33935;
    wire N__33930;
    wire N__33929;
    wire N__33926;
    wire N__33923;
    wire N__33920;
    wire N__33915;
    wire N__33912;
    wire N__33909;
    wire N__33906;
    wire N__33903;
    wire N__33900;
    wire N__33899;
    wire N__33896;
    wire N__33893;
    wire N__33890;
    wire N__33885;
    wire N__33882;
    wire N__33881;
    wire N__33878;
    wire N__33875;
    wire N__33872;
    wire N__33867;
    wire N__33864;
    wire N__33863;
    wire N__33860;
    wire N__33857;
    wire N__33854;
    wire N__33849;
    wire N__33846;
    wire N__33843;
    wire N__33840;
    wire N__33837;
    wire N__33834;
    wire N__33831;
    wire N__33830;
    wire N__33827;
    wire N__33824;
    wire N__33821;
    wire N__33816;
    wire N__33815;
    wire N__33812;
    wire N__33809;
    wire N__33806;
    wire N__33803;
    wire N__33798;
    wire N__33795;
    wire N__33794;
    wire N__33793;
    wire N__33790;
    wire N__33787;
    wire N__33784;
    wire N__33777;
    wire N__33774;
    wire N__33771;
    wire N__33768;
    wire N__33765;
    wire N__33764;
    wire N__33761;
    wire N__33758;
    wire N__33755;
    wire N__33752;
    wire N__33747;
    wire N__33744;
    wire N__33741;
    wire N__33740;
    wire N__33739;
    wire N__33736;
    wire N__33733;
    wire N__33732;
    wire N__33729;
    wire N__33728;
    wire N__33725;
    wire N__33720;
    wire N__33715;
    wire N__33708;
    wire N__33705;
    wire N__33702;
    wire N__33699;
    wire N__33698;
    wire N__33695;
    wire N__33692;
    wire N__33687;
    wire N__33684;
    wire N__33681;
    wire N__33678;
    wire N__33675;
    wire N__33672;
    wire N__33669;
    wire N__33666;
    wire N__33663;
    wire N__33660;
    wire N__33657;
    wire N__33656;
    wire N__33655;
    wire N__33652;
    wire N__33651;
    wire N__33648;
    wire N__33643;
    wire N__33640;
    wire N__33637;
    wire N__33634;
    wire N__33631;
    wire N__33628;
    wire N__33625;
    wire N__33618;
    wire N__33615;
    wire N__33612;
    wire N__33609;
    wire N__33606;
    wire N__33603;
    wire N__33600;
    wire N__33597;
    wire N__33594;
    wire N__33591;
    wire N__33588;
    wire N__33585;
    wire N__33582;
    wire N__33579;
    wire N__33576;
    wire N__33573;
    wire N__33570;
    wire N__33567;
    wire N__33564;
    wire N__33561;
    wire N__33558;
    wire N__33555;
    wire N__33554;
    wire N__33553;
    wire N__33550;
    wire N__33547;
    wire N__33544;
    wire N__33537;
    wire N__33536;
    wire N__33535;
    wire N__33534;
    wire N__33531;
    wire N__33528;
    wire N__33523;
    wire N__33522;
    wire N__33521;
    wire N__33520;
    wire N__33519;
    wire N__33516;
    wire N__33511;
    wire N__33502;
    wire N__33499;
    wire N__33494;
    wire N__33489;
    wire N__33488;
    wire N__33487;
    wire N__33484;
    wire N__33479;
    wire N__33476;
    wire N__33471;
    wire N__33470;
    wire N__33469;
    wire N__33466;
    wire N__33463;
    wire N__33460;
    wire N__33455;
    wire N__33452;
    wire N__33449;
    wire N__33444;
    wire N__33441;
    wire N__33438;
    wire N__33437;
    wire N__33436;
    wire N__33433;
    wire N__33430;
    wire N__33427;
    wire N__33422;
    wire N__33417;
    wire N__33416;
    wire N__33413;
    wire N__33412;
    wire N__33409;
    wire N__33406;
    wire N__33403;
    wire N__33400;
    wire N__33397;
    wire N__33390;
    wire N__33387;
    wire N__33384;
    wire N__33383;
    wire N__33382;
    wire N__33381;
    wire N__33380;
    wire N__33375;
    wire N__33372;
    wire N__33367;
    wire N__33360;
    wire N__33359;
    wire N__33356;
    wire N__33355;
    wire N__33354;
    wire N__33351;
    wire N__33348;
    wire N__33343;
    wire N__33336;
    wire N__33333;
    wire N__33332;
    wire N__33329;
    wire N__33326;
    wire N__33323;
    wire N__33322;
    wire N__33319;
    wire N__33316;
    wire N__33313;
    wire N__33306;
    wire N__33303;
    wire N__33300;
    wire N__33297;
    wire N__33294;
    wire N__33291;
    wire N__33290;
    wire N__33287;
    wire N__33284;
    wire N__33281;
    wire N__33280;
    wire N__33277;
    wire N__33274;
    wire N__33271;
    wire N__33264;
    wire N__33261;
    wire N__33258;
    wire N__33255;
    wire N__33252;
    wire N__33251;
    wire N__33250;
    wire N__33249;
    wire N__33248;
    wire N__33247;
    wire N__33246;
    wire N__33243;
    wire N__33240;
    wire N__33237;
    wire N__33236;
    wire N__33235;
    wire N__33234;
    wire N__33233;
    wire N__33232;
    wire N__33229;
    wire N__33226;
    wire N__33225;
    wire N__33224;
    wire N__33223;
    wire N__33222;
    wire N__33221;
    wire N__33220;
    wire N__33219;
    wire N__33218;
    wire N__33215;
    wire N__33212;
    wire N__33207;
    wire N__33204;
    wire N__33201;
    wire N__33198;
    wire N__33197;
    wire N__33194;
    wire N__33191;
    wire N__33188;
    wire N__33187;
    wire N__33186;
    wire N__33185;
    wire N__33184;
    wire N__33179;
    wire N__33176;
    wire N__33173;
    wire N__33170;
    wire N__33167;
    wire N__33164;
    wire N__33161;
    wire N__33160;
    wire N__33159;
    wire N__33156;
    wire N__33153;
    wire N__33152;
    wire N__33151;
    wire N__33150;
    wire N__33149;
    wire N__33148;
    wire N__33143;
    wire N__33134;
    wire N__33131;
    wire N__33124;
    wire N__33121;
    wire N__33118;
    wire N__33115;
    wire N__33112;
    wire N__33099;
    wire N__33096;
    wire N__33093;
    wire N__33090;
    wire N__33085;
    wire N__33082;
    wire N__33079;
    wire N__33076;
    wire N__33073;
    wire N__33070;
    wire N__33063;
    wire N__33052;
    wire N__33045;
    wire N__33040;
    wire N__33039;
    wire N__33028;
    wire N__33025;
    wire N__33020;
    wire N__33017;
    wire N__33014;
    wire N__33013;
    wire N__33012;
    wire N__33011;
    wire N__33008;
    wire N__33005;
    wire N__33002;
    wire N__32999;
    wire N__32996;
    wire N__32993;
    wire N__32990;
    wire N__32987;
    wire N__32970;
    wire N__32967;
    wire N__32964;
    wire N__32961;
    wire N__32958;
    wire N__32955;
    wire N__32952;
    wire N__32949;
    wire N__32946;
    wire N__32943;
    wire N__32940;
    wire N__32937;
    wire N__32936;
    wire N__32933;
    wire N__32930;
    wire N__32927;
    wire N__32922;
    wire N__32921;
    wire N__32920;
    wire N__32917;
    wire N__32916;
    wire N__32911;
    wire N__32908;
    wire N__32905;
    wire N__32898;
    wire N__32895;
    wire N__32892;
    wire N__32889;
    wire N__32888;
    wire N__32885;
    wire N__32884;
    wire N__32881;
    wire N__32880;
    wire N__32877;
    wire N__32874;
    wire N__32873;
    wire N__32872;
    wire N__32869;
    wire N__32866;
    wire N__32865;
    wire N__32862;
    wire N__32857;
    wire N__32854;
    wire N__32849;
    wire N__32846;
    wire N__32841;
    wire N__32838;
    wire N__32833;
    wire N__32830;
    wire N__32827;
    wire N__32824;
    wire N__32819;
    wire N__32816;
    wire N__32811;
    wire N__32810;
    wire N__32807;
    wire N__32804;
    wire N__32801;
    wire N__32798;
    wire N__32795;
    wire N__32792;
    wire N__32791;
    wire N__32788;
    wire N__32785;
    wire N__32782;
    wire N__32779;
    wire N__32774;
    wire N__32769;
    wire N__32766;
    wire N__32765;
    wire N__32762;
    wire N__32759;
    wire N__32756;
    wire N__32751;
    wire N__32750;
    wire N__32749;
    wire N__32746;
    wire N__32745;
    wire N__32742;
    wire N__32739;
    wire N__32736;
    wire N__32733;
    wire N__32724;
    wire N__32721;
    wire N__32718;
    wire N__32715;
    wire N__32712;
    wire N__32709;
    wire N__32708;
    wire N__32707;
    wire N__32706;
    wire N__32703;
    wire N__32702;
    wire N__32697;
    wire N__32696;
    wire N__32695;
    wire N__32692;
    wire N__32687;
    wire N__32684;
    wire N__32681;
    wire N__32680;
    wire N__32677;
    wire N__32674;
    wire N__32671;
    wire N__32668;
    wire N__32665;
    wire N__32660;
    wire N__32655;
    wire N__32652;
    wire N__32647;
    wire N__32644;
    wire N__32641;
    wire N__32640;
    wire N__32637;
    wire N__32634;
    wire N__32631;
    wire N__32628;
    wire N__32619;
    wire N__32618;
    wire N__32615;
    wire N__32612;
    wire N__32607;
    wire N__32604;
    wire N__32601;
    wire N__32600;
    wire N__32597;
    wire N__32594;
    wire N__32589;
    wire N__32586;
    wire N__32583;
    wire N__32580;
    wire N__32577;
    wire N__32574;
    wire N__32571;
    wire N__32568;
    wire N__32565;
    wire N__32564;
    wire N__32563;
    wire N__32562;
    wire N__32561;
    wire N__32560;
    wire N__32559;
    wire N__32556;
    wire N__32553;
    wire N__32546;
    wire N__32541;
    wire N__32532;
    wire N__32531;
    wire N__32528;
    wire N__32525;
    wire N__32522;
    wire N__32517;
    wire N__32514;
    wire N__32511;
    wire N__32508;
    wire N__32507;
    wire N__32506;
    wire N__32503;
    wire N__32498;
    wire N__32493;
    wire N__32492;
    wire N__32489;
    wire N__32486;
    wire N__32483;
    wire N__32478;
    wire N__32475;
    wire N__32474;
    wire N__32471;
    wire N__32468;
    wire N__32463;
    wire N__32462;
    wire N__32461;
    wire N__32460;
    wire N__32459;
    wire N__32458;
    wire N__32455;
    wire N__32448;
    wire N__32447;
    wire N__32446;
    wire N__32445;
    wire N__32444;
    wire N__32443;
    wire N__32442;
    wire N__32441;
    wire N__32436;
    wire N__32433;
    wire N__32430;
    wire N__32425;
    wire N__32424;
    wire N__32423;
    wire N__32418;
    wire N__32417;
    wire N__32416;
    wire N__32415;
    wire N__32414;
    wire N__32413;
    wire N__32412;
    wire N__32405;
    wire N__32402;
    wire N__32395;
    wire N__32392;
    wire N__32389;
    wire N__32388;
    wire N__32385;
    wire N__32378;
    wire N__32371;
    wire N__32370;
    wire N__32369;
    wire N__32364;
    wire N__32363;
    wire N__32362;
    wire N__32359;
    wire N__32354;
    wire N__32351;
    wire N__32348;
    wire N__32343;
    wire N__32338;
    wire N__32335;
    wire N__32334;
    wire N__32333;
    wire N__32330;
    wire N__32327;
    wire N__32324;
    wire N__32313;
    wire N__32310;
    wire N__32307;
    wire N__32304;
    wire N__32289;
    wire N__32288;
    wire N__32287;
    wire N__32284;
    wire N__32281;
    wire N__32278;
    wire N__32277;
    wire N__32276;
    wire N__32275;
    wire N__32268;
    wire N__32265;
    wire N__32262;
    wire N__32261;
    wire N__32260;
    wire N__32257;
    wire N__32254;
    wire N__32251;
    wire N__32248;
    wire N__32247;
    wire N__32244;
    wire N__32241;
    wire N__32236;
    wire N__32235;
    wire N__32234;
    wire N__32229;
    wire N__32226;
    wire N__32225;
    wire N__32218;
    wire N__32215;
    wire N__32212;
    wire N__32209;
    wire N__32206;
    wire N__32203;
    wire N__32198;
    wire N__32187;
    wire N__32184;
    wire N__32181;
    wire N__32178;
    wire N__32175;
    wire N__32174;
    wire N__32173;
    wire N__32172;
    wire N__32171;
    wire N__32170;
    wire N__32169;
    wire N__32168;
    wire N__32167;
    wire N__32162;
    wire N__32157;
    wire N__32154;
    wire N__32153;
    wire N__32150;
    wire N__32149;
    wire N__32148;
    wire N__32147;
    wire N__32146;
    wire N__32143;
    wire N__32142;
    wire N__32141;
    wire N__32136;
    wire N__32133;
    wire N__32128;
    wire N__32123;
    wire N__32120;
    wire N__32113;
    wire N__32110;
    wire N__32109;
    wire N__32104;
    wire N__32101;
    wire N__32096;
    wire N__32087;
    wire N__32084;
    wire N__32077;
    wire N__32072;
    wire N__32071;
    wire N__32070;
    wire N__32069;
    wire N__32066;
    wire N__32063;
    wire N__32056;
    wire N__32049;
    wire N__32046;
    wire N__32043;
    wire N__32040;
    wire N__32037;
    wire N__32034;
    wire N__32031;
    wire N__32030;
    wire N__32027;
    wire N__32024;
    wire N__32021;
    wire N__32016;
    wire N__32013;
    wire N__32012;
    wire N__32009;
    wire N__32006;
    wire N__32003;
    wire N__32000;
    wire N__31995;
    wire N__31992;
    wire N__31989;
    wire N__31986;
    wire N__31983;
    wire N__31980;
    wire N__31977;
    wire N__31974;
    wire N__31973;
    wire N__31970;
    wire N__31967;
    wire N__31964;
    wire N__31961;
    wire N__31956;
    wire N__31953;
    wire N__31952;
    wire N__31949;
    wire N__31946;
    wire N__31943;
    wire N__31940;
    wire N__31939;
    wire N__31938;
    wire N__31937;
    wire N__31934;
    wire N__31933;
    wire N__31930;
    wire N__31927;
    wire N__31922;
    wire N__31919;
    wire N__31916;
    wire N__31913;
    wire N__31908;
    wire N__31899;
    wire N__31896;
    wire N__31895;
    wire N__31892;
    wire N__31891;
    wire N__31890;
    wire N__31887;
    wire N__31884;
    wire N__31879;
    wire N__31876;
    wire N__31869;
    wire N__31868;
    wire N__31867;
    wire N__31866;
    wire N__31863;
    wire N__31854;
    wire N__31853;
    wire N__31852;
    wire N__31851;
    wire N__31850;
    wire N__31849;
    wire N__31848;
    wire N__31845;
    wire N__31842;
    wire N__31839;
    wire N__31836;
    wire N__31829;
    wire N__31826;
    wire N__31823;
    wire N__31818;
    wire N__31815;
    wire N__31810;
    wire N__31805;
    wire N__31800;
    wire N__31797;
    wire N__31794;
    wire N__31791;
    wire N__31788;
    wire N__31785;
    wire N__31782;
    wire N__31781;
    wire N__31776;
    wire N__31775;
    wire N__31774;
    wire N__31771;
    wire N__31768;
    wire N__31767;
    wire N__31764;
    wire N__31761;
    wire N__31758;
    wire N__31755;
    wire N__31752;
    wire N__31749;
    wire N__31746;
    wire N__31737;
    wire N__31736;
    wire N__31735;
    wire N__31730;
    wire N__31727;
    wire N__31726;
    wire N__31723;
    wire N__31720;
    wire N__31719;
    wire N__31716;
    wire N__31713;
    wire N__31710;
    wire N__31707;
    wire N__31698;
    wire N__31695;
    wire N__31692;
    wire N__31691;
    wire N__31686;
    wire N__31683;
    wire N__31680;
    wire N__31677;
    wire N__31676;
    wire N__31675;
    wire N__31674;
    wire N__31671;
    wire N__31668;
    wire N__31665;
    wire N__31662;
    wire N__31659;
    wire N__31656;
    wire N__31655;
    wire N__31652;
    wire N__31649;
    wire N__31646;
    wire N__31643;
    wire N__31640;
    wire N__31633;
    wire N__31626;
    wire N__31623;
    wire N__31622;
    wire N__31619;
    wire N__31618;
    wire N__31615;
    wire N__31614;
    wire N__31611;
    wire N__31608;
    wire N__31605;
    wire N__31602;
    wire N__31597;
    wire N__31596;
    wire N__31593;
    wire N__31590;
    wire N__31587;
    wire N__31584;
    wire N__31581;
    wire N__31578;
    wire N__31569;
    wire N__31566;
    wire N__31565;
    wire N__31564;
    wire N__31563;
    wire N__31560;
    wire N__31557;
    wire N__31554;
    wire N__31551;
    wire N__31548;
    wire N__31545;
    wire N__31544;
    wire N__31539;
    wire N__31536;
    wire N__31533;
    wire N__31530;
    wire N__31525;
    wire N__31518;
    wire N__31515;
    wire N__31514;
    wire N__31513;
    wire N__31510;
    wire N__31507;
    wire N__31506;
    wire N__31503;
    wire N__31500;
    wire N__31497;
    wire N__31494;
    wire N__31491;
    wire N__31488;
    wire N__31483;
    wire N__31482;
    wire N__31479;
    wire N__31474;
    wire N__31471;
    wire N__31468;
    wire N__31461;
    wire N__31458;
    wire N__31455;
    wire N__31454;
    wire N__31453;
    wire N__31450;
    wire N__31449;
    wire N__31446;
    wire N__31443;
    wire N__31440;
    wire N__31437;
    wire N__31434;
    wire N__31431;
    wire N__31430;
    wire N__31425;
    wire N__31422;
    wire N__31419;
    wire N__31416;
    wire N__31411;
    wire N__31404;
    wire N__31401;
    wire N__31400;
    wire N__31399;
    wire N__31396;
    wire N__31393;
    wire N__31392;
    wire N__31389;
    wire N__31386;
    wire N__31383;
    wire N__31380;
    wire N__31377;
    wire N__31376;
    wire N__31373;
    wire N__31368;
    wire N__31365;
    wire N__31362;
    wire N__31357;
    wire N__31354;
    wire N__31347;
    wire N__31344;
    wire N__31341;
    wire N__31338;
    wire N__31335;
    wire N__31334;
    wire N__31331;
    wire N__31328;
    wire N__31325;
    wire N__31320;
    wire N__31319;
    wire N__31316;
    wire N__31313;
    wire N__31310;
    wire N__31307;
    wire N__31302;
    wire N__31301;
    wire N__31298;
    wire N__31295;
    wire N__31292;
    wire N__31287;
    wire N__31286;
    wire N__31283;
    wire N__31280;
    wire N__31277;
    wire N__31272;
    wire N__31269;
    wire N__31268;
    wire N__31265;
    wire N__31264;
    wire N__31263;
    wire N__31260;
    wire N__31257;
    wire N__31254;
    wire N__31251;
    wire N__31248;
    wire N__31245;
    wire N__31242;
    wire N__31239;
    wire N__31238;
    wire N__31235;
    wire N__31232;
    wire N__31227;
    wire N__31224;
    wire N__31221;
    wire N__31212;
    wire N__31209;
    wire N__31208;
    wire N__31205;
    wire N__31202;
    wire N__31201;
    wire N__31198;
    wire N__31195;
    wire N__31194;
    wire N__31191;
    wire N__31188;
    wire N__31185;
    wire N__31182;
    wire N__31181;
    wire N__31178;
    wire N__31171;
    wire N__31168;
    wire N__31165;
    wire N__31158;
    wire N__31155;
    wire N__31154;
    wire N__31151;
    wire N__31150;
    wire N__31149;
    wire N__31146;
    wire N__31143;
    wire N__31140;
    wire N__31137;
    wire N__31134;
    wire N__31131;
    wire N__31128;
    wire N__31127;
    wire N__31124;
    wire N__31121;
    wire N__31118;
    wire N__31115;
    wire N__31112;
    wire N__31107;
    wire N__31098;
    wire N__31095;
    wire N__31094;
    wire N__31091;
    wire N__31090;
    wire N__31089;
    wire N__31086;
    wire N__31083;
    wire N__31080;
    wire N__31077;
    wire N__31074;
    wire N__31071;
    wire N__31068;
    wire N__31065;
    wire N__31064;
    wire N__31061;
    wire N__31058;
    wire N__31055;
    wire N__31052;
    wire N__31049;
    wire N__31046;
    wire N__31035;
    wire N__31032;
    wire N__31031;
    wire N__31030;
    wire N__31027;
    wire N__31026;
    wire N__31023;
    wire N__31020;
    wire N__31017;
    wire N__31014;
    wire N__31011;
    wire N__31008;
    wire N__31003;
    wire N__31002;
    wire N__30999;
    wire N__30996;
    wire N__30993;
    wire N__30990;
    wire N__30987;
    wire N__30978;
    wire N__30975;
    wire N__30974;
    wire N__30971;
    wire N__30970;
    wire N__30967;
    wire N__30964;
    wire N__30961;
    wire N__30960;
    wire N__30957;
    wire N__30952;
    wire N__30949;
    wire N__30948;
    wire N__30945;
    wire N__30942;
    wire N__30939;
    wire N__30936;
    wire N__30933;
    wire N__30924;
    wire N__30921;
    wire N__30920;
    wire N__30919;
    wire N__30916;
    wire N__30915;
    wire N__30912;
    wire N__30909;
    wire N__30906;
    wire N__30903;
    wire N__30900;
    wire N__30899;
    wire N__30896;
    wire N__30891;
    wire N__30888;
    wire N__30885;
    wire N__30878;
    wire N__30873;
    wire N__30870;
    wire N__30867;
    wire N__30864;
    wire N__30863;
    wire N__30860;
    wire N__30857;
    wire N__30854;
    wire N__30851;
    wire N__30846;
    wire N__30843;
    wire N__30842;
    wire N__30839;
    wire N__30838;
    wire N__30835;
    wire N__30834;
    wire N__30831;
    wire N__30828;
    wire N__30825;
    wire N__30822;
    wire N__30819;
    wire N__30816;
    wire N__30811;
    wire N__30810;
    wire N__30807;
    wire N__30804;
    wire N__30801;
    wire N__30798;
    wire N__30793;
    wire N__30786;
    wire N__30783;
    wire N__30782;
    wire N__30781;
    wire N__30780;
    wire N__30779;
    wire N__30776;
    wire N__30773;
    wire N__30770;
    wire N__30767;
    wire N__30764;
    wire N__30761;
    wire N__30758;
    wire N__30755;
    wire N__30752;
    wire N__30751;
    wire N__30748;
    wire N__30743;
    wire N__30740;
    wire N__30737;
    wire N__30734;
    wire N__30731;
    wire N__30720;
    wire N__30717;
    wire N__30716;
    wire N__30713;
    wire N__30710;
    wire N__30709;
    wire N__30708;
    wire N__30707;
    wire N__30704;
    wire N__30701;
    wire N__30698;
    wire N__30695;
    wire N__30692;
    wire N__30689;
    wire N__30682;
    wire N__30681;
    wire N__30678;
    wire N__30673;
    wire N__30670;
    wire N__30667;
    wire N__30660;
    wire N__30657;
    wire N__30656;
    wire N__30655;
    wire N__30650;
    wire N__30647;
    wire N__30646;
    wire N__30645;
    wire N__30642;
    wire N__30639;
    wire N__30636;
    wire N__30633;
    wire N__30630;
    wire N__30629;
    wire N__30626;
    wire N__30621;
    wire N__30618;
    wire N__30615;
    wire N__30612;
    wire N__30603;
    wire N__30600;
    wire N__30599;
    wire N__30598;
    wire N__30595;
    wire N__30594;
    wire N__30591;
    wire N__30588;
    wire N__30585;
    wire N__30584;
    wire N__30581;
    wire N__30578;
    wire N__30575;
    wire N__30574;
    wire N__30571;
    wire N__30568;
    wire N__30565;
    wire N__30562;
    wire N__30559;
    wire N__30556;
    wire N__30553;
    wire N__30540;
    wire N__30537;
    wire N__30536;
    wire N__30535;
    wire N__30534;
    wire N__30533;
    wire N__30530;
    wire N__30527;
    wire N__30524;
    wire N__30521;
    wire N__30518;
    wire N__30515;
    wire N__30512;
    wire N__30509;
    wire N__30506;
    wire N__30503;
    wire N__30502;
    wire N__30497;
    wire N__30494;
    wire N__30491;
    wire N__30488;
    wire N__30485;
    wire N__30480;
    wire N__30471;
    wire N__30468;
    wire N__30467;
    wire N__30466;
    wire N__30465;
    wire N__30462;
    wire N__30459;
    wire N__30454;
    wire N__30451;
    wire N__30448;
    wire N__30447;
    wire N__30446;
    wire N__30443;
    wire N__30440;
    wire N__30437;
    wire N__30434;
    wire N__30431;
    wire N__30426;
    wire N__30417;
    wire N__30414;
    wire N__30413;
    wire N__30410;
    wire N__30407;
    wire N__30406;
    wire N__30405;
    wire N__30402;
    wire N__30399;
    wire N__30396;
    wire N__30393;
    wire N__30392;
    wire N__30389;
    wire N__30384;
    wire N__30381;
    wire N__30378;
    wire N__30375;
    wire N__30366;
    wire N__30363;
    wire N__30360;
    wire N__30359;
    wire N__30356;
    wire N__30355;
    wire N__30352;
    wire N__30351;
    wire N__30348;
    wire N__30345;
    wire N__30342;
    wire N__30339;
    wire N__30336;
    wire N__30333;
    wire N__30330;
    wire N__30329;
    wire N__30326;
    wire N__30321;
    wire N__30318;
    wire N__30315;
    wire N__30310;
    wire N__30303;
    wire N__30300;
    wire N__30299;
    wire N__30296;
    wire N__30293;
    wire N__30290;
    wire N__30287;
    wire N__30282;
    wire N__30279;
    wire N__30278;
    wire N__30275;
    wire N__30274;
    wire N__30271;
    wire N__30268;
    wire N__30265;
    wire N__30264;
    wire N__30261;
    wire N__30258;
    wire N__30257;
    wire N__30254;
    wire N__30251;
    wire N__30250;
    wire N__30247;
    wire N__30244;
    wire N__30241;
    wire N__30236;
    wire N__30233;
    wire N__30228;
    wire N__30219;
    wire N__30216;
    wire N__30215;
    wire N__30212;
    wire N__30211;
    wire N__30210;
    wire N__30209;
    wire N__30206;
    wire N__30205;
    wire N__30202;
    wire N__30197;
    wire N__30194;
    wire N__30191;
    wire N__30188;
    wire N__30185;
    wire N__30174;
    wire N__30171;
    wire N__30170;
    wire N__30169;
    wire N__30166;
    wire N__30163;
    wire N__30162;
    wire N__30159;
    wire N__30158;
    wire N__30153;
    wire N__30150;
    wire N__30147;
    wire N__30144;
    wire N__30143;
    wire N__30140;
    wire N__30137;
    wire N__30134;
    wire N__30131;
    wire N__30128;
    wire N__30123;
    wire N__30114;
    wire N__30111;
    wire N__30110;
    wire N__30109;
    wire N__30106;
    wire N__30105;
    wire N__30104;
    wire N__30101;
    wire N__30098;
    wire N__30095;
    wire N__30092;
    wire N__30089;
    wire N__30088;
    wire N__30083;
    wire N__30080;
    wire N__30077;
    wire N__30074;
    wire N__30071;
    wire N__30066;
    wire N__30057;
    wire N__30054;
    wire N__30053;
    wire N__30050;
    wire N__30049;
    wire N__30046;
    wire N__30043;
    wire N__30040;
    wire N__30039;
    wire N__30036;
    wire N__30033;
    wire N__30032;
    wire N__30031;
    wire N__30028;
    wire N__30025;
    wire N__30022;
    wire N__30019;
    wire N__30016;
    wire N__30013;
    wire N__30006;
    wire N__29997;
    wire N__29994;
    wire N__29993;
    wire N__29992;
    wire N__29991;
    wire N__29988;
    wire N__29985;
    wire N__29982;
    wire N__29979;
    wire N__29976;
    wire N__29973;
    wire N__29970;
    wire N__29967;
    wire N__29966;
    wire N__29965;
    wire N__29962;
    wire N__29959;
    wire N__29954;
    wire N__29951;
    wire N__29948;
    wire N__29945;
    wire N__29934;
    wire N__29931;
    wire N__29930;
    wire N__29929;
    wire N__29926;
    wire N__29923;
    wire N__29920;
    wire N__29917;
    wire N__29916;
    wire N__29913;
    wire N__29912;
    wire N__29907;
    wire N__29904;
    wire N__29903;
    wire N__29900;
    wire N__29897;
    wire N__29892;
    wire N__29889;
    wire N__29886;
    wire N__29877;
    wire N__29874;
    wire N__29873;
    wire N__29872;
    wire N__29869;
    wire N__29866;
    wire N__29863;
    wire N__29862;
    wire N__29861;
    wire N__29858;
    wire N__29855;
    wire N__29852;
    wire N__29847;
    wire N__29846;
    wire N__29843;
    wire N__29840;
    wire N__29835;
    wire N__29832;
    wire N__29827;
    wire N__29820;
    wire N__29817;
    wire N__29816;
    wire N__29813;
    wire N__29812;
    wire N__29811;
    wire N__29810;
    wire N__29807;
    wire N__29804;
    wire N__29799;
    wire N__29796;
    wire N__29793;
    wire N__29790;
    wire N__29787;
    wire N__29784;
    wire N__29783;
    wire N__29780;
    wire N__29775;
    wire N__29772;
    wire N__29769;
    wire N__29766;
    wire N__29757;
    wire N__29754;
    wire N__29753;
    wire N__29750;
    wire N__29747;
    wire N__29744;
    wire N__29741;
    wire N__29736;
    wire N__29733;
    wire N__29732;
    wire N__29731;
    wire N__29730;
    wire N__29727;
    wire N__29724;
    wire N__29719;
    wire N__29712;
    wire N__29711;
    wire N__29710;
    wire N__29707;
    wire N__29704;
    wire N__29701;
    wire N__29698;
    wire N__29695;
    wire N__29692;
    wire N__29689;
    wire N__29686;
    wire N__29683;
    wire N__29680;
    wire N__29679;
    wire N__29676;
    wire N__29673;
    wire N__29670;
    wire N__29667;
    wire N__29662;
    wire N__29655;
    wire N__29652;
    wire N__29651;
    wire N__29648;
    wire N__29647;
    wire N__29646;
    wire N__29643;
    wire N__29640;
    wire N__29637;
    wire N__29634;
    wire N__29627;
    wire N__29622;
    wire N__29619;
    wire N__29616;
    wire N__29613;
    wire N__29610;
    wire N__29609;
    wire N__29608;
    wire N__29605;
    wire N__29602;
    wire N__29599;
    wire N__29596;
    wire N__29593;
    wire N__29586;
    wire N__29583;
    wire N__29580;
    wire N__29577;
    wire N__29574;
    wire N__29571;
    wire N__29568;
    wire N__29565;
    wire N__29564;
    wire N__29561;
    wire N__29560;
    wire N__29559;
    wire N__29558;
    wire N__29555;
    wire N__29552;
    wire N__29549;
    wire N__29546;
    wire N__29543;
    wire N__29542;
    wire N__29539;
    wire N__29534;
    wire N__29529;
    wire N__29526;
    wire N__29523;
    wire N__29520;
    wire N__29517;
    wire N__29508;
    wire N__29505;
    wire N__29502;
    wire N__29499;
    wire N__29496;
    wire N__29493;
    wire N__29490;
    wire N__29487;
    wire N__29484;
    wire N__29481;
    wire N__29478;
    wire N__29475;
    wire N__29472;
    wire N__29469;
    wire N__29466;
    wire N__29463;
    wire N__29460;
    wire N__29459;
    wire N__29458;
    wire N__29455;
    wire N__29454;
    wire N__29453;
    wire N__29450;
    wire N__29447;
    wire N__29444;
    wire N__29441;
    wire N__29438;
    wire N__29435;
    wire N__29432;
    wire N__29431;
    wire N__29428;
    wire N__29425;
    wire N__29420;
    wire N__29417;
    wire N__29414;
    wire N__29411;
    wire N__29400;
    wire N__29397;
    wire N__29394;
    wire N__29393;
    wire N__29392;
    wire N__29391;
    wire N__29388;
    wire N__29381;
    wire N__29376;
    wire N__29375;
    wire N__29372;
    wire N__29369;
    wire N__29366;
    wire N__29361;
    wire N__29358;
    wire N__29355;
    wire N__29352;
    wire N__29349;
    wire N__29346;
    wire N__29343;
    wire N__29340;
    wire N__29337;
    wire N__29334;
    wire N__29333;
    wire N__29330;
    wire N__29329;
    wire N__29328;
    wire N__29325;
    wire N__29322;
    wire N__29317;
    wire N__29310;
    wire N__29307;
    wire N__29304;
    wire N__29301;
    wire N__29300;
    wire N__29297;
    wire N__29294;
    wire N__29291;
    wire N__29288;
    wire N__29285;
    wire N__29280;
    wire N__29279;
    wire N__29278;
    wire N__29275;
    wire N__29270;
    wire N__29265;
    wire N__29262;
    wire N__29259;
    wire N__29256;
    wire N__29253;
    wire N__29252;
    wire N__29249;
    wire N__29246;
    wire N__29241;
    wire N__29240;
    wire N__29237;
    wire N__29234;
    wire N__29233;
    wire N__29232;
    wire N__29229;
    wire N__29226;
    wire N__29221;
    wire N__29214;
    wire N__29213;
    wire N__29212;
    wire N__29211;
    wire N__29206;
    wire N__29203;
    wire N__29200;
    wire N__29193;
    wire N__29190;
    wire N__29187;
    wire N__29184;
    wire N__29181;
    wire N__29180;
    wire N__29177;
    wire N__29176;
    wire N__29175;
    wire N__29172;
    wire N__29169;
    wire N__29166;
    wire N__29163;
    wire N__29154;
    wire N__29153;
    wire N__29150;
    wire N__29149;
    wire N__29144;
    wire N__29141;
    wire N__29140;
    wire N__29135;
    wire N__29132;
    wire N__29129;
    wire N__29124;
    wire N__29121;
    wire N__29118;
    wire N__29115;
    wire N__29112;
    wire N__29109;
    wire N__29108;
    wire N__29105;
    wire N__29102;
    wire N__29097;
    wire N__29094;
    wire N__29091;
    wire N__29088;
    wire N__29085;
    wire N__29082;
    wire N__29079;
    wire N__29076;
    wire N__29073;
    wire N__29070;
    wire N__29067;
    wire N__29066;
    wire N__29063;
    wire N__29060;
    wire N__29059;
    wire N__29058;
    wire N__29057;
    wire N__29056;
    wire N__29055;
    wire N__29054;
    wire N__29053;
    wire N__29052;
    wire N__29051;
    wire N__29050;
    wire N__29049;
    wire N__29048;
    wire N__29047;
    wire N__29044;
    wire N__29041;
    wire N__29036;
    wire N__29033;
    wire N__29028;
    wire N__29025;
    wire N__29024;
    wire N__29023;
    wire N__29022;
    wire N__29019;
    wire N__29014;
    wire N__29009;
    wire N__29008;
    wire N__29007;
    wire N__29006;
    wire N__29005;
    wire N__29004;
    wire N__29003;
    wire N__29000;
    wire N__28999;
    wire N__28998;
    wire N__28997;
    wire N__28994;
    wire N__28989;
    wire N__28986;
    wire N__28981;
    wire N__28978;
    wire N__28973;
    wire N__28972;
    wire N__28971;
    wire N__28970;
    wire N__28969;
    wire N__28968;
    wire N__28967;
    wire N__28966;
    wire N__28963;
    wire N__28962;
    wire N__28961;
    wire N__28960;
    wire N__28959;
    wire N__28954;
    wire N__28951;
    wire N__28944;
    wire N__28939;
    wire N__28938;
    wire N__28935;
    wire N__28934;
    wire N__28933;
    wire N__28932;
    wire N__28929;
    wire N__28926;
    wire N__28925;
    wire N__28924;
    wire N__28923;
    wire N__28920;
    wire N__28917;
    wire N__28914;
    wire N__28911;
    wire N__28902;
    wire N__28901;
    wire N__28896;
    wire N__28893;
    wire N__28892;
    wire N__28891;
    wire N__28888;
    wire N__28881;
    wire N__28878;
    wire N__28873;
    wire N__28870;
    wire N__28867;
    wire N__28862;
    wire N__28857;
    wire N__28854;
    wire N__28851;
    wire N__28846;
    wire N__28843;
    wire N__28838;
    wire N__28831;
    wire N__28826;
    wire N__28819;
    wire N__28818;
    wire N__28817;
    wire N__28816;
    wire N__28813;
    wire N__28808;
    wire N__28803;
    wire N__28794;
    wire N__28791;
    wire N__28784;
    wire N__28783;
    wire N__28776;
    wire N__28773;
    wire N__28764;
    wire N__28757;
    wire N__28748;
    wire N__28743;
    wire N__28740;
    wire N__28735;
    wire N__28732;
    wire N__28725;
    wire N__28716;
    wire N__28713;
    wire N__28710;
    wire N__28707;
    wire N__28704;
    wire N__28701;
    wire N__28700;
    wire N__28699;
    wire N__28696;
    wire N__28695;
    wire N__28694;
    wire N__28689;
    wire N__28686;
    wire N__28685;
    wire N__28684;
    wire N__28683;
    wire N__28680;
    wire N__28677;
    wire N__28676;
    wire N__28675;
    wire N__28672;
    wire N__28669;
    wire N__28664;
    wire N__28663;
    wire N__28662;
    wire N__28661;
    wire N__28660;
    wire N__28659;
    wire N__28656;
    wire N__28655;
    wire N__28654;
    wire N__28653;
    wire N__28652;
    wire N__28651;
    wire N__28650;
    wire N__28649;
    wire N__28648;
    wire N__28647;
    wire N__28642;
    wire N__28641;
    wire N__28640;
    wire N__28639;
    wire N__28638;
    wire N__28637;
    wire N__28636;
    wire N__28633;
    wire N__28632;
    wire N__28631;
    wire N__28628;
    wire N__28621;
    wire N__28616;
    wire N__28615;
    wire N__28614;
    wire N__28613;
    wire N__28612;
    wire N__28611;
    wire N__28610;
    wire N__28607;
    wire N__28602;
    wire N__28601;
    wire N__28600;
    wire N__28599;
    wire N__28598;
    wire N__28597;
    wire N__28596;
    wire N__28591;
    wire N__28590;
    wire N__28589;
    wire N__28586;
    wire N__28585;
    wire N__28580;
    wire N__28577;
    wire N__28572;
    wire N__28567;
    wire N__28564;
    wire N__28561;
    wire N__28556;
    wire N__28551;
    wire N__28550;
    wire N__28549;
    wire N__28548;
    wire N__28547;
    wire N__28546;
    wire N__28539;
    wire N__28534;
    wire N__28531;
    wire N__28528;
    wire N__28523;
    wire N__28520;
    wire N__28517;
    wire N__28510;
    wire N__28507;
    wire N__28506;
    wire N__28505;
    wire N__28504;
    wire N__28503;
    wire N__28500;
    wire N__28499;
    wire N__28498;
    wire N__28497;
    wire N__28494;
    wire N__28493;
    wire N__28490;
    wire N__28487;
    wire N__28484;
    wire N__28483;
    wire N__28480;
    wire N__28477;
    wire N__28474;
    wire N__28469;
    wire N__28466;
    wire N__28465;
    wire N__28462;
    wire N__28455;
    wire N__28450;
    wire N__28449;
    wire N__28448;
    wire N__28447;
    wire N__28442;
    wire N__28431;
    wire N__28426;
    wire N__28423;
    wire N__28420;
    wire N__28411;
    wire N__28408;
    wire N__28401;
    wire N__28394;
    wire N__28387;
    wire N__28384;
    wire N__28381;
    wire N__28378;
    wire N__28373;
    wire N__28368;
    wire N__28363;
    wire N__28362;
    wire N__28361;
    wire N__28360;
    wire N__28357;
    wire N__28354;
    wire N__28347;
    wire N__28340;
    wire N__28329;
    wire N__28314;
    wire N__28305;
    wire N__28302;
    wire N__28299;
    wire N__28296;
    wire N__28293;
    wire N__28288;
    wire N__28281;
    wire N__28278;
    wire N__28263;
    wire N__28260;
    wire N__28257;
    wire N__28256;
    wire N__28251;
    wire N__28248;
    wire N__28245;
    wire N__28242;
    wire N__28239;
    wire N__28236;
    wire N__28233;
    wire N__28230;
    wire N__28227;
    wire N__28224;
    wire N__28221;
    wire N__28218;
    wire N__28215;
    wire N__28212;
    wire N__28209;
    wire N__28206;
    wire N__28203;
    wire N__28200;
    wire N__28197;
    wire N__28194;
    wire N__28191;
    wire N__28188;
    wire N__28185;
    wire N__28182;
    wire N__28179;
    wire N__28176;
    wire N__28173;
    wire N__28170;
    wire N__28167;
    wire N__28164;
    wire N__28161;
    wire N__28158;
    wire N__28155;
    wire N__28152;
    wire N__28149;
    wire N__28146;
    wire N__28143;
    wire N__28140;
    wire N__28137;
    wire N__28134;
    wire N__28131;
    wire N__28128;
    wire N__28125;
    wire N__28122;
    wire N__28119;
    wire N__28116;
    wire N__28113;
    wire N__28110;
    wire N__28107;
    wire N__28104;
    wire N__28101;
    wire N__28098;
    wire N__28095;
    wire N__28092;
    wire N__28089;
    wire N__28086;
    wire N__28083;
    wire N__28080;
    wire N__28077;
    wire N__28074;
    wire N__28071;
    wire N__28068;
    wire N__28065;
    wire N__28062;
    wire N__28059;
    wire N__28056;
    wire N__28055;
    wire N__28054;
    wire N__28049;
    wire N__28048;
    wire N__28045;
    wire N__28042;
    wire N__28039;
    wire N__28034;
    wire N__28029;
    wire N__28026;
    wire N__28023;
    wire N__28020;
    wire N__28017;
    wire N__28014;
    wire N__28011;
    wire N__28008;
    wire N__28005;
    wire N__28002;
    wire N__28001;
    wire N__28000;
    wire N__27997;
    wire N__27996;
    wire N__27993;
    wire N__27990;
    wire N__27987;
    wire N__27984;
    wire N__27979;
    wire N__27974;
    wire N__27969;
    wire N__27966;
    wire N__27963;
    wire N__27960;
    wire N__27957;
    wire N__27954;
    wire N__27951;
    wire N__27948;
    wire N__27945;
    wire N__27942;
    wire N__27941;
    wire N__27938;
    wire N__27937;
    wire N__27934;
    wire N__27929;
    wire N__27928;
    wire N__27925;
    wire N__27922;
    wire N__27919;
    wire N__27916;
    wire N__27911;
    wire N__27906;
    wire N__27903;
    wire N__27900;
    wire N__27897;
    wire N__27894;
    wire N__27891;
    wire N__27890;
    wire N__27889;
    wire N__27886;
    wire N__27883;
    wire N__27880;
    wire N__27877;
    wire N__27874;
    wire N__27873;
    wire N__27870;
    wire N__27867;
    wire N__27864;
    wire N__27861;
    wire N__27858;
    wire N__27855;
    wire N__27852;
    wire N__27843;
    wire N__27842;
    wire N__27841;
    wire N__27840;
    wire N__27839;
    wire N__27836;
    wire N__27835;
    wire N__27834;
    wire N__27833;
    wire N__27832;
    wire N__27831;
    wire N__27830;
    wire N__27823;
    wire N__27822;
    wire N__27821;
    wire N__27820;
    wire N__27819;
    wire N__27818;
    wire N__27817;
    wire N__27816;
    wire N__27813;
    wire N__27808;
    wire N__27805;
    wire N__27802;
    wire N__27801;
    wire N__27800;
    wire N__27799;
    wire N__27798;
    wire N__27797;
    wire N__27796;
    wire N__27795;
    wire N__27794;
    wire N__27793;
    wire N__27790;
    wire N__27787;
    wire N__27786;
    wire N__27783;
    wire N__27782;
    wire N__27781;
    wire N__27780;
    wire N__27777;
    wire N__27770;
    wire N__27761;
    wire N__27756;
    wire N__27753;
    wire N__27748;
    wire N__27739;
    wire N__27730;
    wire N__27721;
    wire N__27714;
    wire N__27709;
    wire N__27702;
    wire N__27687;
    wire N__27684;
    wire N__27681;
    wire N__27678;
    wire N__27675;
    wire N__27672;
    wire N__27669;
    wire N__27666;
    wire N__27663;
    wire N__27660;
    wire N__27657;
    wire N__27656;
    wire N__27655;
    wire N__27652;
    wire N__27649;
    wire N__27648;
    wire N__27645;
    wire N__27642;
    wire N__27639;
    wire N__27636;
    wire N__27635;
    wire N__27632;
    wire N__27627;
    wire N__27624;
    wire N__27621;
    wire N__27616;
    wire N__27613;
    wire N__27606;
    wire N__27603;
    wire N__27600;
    wire N__27597;
    wire N__27596;
    wire N__27595;
    wire N__27592;
    wire N__27589;
    wire N__27586;
    wire N__27579;
    wire N__27576;
    wire N__27573;
    wire N__27570;
    wire N__27567;
    wire N__27566;
    wire N__27563;
    wire N__27562;
    wire N__27557;
    wire N__27554;
    wire N__27551;
    wire N__27546;
    wire N__27545;
    wire N__27542;
    wire N__27539;
    wire N__27536;
    wire N__27531;
    wire N__27530;
    wire N__27527;
    wire N__27524;
    wire N__27521;
    wire N__27516;
    wire N__27515;
    wire N__27514;
    wire N__27511;
    wire N__27506;
    wire N__27503;
    wire N__27498;
    wire N__27495;
    wire N__27492;
    wire N__27489;
    wire N__27486;
    wire N__27483;
    wire N__27482;
    wire N__27481;
    wire N__27478;
    wire N__27475;
    wire N__27472;
    wire N__27467;
    wire N__27462;
    wire N__27459;
    wire N__27456;
    wire N__27453;
    wire N__27452;
    wire N__27451;
    wire N__27444;
    wire N__27441;
    wire N__27438;
    wire N__27435;
    wire N__27432;
    wire N__27431;
    wire N__27430;
    wire N__27425;
    wire N__27422;
    wire N__27419;
    wire N__27416;
    wire N__27413;
    wire N__27408;
    wire N__27405;
    wire N__27402;
    wire N__27399;
    wire N__27396;
    wire N__27395;
    wire N__27392;
    wire N__27391;
    wire N__27388;
    wire N__27385;
    wire N__27382;
    wire N__27379;
    wire N__27374;
    wire N__27371;
    wire N__27368;
    wire N__27363;
    wire N__27360;
    wire N__27357;
    wire N__27354;
    wire N__27351;
    wire N__27348;
    wire N__27347;
    wire N__27346;
    wire N__27343;
    wire N__27338;
    wire N__27333;
    wire N__27330;
    wire N__27327;
    wire N__27324;
    wire N__27323;
    wire N__27322;
    wire N__27319;
    wire N__27316;
    wire N__27313;
    wire N__27308;
    wire N__27305;
    wire N__27302;
    wire N__27297;
    wire N__27294;
    wire N__27291;
    wire N__27288;
    wire N__27285;
    wire N__27282;
    wire N__27281;
    wire N__27278;
    wire N__27277;
    wire N__27272;
    wire N__27269;
    wire N__27264;
    wire N__27263;
    wire N__27260;
    wire N__27259;
    wire N__27258;
    wire N__27255;
    wire N__27252;
    wire N__27249;
    wire N__27246;
    wire N__27243;
    wire N__27240;
    wire N__27235;
    wire N__27232;
    wire N__27227;
    wire N__27222;
    wire N__27219;
    wire N__27216;
    wire N__27213;
    wire N__27210;
    wire N__27207;
    wire N__27206;
    wire N__27203;
    wire N__27202;
    wire N__27199;
    wire N__27198;
    wire N__27195;
    wire N__27192;
    wire N__27189;
    wire N__27186;
    wire N__27179;
    wire N__27174;
    wire N__27171;
    wire N__27168;
    wire N__27165;
    wire N__27162;
    wire N__27159;
    wire N__27158;
    wire N__27155;
    wire N__27152;
    wire N__27151;
    wire N__27148;
    wire N__27147;
    wire N__27144;
    wire N__27141;
    wire N__27138;
    wire N__27135;
    wire N__27132;
    wire N__27125;
    wire N__27122;
    wire N__27119;
    wire N__27114;
    wire N__27111;
    wire N__27108;
    wire N__27105;
    wire N__27102;
    wire N__27099;
    wire N__27096;
    wire N__27095;
    wire N__27092;
    wire N__27089;
    wire N__27086;
    wire N__27083;
    wire N__27082;
    wire N__27081;
    wire N__27078;
    wire N__27075;
    wire N__27070;
    wire N__27063;
    wire N__27060;
    wire N__27057;
    wire N__27054;
    wire N__27051;
    wire N__27048;
    wire N__27045;
    wire N__27042;
    wire N__27039;
    wire N__27036;
    wire N__27033;
    wire N__27030;
    wire N__27027;
    wire N__27026;
    wire N__27025;
    wire N__27024;
    wire N__27021;
    wire N__27016;
    wire N__27013;
    wire N__27008;
    wire N__27005;
    wire N__27002;
    wire N__26997;
    wire N__26994;
    wire N__26991;
    wire N__26988;
    wire N__26985;
    wire N__26982;
    wire N__26979;
    wire N__26976;
    wire N__26973;
    wire N__26970;
    wire N__26967;
    wire N__26964;
    wire N__26963;
    wire N__26962;
    wire N__26959;
    wire N__26956;
    wire N__26953;
    wire N__26948;
    wire N__26943;
    wire N__26940;
    wire N__26937;
    wire N__26936;
    wire N__26935;
    wire N__26932;
    wire N__26927;
    wire N__26922;
    wire N__26919;
    wire N__26916;
    wire N__26913;
    wire N__26910;
    wire N__26907;
    wire N__26904;
    wire N__26901;
    wire N__26900;
    wire N__26899;
    wire N__26892;
    wire N__26889;
    wire N__26886;
    wire N__26883;
    wire N__26880;
    wire N__26879;
    wire N__26876;
    wire N__26873;
    wire N__26868;
    wire N__26867;
    wire N__26866;
    wire N__26861;
    wire N__26858;
    wire N__26853;
    wire N__26852;
    wire N__26849;
    wire N__26848;
    wire N__26847;
    wire N__26844;
    wire N__26841;
    wire N__26840;
    wire N__26839;
    wire N__26836;
    wire N__26833;
    wire N__26830;
    wire N__26827;
    wire N__26826;
    wire N__26823;
    wire N__26820;
    wire N__26819;
    wire N__26818;
    wire N__26815;
    wire N__26810;
    wire N__26807;
    wire N__26804;
    wire N__26799;
    wire N__26794;
    wire N__26791;
    wire N__26788;
    wire N__26785;
    wire N__26780;
    wire N__26769;
    wire N__26766;
    wire N__26763;
    wire N__26760;
    wire N__26757;
    wire N__26754;
    wire N__26753;
    wire N__26752;
    wire N__26751;
    wire N__26750;
    wire N__26747;
    wire N__26746;
    wire N__26743;
    wire N__26742;
    wire N__26741;
    wire N__26740;
    wire N__26735;
    wire N__26730;
    wire N__26727;
    wire N__26724;
    wire N__26721;
    wire N__26720;
    wire N__26717;
    wire N__26714;
    wire N__26711;
    wire N__26708;
    wire N__26705;
    wire N__26702;
    wire N__26699;
    wire N__26696;
    wire N__26691;
    wire N__26686;
    wire N__26679;
    wire N__26670;
    wire N__26667;
    wire N__26664;
    wire N__26661;
    wire N__26658;
    wire N__26655;
    wire N__26652;
    wire N__26649;
    wire N__26646;
    wire N__26645;
    wire N__26640;
    wire N__26639;
    wire N__26636;
    wire N__26633;
    wire N__26632;
    wire N__26629;
    wire N__26626;
    wire N__26623;
    wire N__26618;
    wire N__26613;
    wire N__26612;
    wire N__26611;
    wire N__26610;
    wire N__26609;
    wire N__26608;
    wire N__26607;
    wire N__26602;
    wire N__26601;
    wire N__26600;
    wire N__26599;
    wire N__26598;
    wire N__26597;
    wire N__26596;
    wire N__26593;
    wire N__26590;
    wire N__26589;
    wire N__26588;
    wire N__26587;
    wire N__26586;
    wire N__26585;
    wire N__26584;
    wire N__26583;
    wire N__26582;
    wire N__26581;
    wire N__26580;
    wire N__26579;
    wire N__26578;
    wire N__26577;
    wire N__26576;
    wire N__26575;
    wire N__26574;
    wire N__26573;
    wire N__26572;
    wire N__26571;
    wire N__26568;
    wire N__26567;
    wire N__26566;
    wire N__26565;
    wire N__26564;
    wire N__26563;
    wire N__26562;
    wire N__26561;
    wire N__26560;
    wire N__26559;
    wire N__26558;
    wire N__26557;
    wire N__26556;
    wire N__26555;
    wire N__26554;
    wire N__26551;
    wire N__26548;
    wire N__26547;
    wire N__26546;
    wire N__26545;
    wire N__26544;
    wire N__26543;
    wire N__26542;
    wire N__26539;
    wire N__26538;
    wire N__26531;
    wire N__26524;
    wire N__26519;
    wire N__26518;
    wire N__26517;
    wire N__26516;
    wire N__26515;
    wire N__26514;
    wire N__26513;
    wire N__26512;
    wire N__26511;
    wire N__26510;
    wire N__26509;
    wire N__26508;
    wire N__26501;
    wire N__26494;
    wire N__26491;
    wire N__26484;
    wire N__26475;
    wire N__26464;
    wire N__26461;
    wire N__26460;
    wire N__26459;
    wire N__26452;
    wire N__26449;
    wire N__26446;
    wire N__26443;
    wire N__26440;
    wire N__26433;
    wire N__26424;
    wire N__26419;
    wire N__26416;
    wire N__26415;
    wire N__26410;
    wire N__26407;
    wire N__26404;
    wire N__26401;
    wire N__26398;
    wire N__26395;
    wire N__26390;
    wire N__26387;
    wire N__26386;
    wire N__26385;
    wire N__26384;
    wire N__26383;
    wire N__26382;
    wire N__26381;
    wire N__26380;
    wire N__26379;
    wire N__26378;
    wire N__26377;
    wire N__26376;
    wire N__26375;
    wire N__26374;
    wire N__26373;
    wire N__26372;
    wire N__26371;
    wire N__26370;
    wire N__26369;
    wire N__26368;
    wire N__26367;
    wire N__26366;
    wire N__26365;
    wire N__26364;
    wire N__26363;
    wire N__26362;
    wire N__26361;
    wire N__26360;
    wire N__26359;
    wire N__26358;
    wire N__26357;
    wire N__26356;
    wire N__26355;
    wire N__26354;
    wire N__26353;
    wire N__26352;
    wire N__26351;
    wire N__26350;
    wire N__26349;
    wire N__26348;
    wire N__26347;
    wire N__26346;
    wire N__26345;
    wire N__26344;
    wire N__26343;
    wire N__26342;
    wire N__26341;
    wire N__26340;
    wire N__26339;
    wire N__26338;
    wire N__26337;
    wire N__26336;
    wire N__26335;
    wire N__26334;
    wire N__26333;
    wire N__26330;
    wire N__26327;
    wire N__26318;
    wire N__26307;
    wire N__26304;
    wire N__26301;
    wire N__26290;
    wire N__26285;
    wire N__26282;
    wire N__26279;
    wire N__26270;
    wire N__26265;
    wire N__26260;
    wire N__26255;
    wire N__26250;
    wire N__26241;
    wire N__26236;
    wire N__26219;
    wire N__26208;
    wire N__26193;
    wire N__26180;
    wire N__26167;
    wire N__26152;
    wire N__26135;
    wire N__26124;
    wire N__26121;
    wire N__26118;
    wire N__26115;
    wire N__26106;
    wire N__26095;
    wire N__26086;
    wire N__26055;
    wire N__26054;
    wire N__26053;
    wire N__26052;
    wire N__26049;
    wire N__26046;
    wire N__26043;
    wire N__26042;
    wire N__26039;
    wire N__26036;
    wire N__26033;
    wire N__26032;
    wire N__26029;
    wire N__26026;
    wire N__26023;
    wire N__26022;
    wire N__26017;
    wire N__26014;
    wire N__26011;
    wire N__26006;
    wire N__26003;
    wire N__26000;
    wire N__25993;
    wire N__25986;
    wire N__25985;
    wire N__25984;
    wire N__25983;
    wire N__25978;
    wire N__25975;
    wire N__25972;
    wire N__25969;
    wire N__25968;
    wire N__25963;
    wire N__25962;
    wire N__25959;
    wire N__25956;
    wire N__25953;
    wire N__25950;
    wire N__25941;
    wire N__25940;
    wire N__25939;
    wire N__25938;
    wire N__25937;
    wire N__25936;
    wire N__25935;
    wire N__25934;
    wire N__25931;
    wire N__25928;
    wire N__25925;
    wire N__25920;
    wire N__25917;
    wire N__25912;
    wire N__25907;
    wire N__25904;
    wire N__25901;
    wire N__25898;
    wire N__25893;
    wire N__25884;
    wire N__25881;
    wire N__25878;
    wire N__25875;
    wire N__25872;
    wire N__25869;
    wire N__25868;
    wire N__25867;
    wire N__25866;
    wire N__25863;
    wire N__25858;
    wire N__25855;
    wire N__25852;
    wire N__25849;
    wire N__25846;
    wire N__25843;
    wire N__25840;
    wire N__25833;
    wire N__25830;
    wire N__25827;
    wire N__25824;
    wire N__25821;
    wire N__25818;
    wire N__25815;
    wire N__25812;
    wire N__25809;
    wire N__25806;
    wire N__25803;
    wire N__25800;
    wire N__25797;
    wire N__25794;
    wire N__25793;
    wire N__25792;
    wire N__25791;
    wire N__25788;
    wire N__25785;
    wire N__25782;
    wire N__25777;
    wire N__25774;
    wire N__25773;
    wire N__25772;
    wire N__25771;
    wire N__25768;
    wire N__25765;
    wire N__25762;
    wire N__25759;
    wire N__25754;
    wire N__25749;
    wire N__25740;
    wire N__25737;
    wire N__25736;
    wire N__25735;
    wire N__25734;
    wire N__25731;
    wire N__25730;
    wire N__25729;
    wire N__25726;
    wire N__25721;
    wire N__25718;
    wire N__25713;
    wire N__25710;
    wire N__25701;
    wire N__25698;
    wire N__25695;
    wire N__25692;
    wire N__25689;
    wire N__25686;
    wire N__25683;
    wire N__25680;
    wire N__25677;
    wire N__25676;
    wire N__25673;
    wire N__25672;
    wire N__25669;
    wire N__25666;
    wire N__25663;
    wire N__25660;
    wire N__25655;
    wire N__25650;
    wire N__25647;
    wire N__25644;
    wire N__25641;
    wire N__25638;
    wire N__25635;
    wire N__25632;
    wire N__25629;
    wire N__25626;
    wire N__25625;
    wire N__25624;
    wire N__25623;
    wire N__25620;
    wire N__25613;
    wire N__25608;
    wire N__25605;
    wire N__25602;
    wire N__25599;
    wire N__25598;
    wire N__25595;
    wire N__25592;
    wire N__25591;
    wire N__25588;
    wire N__25585;
    wire N__25584;
    wire N__25581;
    wire N__25578;
    wire N__25575;
    wire N__25570;
    wire N__25563;
    wire N__25562;
    wire N__25561;
    wire N__25560;
    wire N__25553;
    wire N__25552;
    wire N__25551;
    wire N__25550;
    wire N__25547;
    wire N__25546;
    wire N__25545;
    wire N__25544;
    wire N__25541;
    wire N__25534;
    wire N__25531;
    wire N__25524;
    wire N__25521;
    wire N__25512;
    wire N__25509;
    wire N__25508;
    wire N__25507;
    wire N__25504;
    wire N__25503;
    wire N__25502;
    wire N__25499;
    wire N__25496;
    wire N__25489;
    wire N__25488;
    wire N__25487;
    wire N__25486;
    wire N__25485;
    wire N__25484;
    wire N__25479;
    wire N__25476;
    wire N__25469;
    wire N__25464;
    wire N__25461;
    wire N__25458;
    wire N__25449;
    wire N__25446;
    wire N__25443;
    wire N__25440;
    wire N__25437;
    wire N__25434;
    wire N__25433;
    wire N__25432;
    wire N__25431;
    wire N__25426;
    wire N__25423;
    wire N__25420;
    wire N__25417;
    wire N__25414;
    wire N__25411;
    wire N__25404;
    wire N__25401;
    wire N__25398;
    wire N__25395;
    wire N__25392;
    wire N__25389;
    wire N__25386;
    wire N__25383;
    wire N__25380;
    wire N__25377;
    wire N__25374;
    wire N__25371;
    wire N__25368;
    wire N__25365;
    wire N__25362;
    wire N__25359;
    wire N__25356;
    wire N__25353;
    wire N__25350;
    wire N__25347;
    wire N__25344;
    wire N__25343;
    wire N__25342;
    wire N__25337;
    wire N__25334;
    wire N__25331;
    wire N__25328;
    wire N__25327;
    wire N__25322;
    wire N__25319;
    wire N__25316;
    wire N__25311;
    wire N__25308;
    wire N__25305;
    wire N__25302;
    wire N__25299;
    wire N__25298;
    wire N__25295;
    wire N__25292;
    wire N__25289;
    wire N__25288;
    wire N__25285;
    wire N__25282;
    wire N__25281;
    wire N__25278;
    wire N__25275;
    wire N__25272;
    wire N__25269;
    wire N__25266;
    wire N__25257;
    wire N__25254;
    wire N__25251;
    wire N__25248;
    wire N__25245;
    wire N__25242;
    wire N__25239;
    wire N__25236;
    wire N__25233;
    wire N__25230;
    wire N__25227;
    wire N__25224;
    wire N__25221;
    wire N__25220;
    wire N__25219;
    wire N__25218;
    wire N__25215;
    wire N__25212;
    wire N__25207;
    wire N__25204;
    wire N__25201;
    wire N__25198;
    wire N__25195;
    wire N__25192;
    wire N__25189;
    wire N__25182;
    wire N__25179;
    wire N__25176;
    wire N__25173;
    wire N__25170;
    wire N__25169;
    wire N__25166;
    wire N__25163;
    wire N__25160;
    wire N__25159;
    wire N__25158;
    wire N__25155;
    wire N__25152;
    wire N__25147;
    wire N__25140;
    wire N__25137;
    wire N__25134;
    wire N__25131;
    wire N__25128;
    wire N__25125;
    wire N__25124;
    wire N__25121;
    wire N__25120;
    wire N__25119;
    wire N__25116;
    wire N__25113;
    wire N__25110;
    wire N__25107;
    wire N__25104;
    wire N__25101;
    wire N__25096;
    wire N__25093;
    wire N__25090;
    wire N__25087;
    wire N__25082;
    wire N__25079;
    wire N__25074;
    wire N__25071;
    wire N__25068;
    wire N__25065;
    wire N__25062;
    wire N__25059;
    wire N__25056;
    wire N__25055;
    wire N__25054;
    wire N__25053;
    wire N__25050;
    wire N__25045;
    wire N__25042;
    wire N__25039;
    wire N__25036;
    wire N__25033;
    wire N__25030;
    wire N__25027;
    wire N__25020;
    wire N__25017;
    wire N__25014;
    wire N__25011;
    wire N__25008;
    wire N__25007;
    wire N__25004;
    wire N__25001;
    wire N__24998;
    wire N__24995;
    wire N__24994;
    wire N__24993;
    wire N__24990;
    wire N__24987;
    wire N__24982;
    wire N__24979;
    wire N__24974;
    wire N__24969;
    wire N__24966;
    wire N__24963;
    wire N__24960;
    wire N__24957;
    wire N__24954;
    wire N__24951;
    wire N__24948;
    wire N__24945;
    wire N__24942;
    wire N__24941;
    wire N__24938;
    wire N__24937;
    wire N__24936;
    wire N__24933;
    wire N__24930;
    wire N__24927;
    wire N__24924;
    wire N__24921;
    wire N__24916;
    wire N__24915;
    wire N__24912;
    wire N__24909;
    wire N__24906;
    wire N__24905;
    wire N__24904;
    wire N__24901;
    wire N__24896;
    wire N__24893;
    wire N__24888;
    wire N__24879;
    wire N__24876;
    wire N__24873;
    wire N__24870;
    wire N__24869;
    wire N__24866;
    wire N__24863;
    wire N__24860;
    wire N__24857;
    wire N__24852;
    wire N__24851;
    wire N__24850;
    wire N__24847;
    wire N__24846;
    wire N__24845;
    wire N__24842;
    wire N__24839;
    wire N__24836;
    wire N__24833;
    wire N__24832;
    wire N__24829;
    wire N__24826;
    wire N__24823;
    wire N__24818;
    wire N__24815;
    wire N__24812;
    wire N__24805;
    wire N__24798;
    wire N__24795;
    wire N__24792;
    wire N__24789;
    wire N__24786;
    wire N__24783;
    wire N__24782;
    wire N__24779;
    wire N__24778;
    wire N__24775;
    wire N__24774;
    wire N__24771;
    wire N__24768;
    wire N__24765;
    wire N__24762;
    wire N__24759;
    wire N__24750;
    wire N__24749;
    wire N__24748;
    wire N__24745;
    wire N__24744;
    wire N__24743;
    wire N__24740;
    wire N__24737;
    wire N__24734;
    wire N__24731;
    wire N__24728;
    wire N__24725;
    wire N__24722;
    wire N__24719;
    wire N__24716;
    wire N__24705;
    wire N__24702;
    wire N__24699;
    wire N__24698;
    wire N__24695;
    wire N__24692;
    wire N__24689;
    wire N__24686;
    wire N__24681;
    wire N__24678;
    wire N__24675;
    wire N__24674;
    wire N__24673;
    wire N__24672;
    wire N__24669;
    wire N__24662;
    wire N__24657;
    wire N__24654;
    wire N__24653;
    wire N__24652;
    wire N__24651;
    wire N__24648;
    wire N__24643;
    wire N__24640;
    wire N__24637;
    wire N__24636;
    wire N__24633;
    wire N__24630;
    wire N__24627;
    wire N__24624;
    wire N__24621;
    wire N__24616;
    wire N__24609;
    wire N__24606;
    wire N__24603;
    wire N__24600;
    wire N__24597;
    wire N__24596;
    wire N__24593;
    wire N__24590;
    wire N__24587;
    wire N__24584;
    wire N__24583;
    wire N__24582;
    wire N__24579;
    wire N__24576;
    wire N__24573;
    wire N__24570;
    wire N__24567;
    wire N__24562;
    wire N__24555;
    wire N__24552;
    wire N__24551;
    wire N__24548;
    wire N__24545;
    wire N__24542;
    wire N__24539;
    wire N__24536;
    wire N__24533;
    wire N__24528;
    wire N__24527;
    wire N__24526;
    wire N__24525;
    wire N__24522;
    wire N__24519;
    wire N__24516;
    wire N__24513;
    wire N__24510;
    wire N__24507;
    wire N__24498;
    wire N__24495;
    wire N__24492;
    wire N__24489;
    wire N__24486;
    wire N__24483;
    wire N__24482;
    wire N__24481;
    wire N__24478;
    wire N__24475;
    wire N__24472;
    wire N__24471;
    wire N__24468;
    wire N__24465;
    wire N__24464;
    wire N__24461;
    wire N__24458;
    wire N__24453;
    wire N__24450;
    wire N__24447;
    wire N__24442;
    wire N__24435;
    wire N__24434;
    wire N__24433;
    wire N__24430;
    wire N__24427;
    wire N__24426;
    wire N__24423;
    wire N__24422;
    wire N__24419;
    wire N__24416;
    wire N__24411;
    wire N__24408;
    wire N__24401;
    wire N__24396;
    wire N__24393;
    wire N__24390;
    wire N__24387;
    wire N__24384;
    wire N__24381;
    wire N__24380;
    wire N__24377;
    wire N__24374;
    wire N__24371;
    wire N__24368;
    wire N__24367;
    wire N__24362;
    wire N__24359;
    wire N__24358;
    wire N__24357;
    wire N__24354;
    wire N__24351;
    wire N__24350;
    wire N__24347;
    wire N__24344;
    wire N__24339;
    wire N__24336;
    wire N__24327;
    wire N__24324;
    wire N__24323;
    wire N__24320;
    wire N__24317;
    wire N__24316;
    wire N__24315;
    wire N__24312;
    wire N__24309;
    wire N__24308;
    wire N__24305;
    wire N__24302;
    wire N__24299;
    wire N__24296;
    wire N__24293;
    wire N__24282;
    wire N__24279;
    wire N__24276;
    wire N__24273;
    wire N__24272;
    wire N__24271;
    wire N__24270;
    wire N__24269;
    wire N__24266;
    wire N__24265;
    wire N__24264;
    wire N__24261;
    wire N__24258;
    wire N__24255;
    wire N__24254;
    wire N__24251;
    wire N__24248;
    wire N__24245;
    wire N__24242;
    wire N__24239;
    wire N__24236;
    wire N__24233;
    wire N__24230;
    wire N__24227;
    wire N__24224;
    wire N__24221;
    wire N__24218;
    wire N__24209;
    wire N__24206;
    wire N__24201;
    wire N__24198;
    wire N__24195;
    wire N__24192;
    wire N__24189;
    wire N__24184;
    wire N__24177;
    wire N__24176;
    wire N__24173;
    wire N__24170;
    wire N__24167;
    wire N__24164;
    wire N__24163;
    wire N__24160;
    wire N__24157;
    wire N__24156;
    wire N__24153;
    wire N__24148;
    wire N__24145;
    wire N__24138;
    wire N__24137;
    wire N__24134;
    wire N__24133;
    wire N__24130;
    wire N__24129;
    wire N__24126;
    wire N__24123;
    wire N__24120;
    wire N__24117;
    wire N__24114;
    wire N__24105;
    wire N__24102;
    wire N__24099;
    wire N__24098;
    wire N__24095;
    wire N__24092;
    wire N__24089;
    wire N__24086;
    wire N__24081;
    wire N__24080;
    wire N__24079;
    wire N__24074;
    wire N__24073;
    wire N__24070;
    wire N__24067;
    wire N__24064;
    wire N__24063;
    wire N__24060;
    wire N__24057;
    wire N__24054;
    wire N__24051;
    wire N__24048;
    wire N__24043;
    wire N__24036;
    wire N__24033;
    wire N__24032;
    wire N__24031;
    wire N__24028;
    wire N__24025;
    wire N__24024;
    wire N__24021;
    wire N__24018;
    wire N__24015;
    wire N__24012;
    wire N__24003;
    wire N__24000;
    wire N__23999;
    wire N__23996;
    wire N__23993;
    wire N__23992;
    wire N__23989;
    wire N__23986;
    wire N__23985;
    wire N__23982;
    wire N__23979;
    wire N__23976;
    wire N__23973;
    wire N__23964;
    wire N__23961;
    wire N__23960;
    wire N__23959;
    wire N__23958;
    wire N__23955;
    wire N__23952;
    wire N__23949;
    wire N__23946;
    wire N__23943;
    wire N__23940;
    wire N__23931;
    wire N__23928;
    wire N__23925;
    wire N__23922;
    wire N__23919;
    wire N__23918;
    wire N__23917;
    wire N__23916;
    wire N__23911;
    wire N__23910;
    wire N__23907;
    wire N__23904;
    wire N__23903;
    wire N__23902;
    wire N__23899;
    wire N__23896;
    wire N__23893;
    wire N__23890;
    wire N__23887;
    wire N__23884;
    wire N__23881;
    wire N__23878;
    wire N__23873;
    wire N__23870;
    wire N__23859;
    wire N__23856;
    wire N__23853;
    wire N__23852;
    wire N__23851;
    wire N__23848;
    wire N__23845;
    wire N__23844;
    wire N__23841;
    wire N__23836;
    wire N__23833;
    wire N__23830;
    wire N__23827;
    wire N__23820;
    wire N__23819;
    wire N__23816;
    wire N__23815;
    wire N__23814;
    wire N__23811;
    wire N__23808;
    wire N__23805;
    wire N__23802;
    wire N__23799;
    wire N__23794;
    wire N__23787;
    wire N__23784;
    wire N__23781;
    wire N__23778;
    wire N__23775;
    wire N__23772;
    wire N__23771;
    wire N__23768;
    wire N__23763;
    wire N__23762;
    wire N__23759;
    wire N__23756;
    wire N__23751;
    wire N__23748;
    wire N__23745;
    wire N__23744;
    wire N__23741;
    wire N__23738;
    wire N__23735;
    wire N__23732;
    wire N__23729;
    wire N__23726;
    wire N__23725;
    wire N__23724;
    wire N__23723;
    wire N__23718;
    wire N__23715;
    wire N__23712;
    wire N__23709;
    wire N__23706;
    wire N__23703;
    wire N__23694;
    wire N__23691;
    wire N__23688;
    wire N__23687;
    wire N__23684;
    wire N__23681;
    wire N__23676;
    wire N__23673;
    wire N__23670;
    wire N__23667;
    wire N__23666;
    wire N__23663;
    wire N__23660;
    wire N__23655;
    wire N__23654;
    wire N__23653;
    wire N__23652;
    wire N__23649;
    wire N__23646;
    wire N__23643;
    wire N__23640;
    wire N__23637;
    wire N__23634;
    wire N__23631;
    wire N__23622;
    wire N__23621;
    wire N__23618;
    wire N__23615;
    wire N__23614;
    wire N__23613;
    wire N__23612;
    wire N__23609;
    wire N__23606;
    wire N__23603;
    wire N__23602;
    wire N__23599;
    wire N__23596;
    wire N__23589;
    wire N__23586;
    wire N__23577;
    wire N__23574;
    wire N__23571;
    wire N__23568;
    wire N__23565;
    wire N__23564;
    wire N__23563;
    wire N__23558;
    wire N__23555;
    wire N__23554;
    wire N__23551;
    wire N__23548;
    wire N__23547;
    wire N__23546;
    wire N__23543;
    wire N__23540;
    wire N__23537;
    wire N__23532;
    wire N__23523;
    wire N__23522;
    wire N__23519;
    wire N__23516;
    wire N__23513;
    wire N__23510;
    wire N__23505;
    wire N__23504;
    wire N__23503;
    wire N__23500;
    wire N__23495;
    wire N__23490;
    wire N__23487;
    wire N__23484;
    wire N__23483;
    wire N__23482;
    wire N__23479;
    wire N__23476;
    wire N__23475;
    wire N__23472;
    wire N__23469;
    wire N__23462;
    wire N__23459;
    wire N__23454;
    wire N__23453;
    wire N__23450;
    wire N__23449;
    wire N__23448;
    wire N__23447;
    wire N__23444;
    wire N__23441;
    wire N__23438;
    wire N__23435;
    wire N__23432;
    wire N__23429;
    wire N__23426;
    wire N__23423;
    wire N__23412;
    wire N__23409;
    wire N__23406;
    wire N__23403;
    wire N__23400;
    wire N__23397;
    wire N__23396;
    wire N__23393;
    wire N__23390;
    wire N__23389;
    wire N__23388;
    wire N__23385;
    wire N__23382;
    wire N__23381;
    wire N__23378;
    wire N__23375;
    wire N__23370;
    wire N__23367;
    wire N__23364;
    wire N__23361;
    wire N__23358;
    wire N__23349;
    wire N__23346;
    wire N__23343;
    wire N__23340;
    wire N__23337;
    wire N__23334;
    wire N__23331;
    wire N__23328;
    wire N__23325;
    wire N__23322;
    wire N__23319;
    wire N__23316;
    wire N__23313;
    wire N__23310;
    wire N__23307;
    wire N__23304;
    wire N__23303;
    wire N__23300;
    wire N__23297;
    wire N__23296;
    wire N__23295;
    wire N__23292;
    wire N__23289;
    wire N__23286;
    wire N__23283;
    wire N__23280;
    wire N__23275;
    wire N__23268;
    wire N__23265;
    wire N__23262;
    wire N__23261;
    wire N__23260;
    wire N__23259;
    wire N__23256;
    wire N__23255;
    wire N__23250;
    wire N__23247;
    wire N__23244;
    wire N__23241;
    wire N__23240;
    wire N__23239;
    wire N__23234;
    wire N__23229;
    wire N__23226;
    wire N__23223;
    wire N__23218;
    wire N__23211;
    wire N__23208;
    wire N__23207;
    wire N__23202;
    wire N__23199;
    wire N__23196;
    wire N__23193;
    wire N__23190;
    wire N__23187;
    wire N__23186;
    wire N__23185;
    wire N__23184;
    wire N__23181;
    wire N__23180;
    wire N__23177;
    wire N__23174;
    wire N__23171;
    wire N__23168;
    wire N__23165;
    wire N__23160;
    wire N__23151;
    wire N__23150;
    wire N__23147;
    wire N__23144;
    wire N__23141;
    wire N__23138;
    wire N__23137;
    wire N__23136;
    wire N__23131;
    wire N__23128;
    wire N__23125;
    wire N__23124;
    wire N__23123;
    wire N__23120;
    wire N__23115;
    wire N__23110;
    wire N__23103;
    wire N__23100;
    wire N__23097;
    wire N__23094;
    wire N__23091;
    wire N__23088;
    wire N__23085;
    wire N__23084;
    wire N__23081;
    wire N__23078;
    wire N__23073;
    wire N__23070;
    wire N__23067;
    wire N__23064;
    wire N__23061;
    wire N__23058;
    wire N__23055;
    wire N__23052;
    wire N__23049;
    wire N__23046;
    wire N__23045;
    wire N__23042;
    wire N__23039;
    wire N__23036;
    wire N__23031;
    wire N__23028;
    wire N__23025;
    wire N__23024;
    wire N__23023;
    wire N__23020;
    wire N__23019;
    wire N__23016;
    wire N__23013;
    wire N__23012;
    wire N__23009;
    wire N__23006;
    wire N__23003;
    wire N__23000;
    wire N__22997;
    wire N__22994;
    wire N__22991;
    wire N__22988;
    wire N__22985;
    wire N__22974;
    wire N__22973;
    wire N__22972;
    wire N__22969;
    wire N__22966;
    wire N__22963;
    wire N__22962;
    wire N__22959;
    wire N__22954;
    wire N__22951;
    wire N__22946;
    wire N__22941;
    wire N__22938;
    wire N__22937;
    wire N__22934;
    wire N__22931;
    wire N__22928;
    wire N__22927;
    wire N__22922;
    wire N__22921;
    wire N__22918;
    wire N__22915;
    wire N__22912;
    wire N__22905;
    wire N__22902;
    wire N__22899;
    wire N__22896;
    wire N__22893;
    wire N__22890;
    wire N__22887;
    wire N__22884;
    wire N__22881;
    wire N__22880;
    wire N__22875;
    wire N__22872;
    wire N__22869;
    wire N__22868;
    wire N__22867;
    wire N__22864;
    wire N__22859;
    wire N__22854;
    wire N__22853;
    wire N__22852;
    wire N__22849;
    wire N__22844;
    wire N__22839;
    wire N__22836;
    wire N__22833;
    wire N__22830;
    wire N__22827;
    wire N__22824;
    wire N__22821;
    wire N__22818;
    wire N__22815;
    wire N__22812;
    wire N__22809;
    wire N__22806;
    wire N__22803;
    wire N__22800;
    wire N__22797;
    wire N__22794;
    wire N__22791;
    wire N__22788;
    wire N__22785;
    wire N__22782;
    wire N__22779;
    wire N__22776;
    wire N__22773;
    wire N__22770;
    wire N__22767;
    wire N__22764;
    wire N__22761;
    wire N__22758;
    wire N__22755;
    wire N__22752;
    wire N__22749;
    wire N__22746;
    wire N__22743;
    wire N__22740;
    wire N__22737;
    wire N__22734;
    wire N__22731;
    wire N__22728;
    wire N__22725;
    wire N__22722;
    wire N__22719;
    wire N__22716;
    wire N__22713;
    wire N__22710;
    wire N__22707;
    wire N__22704;
    wire N__22701;
    wire N__22698;
    wire N__22695;
    wire N__22694;
    wire N__22693;
    wire N__22690;
    wire N__22687;
    wire N__22684;
    wire N__22683;
    wire N__22680;
    wire N__22677;
    wire N__22672;
    wire N__22669;
    wire N__22666;
    wire N__22659;
    wire N__22656;
    wire N__22653;
    wire N__22650;
    wire N__22647;
    wire N__22644;
    wire N__22641;
    wire N__22638;
    wire N__22635;
    wire N__22632;
    wire N__22631;
    wire N__22630;
    wire N__22627;
    wire N__22626;
    wire N__22621;
    wire N__22618;
    wire N__22615;
    wire N__22612;
    wire N__22609;
    wire N__22606;
    wire N__22599;
    wire N__22596;
    wire N__22593;
    wire N__22590;
    wire N__22587;
    wire N__22584;
    wire N__22581;
    wire N__22578;
    wire N__22575;
    wire N__22574;
    wire N__22571;
    wire N__22568;
    wire N__22565;
    wire N__22560;
    wire N__22559;
    wire N__22556;
    wire N__22553;
    wire N__22550;
    wire N__22545;
    wire N__22542;
    wire N__22541;
    wire N__22538;
    wire N__22535;
    wire N__22532;
    wire N__22527;
    wire N__22524;
    wire N__22521;
    wire N__22518;
    wire N__22515;
    wire N__22512;
    wire N__22509;
    wire N__22506;
    wire N__22503;
    wire N__22500;
    wire N__22497;
    wire N__22494;
    wire N__22491;
    wire N__22488;
    wire N__22485;
    wire N__22482;
    wire N__22479;
    wire N__22476;
    wire N__22473;
    wire N__22470;
    wire N__22467;
    wire N__22464;
    wire N__22461;
    wire N__22458;
    wire N__22455;
    wire N__22452;
    wire N__22449;
    wire N__22446;
    wire N__22443;
    wire N__22440;
    wire N__22437;
    wire N__22434;
    wire N__22431;
    wire N__22428;
    wire N__22425;
    wire N__22422;
    wire N__22419;
    wire N__22416;
    wire N__22413;
    wire N__22410;
    wire N__22407;
    wire N__22404;
    wire N__22401;
    wire N__22398;
    wire N__22395;
    wire N__22392;
    wire N__22389;
    wire N__22386;
    wire N__22383;
    wire N__22380;
    wire N__22377;
    wire N__22374;
    wire N__22373;
    wire N__22370;
    wire N__22367;
    wire N__22362;
    wire N__22359;
    wire N__22356;
    wire N__22353;
    wire N__22350;
    wire N__22347;
    wire N__22344;
    wire N__22341;
    wire N__22338;
    wire N__22335;
    wire N__22332;
    wire N__22329;
    wire N__22326;
    wire N__22323;
    wire N__22322;
    wire N__22319;
    wire N__22316;
    wire N__22313;
    wire N__22308;
    wire N__22305;
    wire N__22304;
    wire N__22301;
    wire N__22298;
    wire N__22295;
    wire N__22290;
    wire N__22287;
    wire N__22284;
    wire N__22283;
    wire N__22282;
    wire N__22277;
    wire N__22274;
    wire N__22271;
    wire N__22266;
    wire N__22263;
    wire N__22262;
    wire N__22259;
    wire N__22256;
    wire N__22251;
    wire N__22248;
    wire N__22247;
    wire N__22244;
    wire N__22241;
    wire N__22236;
    wire N__22233;
    wire N__22230;
    wire N__22229;
    wire N__22226;
    wire N__22223;
    wire N__22220;
    wire N__22215;
    wire N__22214;
    wire N__22211;
    wire N__22208;
    wire N__22205;
    wire N__22202;
    wire N__22199;
    wire N__22194;
    wire N__22193;
    wire N__22192;
    wire N__22189;
    wire N__22186;
    wire N__22183;
    wire N__22182;
    wire N__22177;
    wire N__22174;
    wire N__22171;
    wire N__22166;
    wire N__22163;
    wire N__22160;
    wire N__22157;
    wire N__22154;
    wire N__22151;
    wire N__22146;
    wire N__22145;
    wire N__22142;
    wire N__22139;
    wire N__22136;
    wire N__22131;
    wire N__22128;
    wire N__22125;
    wire N__22122;
    wire N__22121;
    wire N__22118;
    wire N__22115;
    wire N__22114;
    wire N__22109;
    wire N__22106;
    wire N__22103;
    wire N__22100;
    wire N__22095;
    wire N__22094;
    wire N__22093;
    wire N__22090;
    wire N__22087;
    wire N__22084;
    wire N__22081;
    wire N__22074;
    wire N__22071;
    wire N__22068;
    wire N__22067;
    wire N__22062;
    wire N__22059;
    wire N__22058;
    wire N__22055;
    wire N__22052;
    wire N__22047;
    wire N__22044;
    wire N__22043;
    wire N__22042;
    wire N__22037;
    wire N__22034;
    wire N__22031;
    wire N__22026;
    wire N__22023;
    wire N__22022;
    wire N__22019;
    wire N__22016;
    wire N__22011;
    wire N__22008;
    wire N__22005;
    wire N__22002;
    wire N__22001;
    wire N__21998;
    wire N__21995;
    wire N__21992;
    wire N__21987;
    wire N__21984;
    wire N__21981;
    wire N__21978;
    wire N__21977;
    wire N__21974;
    wire N__21971;
    wire N__21968;
    wire N__21963;
    wire N__21962;
    wire N__21959;
    wire N__21958;
    wire N__21957;
    wire N__21956;
    wire N__21955;
    wire N__21952;
    wire N__21949;
    wire N__21946;
    wire N__21943;
    wire N__21940;
    wire N__21937;
    wire N__21934;
    wire N__21931;
    wire N__21928;
    wire N__21925;
    wire N__21922;
    wire N__21919;
    wire N__21914;
    wire N__21911;
    wire N__21906;
    wire N__21897;
    wire N__21896;
    wire N__21895;
    wire N__21894;
    wire N__21893;
    wire N__21890;
    wire N__21887;
    wire N__21882;
    wire N__21879;
    wire N__21870;
    wire N__21869;
    wire N__21868;
    wire N__21867;
    wire N__21866;
    wire N__21861;
    wire N__21860;
    wire N__21857;
    wire N__21854;
    wire N__21851;
    wire N__21848;
    wire N__21845;
    wire N__21842;
    wire N__21839;
    wire N__21828;
    wire N__21825;
    wire N__21824;
    wire N__21821;
    wire N__21820;
    wire N__21817;
    wire N__21814;
    wire N__21811;
    wire N__21808;
    wire N__21805;
    wire N__21800;
    wire N__21795;
    wire N__21794;
    wire N__21791;
    wire N__21788;
    wire N__21787;
    wire N__21784;
    wire N__21783;
    wire N__21780;
    wire N__21777;
    wire N__21774;
    wire N__21771;
    wire N__21768;
    wire N__21765;
    wire N__21762;
    wire N__21753;
    wire N__21752;
    wire N__21749;
    wire N__21746;
    wire N__21745;
    wire N__21742;
    wire N__21741;
    wire N__21740;
    wire N__21737;
    wire N__21734;
    wire N__21731;
    wire N__21726;
    wire N__21717;
    wire N__21714;
    wire N__21713;
    wire N__21710;
    wire N__21707;
    wire N__21704;
    wire N__21699;
    wire N__21696;
    wire N__21693;
    wire N__21690;
    wire N__21687;
    wire N__21684;
    wire N__21681;
    wire N__21680;
    wire N__21677;
    wire N__21674;
    wire N__21671;
    wire N__21666;
    wire N__21665;
    wire N__21664;
    wire N__21661;
    wire N__21660;
    wire N__21657;
    wire N__21654;
    wire N__21651;
    wire N__21648;
    wire N__21645;
    wire N__21642;
    wire N__21639;
    wire N__21630;
    wire N__21627;
    wire N__21624;
    wire N__21621;
    wire N__21618;
    wire N__21615;
    wire N__21612;
    wire N__21609;
    wire N__21606;
    wire N__21603;
    wire N__21600;
    wire N__21597;
    wire N__21594;
    wire N__21591;
    wire N__21588;
    wire N__21585;
    wire N__21582;
    wire N__21579;
    wire N__21576;
    wire N__21573;
    wire N__21572;
    wire N__21571;
    wire N__21568;
    wire N__21565;
    wire N__21564;
    wire N__21561;
    wire N__21558;
    wire N__21555;
    wire N__21552;
    wire N__21547;
    wire N__21544;
    wire N__21537;
    wire N__21534;
    wire N__21531;
    wire N__21528;
    wire N__21525;
    wire N__21524;
    wire N__21523;
    wire N__21522;
    wire N__21519;
    wire N__21516;
    wire N__21513;
    wire N__21510;
    wire N__21509;
    wire N__21506;
    wire N__21503;
    wire N__21500;
    wire N__21497;
    wire N__21494;
    wire N__21491;
    wire N__21486;
    wire N__21483;
    wire N__21474;
    wire N__21471;
    wire N__21468;
    wire N__21467;
    wire N__21464;
    wire N__21461;
    wire N__21458;
    wire N__21457;
    wire N__21456;
    wire N__21453;
    wire N__21450;
    wire N__21447;
    wire N__21444;
    wire N__21441;
    wire N__21436;
    wire N__21429;
    wire N__21426;
    wire N__21423;
    wire N__21420;
    wire N__21417;
    wire N__21416;
    wire N__21413;
    wire N__21410;
    wire N__21405;
    wire N__21402;
    wire N__21399;
    wire N__21396;
    wire N__21393;
    wire N__21390;
    wire N__21387;
    wire N__21384;
    wire N__21381;
    wire N__21378;
    wire N__21375;
    wire N__21372;
    wire N__21369;
    wire N__21368;
    wire N__21365;
    wire N__21364;
    wire N__21361;
    wire N__21360;
    wire N__21359;
    wire N__21354;
    wire N__21353;
    wire N__21350;
    wire N__21347;
    wire N__21344;
    wire N__21341;
    wire N__21338;
    wire N__21335;
    wire N__21324;
    wire N__21321;
    wire N__21318;
    wire N__21315;
    wire N__21312;
    wire N__21311;
    wire N__21308;
    wire N__21305;
    wire N__21304;
    wire N__21301;
    wire N__21300;
    wire N__21297;
    wire N__21294;
    wire N__21293;
    wire N__21290;
    wire N__21287;
    wire N__21284;
    wire N__21279;
    wire N__21274;
    wire N__21267;
    wire N__21264;
    wire N__21261;
    wire N__21258;
    wire N__21255;
    wire N__21252;
    wire N__21249;
    wire N__21246;
    wire N__21243;
    wire N__21240;
    wire N__21237;
    wire N__21234;
    wire N__21231;
    wire N__21228;
    wire N__21225;
    wire N__21222;
    wire N__21219;
    wire N__21216;
    wire N__21213;
    wire N__21212;
    wire N__21211;
    wire N__21210;
    wire N__21207;
    wire N__21204;
    wire N__21203;
    wire N__21200;
    wire N__21199;
    wire N__21196;
    wire N__21195;
    wire N__21194;
    wire N__21191;
    wire N__21188;
    wire N__21185;
    wire N__21182;
    wire N__21179;
    wire N__21176;
    wire N__21173;
    wire N__21170;
    wire N__21167;
    wire N__21162;
    wire N__21153;
    wire N__21150;
    wire N__21145;
    wire N__21142;
    wire N__21135;
    wire N__21132;
    wire N__21131;
    wire N__21128;
    wire N__21125;
    wire N__21120;
    wire N__21119;
    wire N__21116;
    wire N__21113;
    wire N__21108;
    wire N__21105;
    wire N__21102;
    wire N__21099;
    wire N__21096;
    wire N__21093;
    wire N__21090;
    wire N__21087;
    wire N__21084;
    wire N__21081;
    wire N__21078;
    wire N__21075;
    wire N__21072;
    wire N__21069;
    wire N__21066;
    wire N__21063;
    wire N__21060;
    wire N__21057;
    wire N__21054;
    wire N__21051;
    wire N__21048;
    wire N__21045;
    wire N__21042;
    wire N__21039;
    wire N__21036;
    wire N__21033;
    wire N__21030;
    wire N__21027;
    wire N__21024;
    wire N__21021;
    wire N__21018;
    wire N__21015;
    wire N__21012;
    wire N__21009;
    wire N__21006;
    wire N__21003;
    wire N__21002;
    wire N__20999;
    wire N__20996;
    wire N__20991;
    wire N__20990;
    wire N__20987;
    wire N__20984;
    wire N__20979;
    wire N__20976;
    wire N__20973;
    wire N__20970;
    wire N__20967;
    wire N__20964;
    wire N__20961;
    wire N__20958;
    wire N__20955;
    wire N__20952;
    wire N__20949;
    wire N__20948;
    wire N__20947;
    wire N__20946;
    wire N__20943;
    wire N__20936;
    wire N__20933;
    wire N__20930;
    wire N__20927;
    wire N__20924;
    wire N__20919;
    wire N__20916;
    wire N__20913;
    wire N__20910;
    wire N__20907;
    wire N__20904;
    wire N__20901;
    wire N__20898;
    wire N__20895;
    wire N__20892;
    wire N__20889;
    wire N__20886;
    wire N__20883;
    wire N__20880;
    wire N__20879;
    wire N__20878;
    wire N__20877;
    wire N__20874;
    wire N__20867;
    wire N__20862;
    wire N__20859;
    wire N__20856;
    wire N__20853;
    wire N__20850;
    wire N__20847;
    wire N__20844;
    wire N__20841;
    wire N__20838;
    wire N__20835;
    wire N__20832;
    wire N__20829;
    wire N__20826;
    wire N__20823;
    wire N__20820;
    wire N__20817;
    wire N__20814;
    wire N__20811;
    wire N__20808;
    wire N__20805;
    wire N__20802;
    wire N__20799;
    wire N__20798;
    wire N__20797;
    wire N__20796;
    wire N__20793;
    wire N__20786;
    wire N__20781;
    wire N__20778;
    wire N__20775;
    wire N__20772;
    wire N__20769;
    wire N__20766;
    wire N__20763;
    wire N__20760;
    wire N__20757;
    wire N__20754;
    wire N__20751;
    wire N__20748;
    wire N__20745;
    wire N__20742;
    wire N__20739;
    wire N__20736;
    wire N__20733;
    wire N__20730;
    wire N__20727;
    wire N__20724;
    wire N__20721;
    wire N__20718;
    wire N__20715;
    wire N__20712;
    wire N__20709;
    wire N__20706;
    wire N__20703;
    wire N__20700;
    wire N__20697;
    wire N__20694;
    wire N__20691;
    wire N__20688;
    wire N__20685;
    wire N__20682;
    wire N__20679;
    wire N__20676;
    wire N__20673;
    wire N__20670;
    wire N__20667;
    wire N__20664;
    wire N__20661;
    wire N__20658;
    wire N__20655;
    wire N__20652;
    wire N__20649;
    wire N__20646;
    wire N__20643;
    wire N__20640;
    wire N__20637;
    wire N__20634;
    wire N__20631;
    wire N__20628;
    wire N__20625;
    wire N__20624;
    wire N__20621;
    wire N__20620;
    wire N__20619;
    wire N__20616;
    wire N__20613;
    wire N__20612;
    wire N__20609;
    wire N__20606;
    wire N__20601;
    wire N__20598;
    wire N__20595;
    wire N__20592;
    wire N__20589;
    wire N__20580;
    wire N__20577;
    wire N__20576;
    wire N__20573;
    wire N__20570;
    wire N__20567;
    wire N__20562;
    wire N__20561;
    wire N__20558;
    wire N__20557;
    wire N__20554;
    wire N__20551;
    wire N__20548;
    wire N__20547;
    wire N__20544;
    wire N__20539;
    wire N__20536;
    wire N__20531;
    wire N__20526;
    wire N__20525;
    wire N__20522;
    wire N__20521;
    wire N__20518;
    wire N__20517;
    wire N__20514;
    wire N__20513;
    wire N__20510;
    wire N__20507;
    wire N__20504;
    wire N__20501;
    wire N__20498;
    wire N__20495;
    wire N__20490;
    wire N__20487;
    wire N__20478;
    wire N__20475;
    wire N__20474;
    wire N__20471;
    wire N__20468;
    wire N__20463;
    wire N__20460;
    wire N__20457;
    wire N__20454;
    wire N__20453;
    wire N__20450;
    wire N__20447;
    wire N__20442;
    wire N__20439;
    wire N__20438;
    wire N__20435;
    wire N__20432;
    wire N__20431;
    wire N__20428;
    wire N__20425;
    wire N__20424;
    wire N__20421;
    wire N__20418;
    wire N__20415;
    wire N__20412;
    wire N__20409;
    wire N__20404;
    wire N__20397;
    wire N__20396;
    wire N__20395;
    wire N__20392;
    wire N__20389;
    wire N__20386;
    wire N__20383;
    wire N__20380;
    wire N__20379;
    wire N__20376;
    wire N__20373;
    wire N__20370;
    wire N__20367;
    wire N__20364;
    wire N__20359;
    wire N__20352;
    wire N__20349;
    wire N__20346;
    wire N__20343;
    wire N__20340;
    wire N__20339;
    wire N__20336;
    wire N__20333;
    wire N__20332;
    wire N__20327;
    wire N__20324;
    wire N__20323;
    wire N__20322;
    wire N__20319;
    wire N__20316;
    wire N__20313;
    wire N__20310;
    wire N__20307;
    wire N__20304;
    wire N__20301;
    wire N__20292;
    wire N__20289;
    wire N__20288;
    wire N__20285;
    wire N__20284;
    wire N__20281;
    wire N__20278;
    wire N__20275;
    wire N__20272;
    wire N__20265;
    wire N__20262;
    wire N__20259;
    wire N__20256;
    wire N__20253;
    wire N__20250;
    wire N__20247;
    wire N__20244;
    wire N__20241;
    wire N__20240;
    wire N__20235;
    wire N__20234;
    wire N__20231;
    wire N__20230;
    wire N__20229;
    wire N__20226;
    wire N__20223;
    wire N__20220;
    wire N__20217;
    wire N__20208;
    wire N__20207;
    wire N__20204;
    wire N__20201;
    wire N__20198;
    wire N__20195;
    wire N__20190;
    wire N__20187;
    wire N__20184;
    wire N__20183;
    wire N__20182;
    wire N__20179;
    wire N__20174;
    wire N__20171;
    wire N__20168;
    wire N__20167;
    wire N__20166;
    wire N__20161;
    wire N__20158;
    wire N__20155;
    wire N__20152;
    wire N__20145;
    wire N__20142;
    wire N__20139;
    wire N__20138;
    wire N__20135;
    wire N__20132;
    wire N__20129;
    wire N__20124;
    wire N__20123;
    wire N__20120;
    wire N__20117;
    wire N__20114;
    wire N__20113;
    wire N__20110;
    wire N__20107;
    wire N__20106;
    wire N__20103;
    wire N__20098;
    wire N__20095;
    wire N__20088;
    wire N__20087;
    wire N__20084;
    wire N__20081;
    wire N__20080;
    wire N__20077;
    wire N__20074;
    wire N__20071;
    wire N__20068;
    wire N__20065;
    wire N__20064;
    wire N__20061;
    wire N__20058;
    wire N__20055;
    wire N__20052;
    wire N__20043;
    wire N__20040;
    wire N__20037;
    wire N__20034;
    wire N__20031;
    wire N__20030;
    wire N__20027;
    wire N__20026;
    wire N__20023;
    wire N__20020;
    wire N__20019;
    wire N__20016;
    wire N__20013;
    wire N__20012;
    wire N__20011;
    wire N__20008;
    wire N__20005;
    wire N__20002;
    wire N__19999;
    wire N__19994;
    wire N__19989;
    wire N__19980;
    wire N__19977;
    wire N__19974;
    wire N__19971;
    wire N__19970;
    wire N__19967;
    wire N__19964;
    wire N__19961;
    wire N__19956;
    wire N__19953;
    wire N__19950;
    wire N__19947;
    wire N__19944;
    wire N__19941;
    wire N__19938;
    wire N__19935;
    wire N__19932;
    wire N__19929;
    wire N__19926;
    wire N__19923;
    wire N__19922;
    wire N__19919;
    wire N__19916;
    wire N__19913;
    wire N__19908;
    wire N__19905;
    wire N__19904;
    wire N__19903;
    wire N__19900;
    wire N__19897;
    wire N__19894;
    wire N__19891;
    wire N__19888;
    wire N__19885;
    wire N__19884;
    wire N__19881;
    wire N__19880;
    wire N__19875;
    wire N__19872;
    wire N__19869;
    wire N__19866;
    wire N__19863;
    wire N__19858;
    wire N__19855;
    wire N__19848;
    wire N__19845;
    wire N__19842;
    wire N__19839;
    wire N__19836;
    wire N__19833;
    wire N__19830;
    wire N__19829;
    wire N__19826;
    wire N__19823;
    wire N__19820;
    wire N__19819;
    wire N__19818;
    wire N__19817;
    wire N__19812;
    wire N__19809;
    wire N__19806;
    wire N__19803;
    wire N__19796;
    wire N__19791;
    wire N__19788;
    wire N__19785;
    wire N__19782;
    wire N__19779;
    wire N__19776;
    wire N__19773;
    wire N__19770;
    wire N__19767;
    wire N__19764;
    wire N__19763;
    wire N__19762;
    wire N__19759;
    wire N__19756;
    wire N__19753;
    wire N__19752;
    wire N__19749;
    wire N__19746;
    wire N__19743;
    wire N__19740;
    wire N__19737;
    wire N__19734;
    wire N__19731;
    wire N__19722;
    wire N__19719;
    wire N__19716;
    wire N__19713;
    wire N__19710;
    wire N__19707;
    wire N__19704;
    wire N__19701;
    wire N__19698;
    wire N__19695;
    wire N__19692;
    wire N__19689;
    wire N__19686;
    wire N__19683;
    wire N__19680;
    wire N__19677;
    wire N__19674;
    wire N__19671;
    wire N__19668;
    wire N__19665;
    wire N__19662;
    wire N__19661;
    wire N__19658;
    wire N__19655;
    wire N__19652;
    wire N__19649;
    wire N__19646;
    wire N__19643;
    wire N__19638;
    wire N__19635;
    wire N__19632;
    wire N__19631;
    wire N__19628;
    wire N__19625;
    wire N__19622;
    wire N__19619;
    wire N__19614;
    wire N__19611;
    wire N__19608;
    wire N__19605;
    wire N__19602;
    wire N__19599;
    wire N__19596;
    wire N__19593;
    wire N__19590;
    wire N__19587;
    wire N__19586;
    wire N__19583;
    wire N__19580;
    wire N__19577;
    wire N__19572;
    wire N__19569;
    wire N__19566;
    wire N__19563;
    wire N__19560;
    wire N__19557;
    wire N__19556;
    wire N__19555;
    wire N__19554;
    wire N__19553;
    wire N__19552;
    wire N__19551;
    wire N__19550;
    wire N__19549;
    wire N__19548;
    wire N__19547;
    wire N__19546;
    wire N__19545;
    wire N__19544;
    wire N__19543;
    wire N__19542;
    wire N__19541;
    wire N__19538;
    wire N__19537;
    wire N__19534;
    wire N__19533;
    wire N__19530;
    wire N__19529;
    wire N__19526;
    wire N__19523;
    wire N__19520;
    wire N__19519;
    wire N__19516;
    wire N__19515;
    wire N__19512;
    wire N__19511;
    wire N__19508;
    wire N__19507;
    wire N__19506;
    wire N__19503;
    wire N__19502;
    wire N__19499;
    wire N__19498;
    wire N__19495;
    wire N__19494;
    wire N__19491;
    wire N__19490;
    wire N__19487;
    wire N__19486;
    wire N__19483;
    wire N__19482;
    wire N__19479;
    wire N__19478;
    wire N__19475;
    wire N__19472;
    wire N__19457;
    wire N__19440;
    wire N__19423;
    wire N__19406;
    wire N__19397;
    wire N__19392;
    wire N__19389;
    wire N__19386;
    wire N__19383;
    wire N__19380;
    wire N__19377;
    wire N__19374;
    wire N__19371;
    wire N__19368;
    wire N__19365;
    wire N__19362;
    wire N__19359;
    wire N__19356;
    wire N__19353;
    wire N__19350;
    wire N__19347;
    wire N__19344;
    wire N__19341;
    wire N__19338;
    wire N__19335;
    wire N__19332;
    wire N__19329;
    wire N__19328;
    wire N__19327;
    wire N__19326;
    wire N__19323;
    wire N__19316;
    wire N__19311;
    wire N__19308;
    wire N__19305;
    wire N__19302;
    wire N__19299;
    wire N__19296;
    wire N__19293;
    wire N__19290;
    wire N__19287;
    wire N__19284;
    wire N__19281;
    wire N__19278;
    wire N__19275;
    wire N__19272;
    wire N__19269;
    wire N__19266;
    wire N__19263;
    wire N__19260;
    wire N__19257;
    wire N__19254;
    wire N__19251;
    wire N__19248;
    wire N__19245;
    wire N__19242;
    wire N__19239;
    wire N__19236;
    wire N__19233;
    wire N__19230;
    wire N__19227;
    wire N__19224;
    wire N__19221;
    wire N__19218;
    wire N__19215;
    wire N__19212;
    wire N__19209;
    wire N__19206;
    wire N__19203;
    wire N__19200;
    wire N__19197;
    wire N__19194;
    wire N__19191;
    wire N__19188;
    wire N__19185;
    wire N__19182;
    wire N__19179;
    wire N__19176;
    wire N__19173;
    wire N__19170;
    wire N__19167;
    wire N__19164;
    wire N__19161;
    wire N__19158;
    wire N__19155;
    wire N__19152;
    wire N__19149;
    wire N__19146;
    wire N__19143;
    wire N__19140;
    wire N__19137;
    wire N__19134;
    wire N__19131;
    wire N__19128;
    wire N__19125;
    wire N__19122;
    wire N__19119;
    wire N__19116;
    wire N__19113;
    wire N__19110;
    wire N__19107;
    wire N__19104;
    wire N__19101;
    wire N__19098;
    wire N__19095;
    wire N__19092;
    wire N__19089;
    wire N__19086;
    wire N__19083;
    wire N__19080;
    wire N__19079;
    wire N__19076;
    wire N__19075;
    wire N__19074;
    wire N__19071;
    wire N__19068;
    wire N__19063;
    wire N__19056;
    wire N__19053;
    wire N__19050;
    wire N__19047;
    wire N__19044;
    wire N__19041;
    wire N__19040;
    wire N__19039;
    wire N__19038;
    wire N__19035;
    wire N__19032;
    wire N__19027;
    wire N__19024;
    wire N__19019;
    wire N__19016;
    wire N__19013;
    wire N__19008;
    wire N__19005;
    wire N__19002;
    wire N__18999;
    wire N__18996;
    wire N__18993;
    wire N__18990;
    wire N__18987;
    wire N__18984;
    wire N__18983;
    wire N__18982;
    wire N__18981;
    wire N__18978;
    wire N__18971;
    wire N__18966;
    wire N__18963;
    wire N__18960;
    wire N__18957;
    wire N__18956;
    wire N__18953;
    wire N__18952;
    wire N__18951;
    wire N__18950;
    wire N__18947;
    wire N__18944;
    wire N__18941;
    wire N__18938;
    wire N__18935;
    wire N__18932;
    wire N__18929;
    wire N__18926;
    wire N__18923;
    wire N__18912;
    wire N__18909;
    wire N__18906;
    wire N__18903;
    wire N__18900;
    wire N__18897;
    wire N__18894;
    wire N__18893;
    wire N__18890;
    wire N__18887;
    wire N__18882;
    wire N__18879;
    wire N__18876;
    wire N__18873;
    wire N__18870;
    wire N__18867;
    wire N__18864;
    wire N__18861;
    wire N__18858;
    wire N__18855;
    wire N__18852;
    wire N__18849;
    wire N__18846;
    wire N__18843;
    wire N__18840;
    wire N__18837;
    wire N__18836;
    wire N__18835;
    wire N__18832;
    wire N__18829;
    wire N__18828;
    wire N__18825;
    wire N__18822;
    wire N__18819;
    wire N__18818;
    wire N__18815;
    wire N__18812;
    wire N__18809;
    wire N__18806;
    wire N__18803;
    wire N__18792;
    wire N__18791;
    wire N__18788;
    wire N__18787;
    wire N__18784;
    wire N__18781;
    wire N__18780;
    wire N__18777;
    wire N__18774;
    wire N__18771;
    wire N__18768;
    wire N__18759;
    wire N__18756;
    wire N__18753;
    wire N__18750;
    wire N__18747;
    wire N__18744;
    wire N__18743;
    wire N__18740;
    wire N__18737;
    wire N__18732;
    wire N__18731;
    wire N__18730;
    wire N__18727;
    wire N__18726;
    wire N__18723;
    wire N__18722;
    wire N__18719;
    wire N__18716;
    wire N__18713;
    wire N__18712;
    wire N__18709;
    wire N__18706;
    wire N__18703;
    wire N__18700;
    wire N__18697;
    wire N__18694;
    wire N__18691;
    wire N__18682;
    wire N__18675;
    wire N__18672;
    wire N__18669;
    wire N__18666;
    wire N__18665;
    wire N__18664;
    wire N__18661;
    wire N__18658;
    wire N__18655;
    wire N__18650;
    wire N__18649;
    wire N__18646;
    wire N__18643;
    wire N__18640;
    wire N__18637;
    wire N__18634;
    wire N__18627;
    wire N__18626;
    wire N__18623;
    wire N__18620;
    wire N__18619;
    wire N__18618;
    wire N__18617;
    wire N__18614;
    wire N__18611;
    wire N__18606;
    wire N__18603;
    wire N__18598;
    wire N__18595;
    wire N__18588;
    wire N__18585;
    wire N__18582;
    wire N__18579;
    wire N__18576;
    wire N__18573;
    wire N__18570;
    wire N__18567;
    wire N__18564;
    wire N__18561;
    wire N__18560;
    wire N__18557;
    wire N__18556;
    wire N__18553;
    wire N__18550;
    wire N__18547;
    wire N__18542;
    wire N__18539;
    wire N__18538;
    wire N__18537;
    wire N__18534;
    wire N__18531;
    wire N__18526;
    wire N__18519;
    wire N__18518;
    wire N__18517;
    wire N__18516;
    wire N__18513;
    wire N__18510;
    wire N__18507;
    wire N__18504;
    wire N__18501;
    wire N__18498;
    wire N__18495;
    wire N__18486;
    wire N__18483;
    wire N__18482;
    wire N__18479;
    wire N__18476;
    wire N__18473;
    wire N__18468;
    wire N__18465;
    wire N__18464;
    wire N__18463;
    wire N__18460;
    wire N__18457;
    wire N__18454;
    wire N__18453;
    wire N__18450;
    wire N__18447;
    wire N__18444;
    wire N__18441;
    wire N__18436;
    wire N__18433;
    wire N__18426;
    wire N__18425;
    wire N__18422;
    wire N__18421;
    wire N__18418;
    wire N__18415;
    wire N__18412;
    wire N__18411;
    wire N__18408;
    wire N__18405;
    wire N__18402;
    wire N__18399;
    wire N__18396;
    wire N__18391;
    wire N__18384;
    wire N__18381;
    wire N__18378;
    wire N__18377;
    wire N__18374;
    wire N__18371;
    wire N__18368;
    wire N__18363;
    wire N__18360;
    wire N__18359;
    wire N__18356;
    wire N__18353;
    wire N__18350;
    wire N__18345;
    wire N__18342;
    wire N__18339;
    wire N__18336;
    wire N__18333;
    wire N__18330;
    wire N__18327;
    wire N__18324;
    wire N__18323;
    wire N__18320;
    wire N__18317;
    wire N__18312;
    wire N__18309;
    wire N__18306;
    wire N__18303;
    wire N__18300;
    wire N__18299;
    wire N__18296;
    wire N__18295;
    wire N__18292;
    wire N__18289;
    wire N__18288;
    wire N__18285;
    wire N__18280;
    wire N__18277;
    wire N__18270;
    wire N__18267;
    wire N__18264;
    wire N__18261;
    wire N__18260;
    wire N__18257;
    wire N__18254;
    wire N__18249;
    wire N__18246;
    wire N__18243;
    wire N__18240;
    wire N__18237;
    wire N__18234;
    wire N__18231;
    wire N__18230;
    wire N__18227;
    wire N__18224;
    wire N__18221;
    wire N__18218;
    wire N__18215;
    wire N__18210;
    wire N__18207;
    wire N__18206;
    wire N__18203;
    wire N__18202;
    wire N__18201;
    wire N__18198;
    wire N__18197;
    wire N__18194;
    wire N__18189;
    wire N__18184;
    wire N__18177;
    wire N__18176;
    wire N__18173;
    wire N__18170;
    wire N__18165;
    wire N__18162;
    wire N__18159;
    wire N__18156;
    wire N__18153;
    wire N__18150;
    wire N__18147;
    wire N__18144;
    wire N__18141;
    wire N__18140;
    wire N__18137;
    wire N__18134;
    wire N__18131;
    wire N__18128;
    wire N__18123;
    wire N__18120;
    wire N__18117;
    wire N__18114;
    wire N__18111;
    wire N__18108;
    wire N__18105;
    wire N__18102;
    wire N__18099;
    wire N__18096;
    wire N__18093;
    wire N__18090;
    wire N__18087;
    wire N__18086;
    wire N__18085;
    wire N__18084;
    wire N__18081;
    wire N__18080;
    wire N__18077;
    wire N__18074;
    wire N__18071;
    wire N__18068;
    wire N__18065;
    wire N__18062;
    wire N__18061;
    wire N__18058;
    wire N__18055;
    wire N__18052;
    wire N__18049;
    wire N__18046;
    wire N__18043;
    wire N__18030;
    wire N__18027;
    wire N__18024;
    wire N__18021;
    wire N__18018;
    wire N__18015;
    wire N__18012;
    wire N__18009;
    wire N__18006;
    wire N__18003;
    wire N__18000;
    wire N__17999;
    wire N__17996;
    wire N__17993;
    wire N__17990;
    wire N__17987;
    wire N__17984;
    wire N__17981;
    wire N__17978;
    wire N__17973;
    wire N__17970;
    wire N__17967;
    wire N__17964;
    wire N__17961;
    wire N__17960;
    wire N__17959;
    wire N__17958;
    wire N__17953;
    wire N__17950;
    wire N__17947;
    wire N__17944;
    wire N__17941;
    wire N__17940;
    wire N__17935;
    wire N__17932;
    wire N__17929;
    wire N__17926;
    wire N__17923;
    wire N__17916;
    wire N__17913;
    wire N__17910;
    wire N__17909;
    wire N__17906;
    wire N__17903;
    wire N__17898;
    wire N__17895;
    wire N__17892;
    wire N__17889;
    wire N__17886;
    wire N__17883;
    wire N__17882;
    wire N__17879;
    wire N__17876;
    wire N__17875;
    wire N__17870;
    wire N__17869;
    wire N__17866;
    wire N__17863;
    wire N__17860;
    wire N__17853;
    wire N__17850;
    wire N__17847;
    wire N__17844;
    wire N__17841;
    wire N__17838;
    wire N__17835;
    wire N__17832;
    wire N__17829;
    wire N__17828;
    wire N__17825;
    wire N__17822;
    wire N__17819;
    wire N__17818;
    wire N__17817;
    wire N__17814;
    wire N__17811;
    wire N__17806;
    wire N__17799;
    wire N__17796;
    wire N__17793;
    wire N__17792;
    wire N__17789;
    wire N__17784;
    wire N__17781;
    wire N__17778;
    wire N__17775;
    wire N__17772;
    wire N__17769;
    wire N__17766;
    wire N__17763;
    wire N__17760;
    wire N__17757;
    wire N__17756;
    wire N__17753;
    wire N__17750;
    wire N__17745;
    wire N__17742;
    wire N__17739;
    wire N__17736;
    wire N__17733;
    wire N__17730;
    wire N__17727;
    wire N__17724;
    wire N__17721;
    wire N__17718;
    wire N__17715;
    wire N__17712;
    wire N__17709;
    wire N__17706;
    wire N__17703;
    wire N__17700;
    wire N__17697;
    wire N__17694;
    wire N__17691;
    wire N__17688;
    wire N__17685;
    wire N__17682;
    wire N__17679;
    wire N__17676;
    wire N__17673;
    wire N__17672;
    wire N__17671;
    wire N__17670;
    wire N__17667;
    wire N__17664;
    wire N__17663;
    wire N__17660;
    wire N__17657;
    wire N__17654;
    wire N__17651;
    wire N__17648;
    wire N__17645;
    wire N__17640;
    wire N__17637;
    wire N__17628;
    wire N__17625;
    wire N__17624;
    wire N__17621;
    wire N__17618;
    wire N__17613;
    wire N__17610;
    wire N__17609;
    wire N__17606;
    wire N__17603;
    wire N__17598;
    wire N__17595;
    wire N__17592;
    wire N__17589;
    wire N__17588;
    wire N__17587;
    wire N__17584;
    wire N__17581;
    wire N__17578;
    wire N__17577;
    wire N__17576;
    wire N__17571;
    wire N__17568;
    wire N__17563;
    wire N__17556;
    wire N__17553;
    wire N__17550;
    wire N__17547;
    wire N__17544;
    wire N__17541;
    wire N__17540;
    wire N__17537;
    wire N__17534;
    wire N__17533;
    wire N__17530;
    wire N__17529;
    wire N__17526;
    wire N__17523;
    wire N__17520;
    wire N__17517;
    wire N__17514;
    wire N__17505;
    wire N__17502;
    wire N__17501;
    wire N__17498;
    wire N__17495;
    wire N__17490;
    wire N__17487;
    wire N__17484;
    wire N__17481;
    wire N__17478;
    wire N__17477;
    wire N__17474;
    wire N__17471;
    wire N__17468;
    wire N__17465;
    wire N__17460;
    wire N__17457;
    wire N__17456;
    wire N__17453;
    wire N__17450;
    wire N__17447;
    wire N__17444;
    wire N__17443;
    wire N__17442;
    wire N__17441;
    wire N__17438;
    wire N__17435;
    wire N__17428;
    wire N__17421;
    wire N__17418;
    wire N__17415;
    wire N__17414;
    wire N__17411;
    wire N__17408;
    wire N__17403;
    wire N__17402;
    wire N__17399;
    wire N__17396;
    wire N__17393;
    wire N__17388;
    wire N__17385;
    wire N__17382;
    wire N__17381;
    wire N__17378;
    wire N__17375;
    wire N__17370;
    wire N__17367;
    wire N__17364;
    wire N__17361;
    wire N__17358;
    wire N__17355;
    wire N__17352;
    wire N__17349;
    wire N__17346;
    wire N__17343;
    wire N__17340;
    wire N__17337;
    wire N__17334;
    wire N__17331;
    wire N__17328;
    wire N__17327;
    wire N__17324;
    wire N__17321;
    wire N__17318;
    wire N__17313;
    wire N__17312;
    wire N__17309;
    wire N__17306;
    wire N__17303;
    wire N__17298;
    wire N__17295;
    wire N__17292;
    wire N__17289;
    wire N__17286;
    wire N__17285;
    wire N__17282;
    wire N__17279;
    wire N__17274;
    wire N__17273;
    wire N__17272;
    wire N__17271;
    wire N__17266;
    wire N__17265;
    wire N__17262;
    wire N__17259;
    wire N__17256;
    wire N__17253;
    wire N__17250;
    wire N__17241;
    wire N__17238;
    wire N__17235;
    wire N__17232;
    wire N__17229;
    wire N__17226;
    wire N__17223;
    wire N__17220;
    wire N__17217;
    wire N__17214;
    wire N__17211;
    wire N__17208;
    wire N__17205;
    wire N__17202;
    wire N__17199;
    wire N__17196;
    wire N__17193;
    wire N__17190;
    wire N__17187;
    wire N__17184;
    wire N__17181;
    wire N__17178;
    wire N__17175;
    wire N__17172;
    wire N__17169;
    wire N__17166;
    wire N__17163;
    wire N__17160;
    wire N__17157;
    wire N__17156;
    wire N__17153;
    wire N__17150;
    wire N__17147;
    wire N__17144;
    wire N__17139;
    wire N__17136;
    wire N__17133;
    wire N__17130;
    wire N__17127;
    wire N__17124;
    wire N__17121;
    wire N__17118;
    wire N__17115;
    wire N__17112;
    wire N__17109;
    wire N__17106;
    wire N__17105;
    wire N__17104;
    wire N__17103;
    wire N__17100;
    wire N__17097;
    wire N__17092;
    wire N__17085;
    wire N__17082;
    wire N__17079;
    wire N__17076;
    wire N__17073;
    wire N__17070;
    wire N__17067;
    wire N__17064;
    wire N__17061;
    wire N__17058;
    wire N__17055;
    wire N__17052;
    wire N__17049;
    wire N__17046;
    wire N__17043;
    wire N__17040;
    wire N__17037;
    wire N__17034;
    wire N__17031;
    wire N__17028;
    wire N__17025;
    wire N__17022;
    wire N__17019;
    wire N__17016;
    wire N__17013;
    wire N__17010;
    wire N__17007;
    wire N__17004;
    wire N__17001;
    wire N__16998;
    wire N__16995;
    wire N__16992;
    wire N__16989;
    wire N__16986;
    wire N__16983;
    wire N__16980;
    wire N__16979;
    wire N__16976;
    wire N__16973;
    wire N__16970;
    wire N__16967;
    wire N__16962;
    wire N__16961;
    wire N__16960;
    wire N__16959;
    wire N__16956;
    wire N__16953;
    wire N__16948;
    wire N__16945;
    wire N__16938;
    wire N__16937;
    wire N__16934;
    wire N__16933;
    wire N__16932;
    wire N__16927;
    wire N__16922;
    wire N__16919;
    wire N__16914;
    wire N__16911;
    wire N__16908;
    wire N__16905;
    wire N__16902;
    wire N__16899;
    wire N__16898;
    wire N__16895;
    wire N__16892;
    wire N__16891;
    wire N__16890;
    wire N__16887;
    wire N__16884;
    wire N__16881;
    wire N__16878;
    wire N__16871;
    wire N__16866;
    wire N__16863;
    wire N__16860;
    wire N__16857;
    wire N__16854;
    wire N__16851;
    wire N__16848;
    wire N__16845;
    wire N__16842;
    wire N__16841;
    wire N__16838;
    wire N__16835;
    wire N__16830;
    wire N__16827;
    wire N__16824;
    wire N__16821;
    wire N__16818;
    wire N__16815;
    wire N__16812;
    wire N__16811;
    wire N__16808;
    wire N__16805;
    wire N__16802;
    wire N__16799;
    wire N__16796;
    wire N__16791;
    wire N__16788;
    wire N__16785;
    wire N__16782;
    wire N__16779;
    wire N__16776;
    wire N__16773;
    wire N__16770;
    wire N__16767;
    wire N__16764;
    wire N__16761;
    wire N__16758;
    wire N__16755;
    wire N__16752;
    wire N__16749;
    wire N__16746;
    wire N__16743;
    wire N__16740;
    wire N__16739;
    wire N__16738;
    wire N__16735;
    wire N__16730;
    wire N__16727;
    wire N__16722;
    wire N__16719;
    wire N__16716;
    wire N__16713;
    wire N__16710;
    wire N__16707;
    wire N__16704;
    wire N__16701;
    wire N__16698;
    wire N__16695;
    wire N__16692;
    wire N__16689;
    wire N__16686;
    wire N__16683;
    wire N__16682;
    wire N__16679;
    wire N__16676;
    wire N__16673;
    wire N__16670;
    wire N__16665;
    wire N__16662;
    wire N__16659;
    wire N__16656;
    wire N__16653;
    wire N__16650;
    wire N__16647;
    wire N__16644;
    wire N__16641;
    wire N__16638;
    wire N__16635;
    wire N__16632;
    wire N__16629;
    wire N__16626;
    wire N__16623;
    wire N__16620;
    wire N__16617;
    wire N__16614;
    wire N__16611;
    wire N__16608;
    wire N__16605;
    wire N__16602;
    wire N__16599;
    wire N__16596;
    wire N__16593;
    wire N__16592;
    wire N__16591;
    wire N__16586;
    wire N__16583;
    wire N__16578;
    wire N__16577;
    wire N__16574;
    wire N__16571;
    wire N__16568;
    wire N__16563;
    wire N__16560;
    wire N__16557;
    wire N__16554;
    wire N__16551;
    wire N__16548;
    wire N__16545;
    wire N__16542;
    wire N__16539;
    wire N__16536;
    wire N__16533;
    wire N__16530;
    wire N__16527;
    wire N__16524;
    wire N__16521;
    wire N__16518;
    wire N__16515;
    wire N__16512;
    wire N__16509;
    wire N__16506;
    wire N__16503;
    wire N__16500;
    wire N__16497;
    wire N__16494;
    wire N__16491;
    wire N__16488;
    wire N__16485;
    wire N__16482;
    wire N__16479;
    wire N__16476;
    wire N__16473;
    wire N__16470;
    wire N__16467;
    wire N__16464;
    wire N__16461;
    wire N__16458;
    wire CLK_pad_gb_input;
    wire VCCG0;
    wire GNDG0;
    wire \c0.n17610_cascade_ ;
    wire \c0.n18214 ;
    wire \c0.n18217 ;
    wire \c0.n18094_cascade_ ;
    wire \c0.n18097_cascade_ ;
    wire \c0.n18262_cascade_ ;
    wire \c0.n22_adj_2365 ;
    wire \c0.n18265_cascade_ ;
    wire \c0.n10468_cascade_ ;
    wire \c0.n14 ;
    wire \c0.n15_cascade_ ;
    wire \c0.data_out_frame2_20_5 ;
    wire \c0.n17306_cascade_ ;
    wire data_out_frame2_18_5;
    wire \c0.n24_cascade_ ;
    wire \c0.n22 ;
    wire \c0.n17174 ;
    wire \c0.n17174_cascade_ ;
    wire \c0.n10356_cascade_ ;
    wire \c0.n18139 ;
    wire \c0.n5_adj_2315_cascade_ ;
    wire data_out_frame2_13_7;
    wire \c0.n18022 ;
    wire \c0.n5_adj_2353_cascade_ ;
    wire \c0.n6 ;
    wire \c0.n6_adj_2138 ;
    wire \c0.n17440 ;
    wire \c0.n18037_cascade_ ;
    wire \c0.n18274_cascade_ ;
    wire \c0.data_out_frame2_20_4 ;
    wire \c0.n18277_cascade_ ;
    wire \c0.n22_adj_2367 ;
    wire \c0.n18034 ;
    wire \c0.n17225 ;
    wire \c0.n17135_cascade_ ;
    wire \c0.n21_cascade_ ;
    wire \c0.n20_adj_2223 ;
    wire \c0.n19_adj_2224 ;
    wire \c0.n14_adj_2308_cascade_ ;
    wire \c0.n17135 ;
    wire \c0.n17092_cascade_ ;
    wire \c0.n17_adj_2294_cascade_ ;
    wire \c0.data_out_frame2_19_4 ;
    wire \c0.n12 ;
    wire data_out_frame2_14_0;
    wire \c0.n17237_cascade_ ;
    wire \c0.n16_adj_2293 ;
    wire \c0.n18136 ;
    wire \c0.data_out_frame2_19_2 ;
    wire \c0.n10520_cascade_ ;
    wire \c0.n10349 ;
    wire \c0.n10462 ;
    wire \c0.n15_adj_2312 ;
    wire \c0.n17285 ;
    wire \c0.n10530 ;
    wire \c0.n10530_cascade_ ;
    wire \c0.n10371 ;
    wire data_out_frame2_7_0;
    wire data_out_frame2_6_0;
    wire \c0.n5_adj_2343 ;
    wire data_out_frame2_15_5;
    wire \c0.n18100_cascade_ ;
    wire \c0.n18103 ;
    wire \c0.n18010_cascade_ ;
    wire \c0.n18013_cascade_ ;
    wire \c0.n22_adj_2375 ;
    wire \c0.n18025 ;
    wire \c0.n18238_cascade_ ;
    wire \c0.n18241 ;
    wire data_out_frame2_7_7;
    wire \c0.n5_adj_2137 ;
    wire \c0.n18154 ;
    wire \c0.n18130_cascade_ ;
    wire \c0.data_out_frame2_20_7 ;
    wire \c0.n18133_cascade_ ;
    wire \c0.n22_adj_2363 ;
    wire \c0.n18028 ;
    wire \c0.n18040_cascade_ ;
    wire \c0.n6_adj_2215 ;
    wire \c0.n17219 ;
    wire \c0.n17141 ;
    wire \c0.n17219_cascade_ ;
    wire \c0.n17_cascade_ ;
    wire \c0.n17228 ;
    wire \c0.n17246_cascade_ ;
    wire \c0.n17187 ;
    wire \c0.n33_cascade_ ;
    wire \c0.data_out_frame2_19_7 ;
    wire \c0.n30_adj_2218 ;
    wire \c0.n17300_cascade_ ;
    wire \c0.n34 ;
    wire \c0.n17237 ;
    wire \c0.n10440 ;
    wire \c0.n17569 ;
    wire data_out_frame2_17_5;
    wire \c0.n17138 ;
    wire \c0.n6_adj_2228_cascade_ ;
    wire \c0.n17312 ;
    wire data_out_frame2_14_3;
    wire \c0.n17267 ;
    wire data_out_frame2_13_2;
    wire \c0.n17309 ;
    wire \c0.n17291 ;
    wire \c0.n17303 ;
    wire \c0.n25 ;
    wire \c0.n28_adj_2200_cascade_ ;
    wire \c0.n27_adj_2204 ;
    wire \c0.n10223_cascade_ ;
    wire \c0.n6_adj_2318 ;
    wire data_out_frame2_9_1;
    wire \c0.n10346 ;
    wire \c0.n17231 ;
    wire \c0.n18076 ;
    wire data_out_frame2_9_5;
    wire \c0.n18109 ;
    wire data_out_frame2_6_3;
    wire \c0.n10334_cascade_ ;
    wire \c0.n10533 ;
    wire \c0.n10_adj_2297 ;
    wire \c0.n14_adj_2296_cascade_ ;
    wire tx2_enable;
    wire \c0.n3_adj_2232 ;
    wire \c0.n3_adj_2278 ;
    wire \c0.n3_adj_2266 ;
    wire \c0.data_out_frame2_19_6 ;
    wire \c0.n18178_cascade_ ;
    wire \c0.n6_adj_2161 ;
    wire \c0.n18181 ;
    wire data_out_frame2_16_6;
    wire \c0.n18112 ;
    wire data_out_frame2_17_6;
    wire \c0.data_out_frame2_20_6 ;
    wire \c0.n18115_cascade_ ;
    wire \c0.n22_adj_2364 ;
    wire data_out_frame2_18_6;
    wire \c0.n18031 ;
    wire \c0.n10548 ;
    wire \c0.n10437 ;
    wire \c0.n17249_cascade_ ;
    wire \c0.n12_adj_2298 ;
    wire data_out_frame2_8_1;
    wire \c0.n20 ;
    wire \c0.n17678 ;
    wire \c0.n17279 ;
    wire \c0.data_out_frame2_20_1 ;
    wire data_out_frame2_13_0;
    wire \c0.n10424 ;
    wire \c0.n14_adj_2346 ;
    wire \c0.n15_adj_2341_cascade_ ;
    wire data_out_frame2_14_5;
    wire \c0.n16_adj_2320_cascade_ ;
    wire \c0.n17216 ;
    wire \c0.data_out_frame2_19_1 ;
    wire \c0.n18058 ;
    wire \c0.n6_adj_2175_cascade_ ;
    wire \c0.n17258 ;
    wire data_out_frame2_11_2;
    wire \c0.n17171 ;
    wire \c0.n17132 ;
    wire \c0.n17184 ;
    wire \c0.n32 ;
    wire data_out_frame2_18_4;
    wire data_out_frame2_5_5;
    wire data_out_frame2_7_3;
    wire data_out_frame2_17_4;
    wire data_out_frame2_17_7;
    wire \c0.n10356 ;
    wire \c0.n10572 ;
    wire \c0.n16_adj_2170 ;
    wire data_out_frame2_6_5;
    wire data_out_frame2_6_7;
    wire data_out_frame2_16_1;
    wire \c0.n17153 ;
    wire \c0.n17168 ;
    wire \c0.n17153_cascade_ ;
    wire \c0.n26_adj_2203 ;
    wire data_out_frame2_5_7;
    wire data_out_frame2_13_3;
    wire data_out_frame2_7_6;
    wire data_out_frame2_6_4;
    wire \c0.n6_adj_2339 ;
    wire \c0.n10507 ;
    wire data_out_frame2_15_0;
    wire \c0.n17273 ;
    wire data_out_frame2_9_2;
    wire \c0.n18046 ;
    wire \c0.n17165 ;
    wire \c0.n10334 ;
    wire \c0.n10223 ;
    wire \c0.n10_adj_2190 ;
    wire \c0.n3_adj_2282 ;
    wire \c0.n3_adj_2227 ;
    wire \c0.n3_adj_2179 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_0 ;
    wire bfn_4_27_0_;
    wire \c0.FRAME_MATCHER_i_31_N_1278_1 ;
    wire \c0.n16079 ;
    wire \c0.n16080 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_3 ;
    wire \c0.FRAME_MATCHER_i_3 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_3 ;
    wire \c0.n16081 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_4 ;
    wire \c0.FRAME_MATCHER_i_4 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_4 ;
    wire \c0.n16082 ;
    wire \c0.n43 ;
    wire \c0.FRAME_MATCHER_i_5 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_5 ;
    wire \c0.n16083 ;
    wire \c0.n16084 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_7 ;
    wire \c0.n16085 ;
    wire \c0.n16086 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_8 ;
    wire bfn_4_28_0_;
    wire \c0.n16087 ;
    wire \c0.n16088 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_11 ;
    wire \c0.n16089 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_12 ;
    wire \c0.n16090 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_13 ;
    wire \c0.n16091 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_14 ;
    wire \c0.n16092 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_15 ;
    wire \c0.n16093 ;
    wire \c0.n16094 ;
    wire bfn_4_29_0_;
    wire \c0.n16095 ;
    wire \c0.n16096 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_19 ;
    wire \c0.n16097 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_20 ;
    wire \c0.n16098 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_21 ;
    wire \c0.n16099 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_22 ;
    wire \c0.n16100 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_23 ;
    wire \c0.n16101 ;
    wire \c0.n16102 ;
    wire bfn_4_30_0_;
    wire \c0.n16103 ;
    wire \c0.n16104 ;
    wire \c0.n16105 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_28 ;
    wire \c0.n16106 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_29 ;
    wire \c0.FRAME_MATCHER_i_29 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_29 ;
    wire \c0.n16107 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_30 ;
    wire \c0.n16108 ;
    wire \c0.n16109 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_31 ;
    wire n5244_cascade_;
    wire n11018_cascade_;
    wire \c0.n18008 ;
    wire n13692_cascade_;
    wire bfn_4_32_0_;
    wire \c0.rx.n16125 ;
    wire \c0.rx.n16126 ;
    wire \c0.rx.n16127 ;
    wire \c0.rx.n16128 ;
    wire \c0.rx.n16129 ;
    wire \c0.rx.n16130 ;
    wire \c0.rx.n16131 ;
    wire data_out_frame2_18_1;
    wire data_out_frame2_5_6;
    wire \c0.n14_adj_2188_cascade_ ;
    wire \c0.n15_adj_2185 ;
    wire \c0.data_out_frame2_20_2 ;
    wire data_out_frame2_7_4;
    wire \c0.n17240 ;
    wire \c0.n17240_cascade_ ;
    wire \c0.n14_adj_2206 ;
    wire \c0.n17439 ;
    wire \c0.n17249 ;
    wire \c0.data_out_frame2_19_5 ;
    wire \c0.n17116 ;
    wire \c0.n17234 ;
    wire \c0.n15_adj_2291 ;
    wire \c0.n17288 ;
    wire data_out_frame2_12_4;
    wire \c0.n17288_cascade_ ;
    wire \c0.n14_adj_2292 ;
    wire \c0.n17294 ;
    wire \c0.n10428_cascade_ ;
    wire \c0.n12_adj_2178 ;
    wire \c0.n10504 ;
    wire data_out_frame2_17_1;
    wire data_out_frame2_9_4;
    wire \c0.n17568 ;
    wire \c0.n10554 ;
    wire \c0.n10263 ;
    wire \c0.n15_adj_2205 ;
    wire \c0.n5_adj_2337 ;
    wire data_out_frame2_10_2;
    wire \c0.n10492 ;
    wire data_out_frame2_12_5;
    wire \c0.n17255 ;
    wire data_out_frame2_16_4;
    wire data_out_frame2_11_1;
    wire \c0.n17156 ;
    wire \c0.n6_adj_2182_cascade_ ;
    wire \c0.n10229 ;
    wire n10725_cascade_;
    wire data_out_frame2_12_7;
    wire data_out_frame2_10_3;
    wire \c0.n18106 ;
    wire data_out_frame2_16_2;
    wire data_out_frame2_15_2;
    wire data_out_frame2_18_2;
    wire data_out_frame2_16_5;
    wire data_out_frame2_15_4;
    wire bfn_5_23_0_;
    wire n15979;
    wire n15980;
    wire n15981;
    wire n15982;
    wire n15983;
    wire n15984;
    wire n15985;
    wire n15986;
    wire bfn_5_24_0_;
    wire n15987;
    wire n15988;
    wire n15989;
    wire n15990;
    wire n15991;
    wire n15992;
    wire n15993;
    wire n15994;
    wire bfn_5_25_0_;
    wire n15995;
    wire n15996;
    wire n15997;
    wire n15998;
    wire n15999;
    wire n16000;
    wire n16001;
    wire n16002;
    wire bfn_5_26_0_;
    wire n16003;
    wire n16004;
    wire n16005;
    wire n16006;
    wire n16007;
    wire n16008;
    wire n16009;
    wire \c0.n3 ;
    wire \c0.n26_adj_2373_cascade_ ;
    wire \c0.n3_adj_2280 ;
    wire \c0.FRAME_MATCHER_i_6 ;
    wire \c0.n41 ;
    wire \c0.n3_adj_2261 ;
    wire \c0.n3_adj_2270 ;
    wire \c0.n3_adj_2252 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_17 ;
    wire \c0.n3_adj_2257 ;
    wire \c0.FRAME_MATCHER_i_17 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_17 ;
    wire \c0.n3_adj_2248 ;
    wire \c0.n3_adj_2250 ;
    wire \c0.n3_adj_2244 ;
    wire \c0.FRAME_MATCHER_i_21 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_21 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_27 ;
    wire \c0.n3_adj_2276 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_8 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_9 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_31 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_25 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_26 ;
    wire \c0.rx.n10845 ;
    wire n1;
    wire \c0.rx.r_Clock_Count_4 ;
    wire \c0.rx.r_Clock_Count_1 ;
    wire \c0.rx.n10656 ;
    wire n17708_cascade_;
    wire n5244;
    wire n11018;
    wire \c0.data_out_frame2_20_0 ;
    wire \c0.n18049 ;
    wire \c0.n18043 ;
    wire \c0.n17586 ;
    wire \c0.n18244_cascade_ ;
    wire \c0.n6_adj_2140 ;
    wire \c0.tx2.r_Tx_Data_1 ;
    wire \c0.tx2.n18232_cascade_ ;
    wire \c0.n22_adj_2387 ;
    wire \c0.tx2.r_Tx_Data_0 ;
    wire \c0.n18157 ;
    wire \c0.n17603 ;
    wire \c0.n18226_cascade_ ;
    wire \c0.n18229 ;
    wire data_out_frame2_10_0;
    wire \c0.n18148_cascade_ ;
    wire \c0.n18151 ;
    wire data_out_frame2_5_0;
    wire \c0.n5_adj_2217 ;
    wire \c0.n6_adj_2143 ;
    wire \c0.data_out_frame2_19_3 ;
    wire \c0.n18052_cascade_ ;
    wire \c0.data_out_frame2_20_3 ;
    wire \c0.n18055_cascade_ ;
    wire \c0.n9157 ;
    wire \c0.n18061 ;
    wire \c0.n18256_cascade_ ;
    wire \c0.n6_adj_2139 ;
    wire \c0.n22_adj_2371 ;
    wire \c0.n18259_cascade_ ;
    wire \c0.tx2.r_Tx_Data_3 ;
    wire data_out_frame2_10_1;
    wire \c0.n17203 ;
    wire data_out_frame2_8_6;
    wire data_out_frame2_9_6;
    wire \c0.n18127 ;
    wire data_out_frame2_18_3;
    wire data_out_frame2_17_0;
    wire \c0.n18163 ;
    wire \c0.n18208 ;
    wire data_out_frame2_17_3;
    wire data_out_frame2_14_2;
    wire \c0.n10_adj_2207 ;
    wire data_out_frame2_11_4;
    wire data_out_frame2_11_5;
    wire \c0.n10359 ;
    wire data_out_frame2_5_4;
    wire data_out_frame2_10_7;
    wire \c0.tx2.n13748_cascade_ ;
    wire data_out_frame2_18_7;
    wire data_out_frame2_17_2;
    wire data_out_frame2_7_5;
    wire \c0.tx2.n10 ;
    wire tx2_o;
    wire data_out_frame2_14_7;
    wire \c0.tx2.n17322 ;
    wire \c0.tx2.n17018 ;
    wire \c0.tx2.r_Clock_Count_0 ;
    wire bfn_6_24_0_;
    wire \c0.tx2.r_Clock_Count_1 ;
    wire \c0.tx2.n16132 ;
    wire \c0.tx2.r_Clock_Count_2 ;
    wire \c0.tx2.n16133 ;
    wire \c0.tx2.r_Clock_Count_3 ;
    wire \c0.tx2.n16134 ;
    wire \c0.tx2.r_Clock_Count_4 ;
    wire \c0.tx2.n16135 ;
    wire \c0.tx2.r_Clock_Count_5 ;
    wire \c0.tx2.n16136 ;
    wire \c0.tx2.r_Clock_Count_6 ;
    wire \c0.tx2.n16137 ;
    wire \c0.tx2.r_Clock_Count_7 ;
    wire \c0.tx2.n16138 ;
    wire \c0.tx2.n16139 ;
    wire bfn_6_25_0_;
    wire \c0.tx2.r_Clock_Count_8 ;
    wire \c0.tx2.n10852 ;
    wire \c0.FRAME_MATCHER_i_8 ;
    wire \c0.n42 ;
    wire \c0.n41_adj_2376_cascade_ ;
    wire \c0.n39_adj_2377 ;
    wire \c0.n43_adj_2380 ;
    wire \c0.n48_adj_2379_cascade_ ;
    wire \c0.n44_adj_2378 ;
    wire \c0.n9995_cascade_ ;
    wire \c0.n9995 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_2 ;
    wire \c0.n3_adj_2286 ;
    wire \c0.n3_adj_2226 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_2 ;
    wire \c0.n40 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_24 ;
    wire \c0.n3_adj_2242 ;
    wire \c0.n3_adj_2240 ;
    wire \c0.n3_adj_2234 ;
    wire \c0.n3_adj_2230 ;
    wire \c0.n10009_cascade_ ;
    wire \c0.n3_adj_2181 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_18 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_27 ;
    wire \c0.FRAME_MATCHER_i_27 ;
    wire \c0.n3_adj_2236 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_9 ;
    wire \c0.FRAME_MATCHER_i_9 ;
    wire \c0.n3_adj_2274 ;
    wire \c0.rx.n17636 ;
    wire n17707;
    wire \c0.rx.r_Clock_Count_2 ;
    wire \c0.rx.r_Clock_Count_0 ;
    wire \c0.rx.r_Clock_Count_3 ;
    wire \c0.rx.n6 ;
    wire \c0.rx.n17022_cascade_ ;
    wire \c0.rx.r_SM_Main_2_N_2094_0_cascade_ ;
    wire \c0.rx.n17380_cascade_ ;
    wire \c0.rx.n17635 ;
    wire \c0.rx.r_SM_Main_2_N_2094_0 ;
    wire \c0.rx.n6_adj_2130 ;
    wire \c0.n18247 ;
    wire \c0.n22_adj_2372 ;
    wire \c0.tx2.r_Tx_Data_2 ;
    wire \c0.n17620 ;
    wire \c0.tx2.r_Tx_Data_6 ;
    wire \c0.tx2.r_Tx_Data_7 ;
    wire \c0.tx2.r_Tx_Data_4 ;
    wire \c0.tx2.n18082_cascade_ ;
    wire \c0.tx2.r_Tx_Data_5 ;
    wire \c0.tx2.n18085_cascade_ ;
    wire \c0.tx2.n18235 ;
    wire \c0.tx2.o_Tx_Serial_N_2062_cascade_ ;
    wire n3;
    wire \c0.tx2.n13614_cascade_ ;
    wire \c0.n17587 ;
    wire \c0.n17107 ;
    wire data_out_frame2_15_6;
    wire data_out_frame2_12_6;
    wire \c0.n18118_cascade_ ;
    wire data_out_frame2_13_6;
    wire \c0.n18121 ;
    wire \c0.tx2.n13614 ;
    wire n10976;
    wire n10976_cascade_;
    wire r_Bit_Index_2_adj_2440;
    wire data_out_frame2_5_1;
    wire \c0.n6_adj_2142 ;
    wire \c0.n18064 ;
    wire \c0.n18067 ;
    wire n8191;
    wire data_out_frame2_6_1;
    wire \c0.n5_adj_2289 ;
    wire data_out_frame2_11_7;
    wire \c0.n10413_cascade_ ;
    wire \c0.n17282 ;
    wire data_out_frame2_10_6;
    wire data_out_frame2_11_6;
    wire \c0.n18124 ;
    wire \c0.data_out_frame2_19_0 ;
    wire data_out_frame2_18_0;
    wire \c0.n18160 ;
    wire \c0.n10563 ;
    wire data_out_frame2_13_5;
    wire \c0.n17095 ;
    wire \c0.n31 ;
    wire data_out_frame2_13_1;
    wire data_out_frame2_12_1;
    wire \c0.n18019 ;
    wire data_out_frame2_12_3;
    wire data_out_frame2_5_3;
    wire \c0.n18142 ;
    wire data_out_frame2_8_7;
    wire data_out_frame2_9_7;
    wire \c0.n18145 ;
    wire \c0.tx2.n9269 ;
    wire data_out_frame2_5_2;
    wire data_out_frame2_10_4;
    wire \c0.n10456 ;
    wire data_out_frame2_10_5;
    wire data_out_frame2_11_3;
    wire data_out_frame2_14_1;
    wire data_out_frame2_15_1;
    wire \c0.n18016 ;
    wire data_out_frame2_12_2;
    wire data_out_frame2_7_2;
    wire data_out_frame2_6_2;
    wire \c0.n5_adj_2290 ;
    wire data_out_frame2_14_4;
    wire data_out_frame2_11_0;
    wire \c0.n17276 ;
    wire n17412;
    wire data_out_frame2_9_3;
    wire \c0.n6_adj_2197 ;
    wire data_out_frame2_15_7;
    wire \c0.n17123 ;
    wire data_out_frame2_14_6;
    wire \c0.n10434 ;
    wire data_out_frame2_16_3;
    wire data_out_frame2_15_3;
    wire \c0.n10482 ;
    wire data_out_frame2_8_4;
    wire data_out_frame2_8_0;
    wire \c0.n10513 ;
    wire data_out_frame2_16_0;
    wire \c0.n17098 ;
    wire data_out_frame2_8_3;
    wire \c0.n17_adj_2321 ;
    wire \c0.n30_cascade_ ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_26 ;
    wire \c0.FRAME_MATCHER_i_25 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_25 ;
    wire \c0.FRAME_MATCHER_i_24 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_24 ;
    wire \c0.FRAME_MATCHER_i_23 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_23 ;
    wire \c0.FRAME_MATCHER_i_20 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_20 ;
    wire \c0.FRAME_MATCHER_i_19 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_19 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_16 ;
    wire \c0.n3_adj_2254 ;
    wire \c0.FRAME_MATCHER_i_18 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_18 ;
    wire \c0.n3_adj_2288 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_1 ;
    wire \c0.n3_adj_2246 ;
    wire \c0.FRAME_MATCHER_i_22 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_22 ;
    wire \c0.FRAME_MATCHER_i_26 ;
    wire \c0.n3_adj_2238 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_10 ;
    wire r_Bit_Index_1_adj_2441;
    wire r_Bit_Index_0_adj_2442;
    wire n5266;
    wire tx_enable;
    wire n10674;
    wire \c0.n17574 ;
    wire \c0.rx.n10620 ;
    wire n17361;
    wire \c0.rx.r_SM_Main_2_N_2088_2 ;
    wire r_SM_Main_1;
    wire \c0.rx.r_SM_Main_2_N_2088_2_cascade_ ;
    wire \c0.rx.r_SM_Main_0 ;
    wire \c0.FRAME_MATCHER_i_31_N_1278_12 ;
    wire \c0.FRAME_MATCHER_i_12 ;
    wire \c0.n3_adj_2268 ;
    wire bfn_9_17_0_;
    wire \c0.n15972 ;
    wire \c0.n15973 ;
    wire \c0.n15974 ;
    wire \c0.n17606 ;
    wire \c0.n15975 ;
    wire \c0.n15976 ;
    wire \c0.n15977 ;
    wire \c0.n15978 ;
    wire \c0.n17714 ;
    wire \c0.n17589 ;
    wire data_out_frame2_7_1;
    wire n10725;
    wire data_out_frame2_12_0;
    wire r_SM_Main_2_N_2031_1;
    wire r_SM_Main_0;
    wire r_SM_Main_2_adj_2438;
    wire n4_adj_2484;
    wire r_SM_Main_1_adj_2439;
    wire data_in_0_3;
    wire \c0.n10133_cascade_ ;
    wire \c0.n6_adj_2356_cascade_ ;
    wire \c0.n10027_cascade_ ;
    wire data_in_0_7;
    wire data_in_1_3;
    wire \c0.n17331_cascade_ ;
    wire \c0.n17410 ;
    wire data_in_2_6;
    wire \c0.n12_adj_2355 ;
    wire data_in_2_4;
    wire \c0.n4_adj_2150 ;
    wire \c0.n10133 ;
    wire \c0.n17406 ;
    wire data_in_0_6;
    wire \c0.FRAME_MATCHER_i_15 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_15 ;
    wire \c0.FRAME_MATCHER_i_13 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_13 ;
    wire \c0.FRAME_MATCHER_i_11 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_11 ;
    wire \c0.FRAME_MATCHER_i_7 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_7 ;
    wire \c0.n37 ;
    wire \c0.FRAME_MATCHER_i_28 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_28 ;
    wire \c0.FRAME_MATCHER_state_13 ;
    wire \c0.n8_adj_2332 ;
    wire \c0.FRAME_MATCHER_state_19 ;
    wire \c0.n8_adj_2328 ;
    wire \c0.FRAME_MATCHER_state_6 ;
    wire \c0.n8_adj_2334 ;
    wire \c0.FRAME_MATCHER_state_12 ;
    wire \c0.n16708 ;
    wire \c0.FRAME_MATCHER_state_14 ;
    wire \c0.n8_adj_2331 ;
    wire data_out_frame2_16_7;
    wire \c0.n17194 ;
    wire \c0.n10459 ;
    wire data_in_0_5;
    wire data_in_0_4;
    wire data_in_0_2;
    wire data_in_1_5;
    wire \c0.FRAME_MATCHER_i_31_N_1278_16 ;
    wire \c0.FRAME_MATCHER_state_4 ;
    wire \c0.n16716 ;
    wire data_in_1_2;
    wire \c0.n17388 ;
    wire \c0.n3_adj_2272 ;
    wire \c0.FRAME_MATCHER_i_10 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_10 ;
    wire \c0.n3_adj_2264 ;
    wire \c0.FRAME_MATCHER_i_14 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_14 ;
    wire \c0.FRAME_MATCHER_i_16 ;
    wire \c0.n10009 ;
    wire \c0.n3_adj_2259 ;
    wire n26_adj_2423;
    wire bfn_9_29_0_;
    wire n25_adj_2424;
    wire n16041;
    wire n24;
    wire n16042;
    wire n23_adj_2425;
    wire n16043;
    wire n22_adj_2426;
    wire n16044;
    wire n21;
    wire n16045;
    wire n20;
    wire n16046;
    wire n19;
    wire n16047;
    wire n16048;
    wire n18;
    wire bfn_9_30_0_;
    wire n17;
    wire n16049;
    wire n16;
    wire n16050;
    wire n15;
    wire n16051;
    wire n14;
    wire n16052;
    wire n13;
    wire n16053;
    wire n12;
    wire n16054;
    wire n11;
    wire n16055;
    wire n16056;
    wire n10_adj_2420;
    wire bfn_9_31_0_;
    wire n9_adj_2421;
    wire n16057;
    wire n8_adj_2412;
    wire n16058;
    wire n7;
    wire n16059;
    wire n6_adj_2429;
    wire n16060;
    wire n16061;
    wire n16062;
    wire n16063;
    wire n16064;
    wire bfn_9_32_0_;
    wire n16065;
    wire \c0.n17711 ;
    wire \c0.n17659 ;
    wire \c0.n11867_cascade_ ;
    wire \c0.n4_adj_2187 ;
    wire \c0.n4_adj_2152 ;
    wire \c0.byte_transmit_counter2_0 ;
    wire \c0.n17761 ;
    wire \c0.byte_transmit_counter2_1 ;
    wire \c0.n4_adj_2155 ;
    wire \c0.data_in_frame_3_6 ;
    wire \c0.n15_adj_2310_cascade_ ;
    wire \c0.data_in_frame_3_3 ;
    wire n17075_cascade_;
    wire data_in_2_5;
    wire data_in_2_0;
    wire \c0.n17400_cascade_ ;
    wire \c0.n8_adj_2359_cascade_ ;
    wire \c0.n13450 ;
    wire \c0.data_in_frame_3_4 ;
    wire data_in_0_1;
    wire \c0.n7_adj_2384_cascade_ ;
    wire \c0.n6_adj_2336 ;
    wire \c0.n10136 ;
    wire data_in_1_4;
    wire data_in_2_3;
    wire \c0.n16_adj_2361_cascade_ ;
    wire \c0.n17_adj_2362 ;
    wire n63_cascade_;
    wire data_in_2_7;
    wire \c0.n10141 ;
    wire \c0.n10027 ;
    wire \c0.n17_adj_2370 ;
    wire \c0.n16_adj_2366_cascade_ ;
    wire data_in_1_7;
    wire n9378_cascade_;
    wire \c0.n47_adj_2347_cascade_ ;
    wire \c0.n13146_cascade_ ;
    wire data_in_3_4;
    wire data_in_1_6;
    wire data_in_3_5;
    wire \c0.n17402 ;
    wire \c0.FRAME_MATCHER_state_20 ;
    wire \c0.n8_adj_2327 ;
    wire \c0.FRAME_MATCHER_i_31 ;
    wire \c0.n10161 ;
    wire n2061_cascade_;
    wire \c0.n47_adj_2347 ;
    wire \c0.n9334_cascade_ ;
    wire \c0.n4 ;
    wire \c0.n15821_cascade_ ;
    wire \c0.n8_adj_2335 ;
    wire rand_data_0;
    wire bfn_10_25_0_;
    wire rand_data_1;
    wire n16010;
    wire rand_data_2;
    wire n16011;
    wire rand_data_3;
    wire n16012;
    wire rand_data_4;
    wire n16013;
    wire rand_data_5;
    wire n16014;
    wire rand_data_6;
    wire n16015;
    wire rand_data_7;
    wire n16016;
    wire n16017;
    wire rand_data_8;
    wire bfn_10_26_0_;
    wire rand_data_9;
    wire rand_setpoint_9;
    wire n16018;
    wire rand_data_10;
    wire n16019;
    wire rand_data_11;
    wire n16020;
    wire rand_data_12;
    wire n16021;
    wire rand_data_13;
    wire n16022;
    wire rand_data_14;
    wire n16023;
    wire rand_data_15;
    wire n16024;
    wire n16025;
    wire rand_data_16;
    wire bfn_10_27_0_;
    wire rand_data_17;
    wire rand_setpoint_17;
    wire n16026;
    wire rand_data_18;
    wire n16027;
    wire rand_data_19;
    wire n16028;
    wire rand_data_20;
    wire n16029;
    wire rand_data_21;
    wire n16030;
    wire rand_data_22;
    wire n16031;
    wire rand_data_23;
    wire n16032;
    wire n16033;
    wire rand_data_24;
    wire rand_setpoint_24;
    wire bfn_10_28_0_;
    wire rand_data_25;
    wire n16034;
    wire rand_data_26;
    wire n16035;
    wire rand_data_27;
    wire n16036;
    wire rand_data_28;
    wire n16037;
    wire rand_data_29;
    wire n16038;
    wire rand_data_30;
    wire n16039;
    wire rand_data_31;
    wire n16040;
    wire rand_setpoint_31;
    wire rand_setpoint_26;
    wire rand_setpoint_29;
    wire rand_setpoint_27;
    wire rand_setpoint_28;
    wire rand_setpoint_11;
    wire \c0.n17585 ;
    wire rand_setpoint_10;
    wire \c0.n17583_cascade_ ;
    wire \c0.rx.r_Clock_Count_5 ;
    wire \c0.rx.n17022 ;
    wire r_SM_Main_2;
    wire \c0.rx.n17058 ;
    wire \c0.rx.r_Clock_Count_7 ;
    wire \c0.rx.r_Clock_Count_6 ;
    wire \c0.rx.n17080 ;
    wire \c0.byte_transmit_counter2_3 ;
    wire \c0.byte_transmit_counter2_4 ;
    wire \c0.n17710 ;
    wire \c0.byte_transmit_counter2_2 ;
    wire \c0.n4_adj_2154 ;
    wire \c0.n4_adj_2345 ;
    wire \c0.n2122_cascade_ ;
    wire \c0.data_in_frame_2_5 ;
    wire \c0.data_in_frame_5_6 ;
    wire \c0.n2124_cascade_ ;
    wire \c0.data_in_frame_5_3 ;
    wire \c0.n16475 ;
    wire \c0.data_in_frame_5_5 ;
    wire \c0.n17373 ;
    wire \c0.n19_adj_2303 ;
    wire \c0.n17076_cascade_ ;
    wire n17075;
    wire data_in_frame_6_4;
    wire \c0.n10215 ;
    wire \c0.data_in_frame_0_4 ;
    wire \c0.n10215_cascade_ ;
    wire \c0.n17206_cascade_ ;
    wire \c0.n20_adj_2195 ;
    wire \c0.n39 ;
    wire \c0.n2137 ;
    wire \c0.n23_cascade_ ;
    wire \c0.n26_adj_2210 ;
    wire \c0.n18 ;
    wire \c0.n30_adj_2213_cascade_ ;
    wire \c0.n17_adj_2214 ;
    wire n31_adj_2415_cascade_;
    wire data_in_frame_6_3;
    wire data_in_3_7;
    wire \c0.n6_adj_2358 ;
    wire \c0.FRAME_MATCHER_i_1 ;
    wire \c0.n15164 ;
    wire \c0.n17072_cascade_ ;
    wire \c0.data_in_frame_2_4 ;
    wire FRAME_MATCHER_i_31__N_1273_cascade_;
    wire n17086_cascade_;
    wire n63_adj_2428;
    wire n63;
    wire \c0.FRAME_MATCHER_state_8 ;
    wire \c0.n16666 ;
    wire \c0.FRAME_MATCHER_state_9 ;
    wire \c0.n16674 ;
    wire \c0.n1034 ;
    wire n10140_cascade_;
    wire \c0.n8_adj_2385_cascade_ ;
    wire \c0.n16670 ;
    wire \c0.n17367_cascade_ ;
    wire n9_cascade_;
    wire \c0.n10139 ;
    wire \c0.n11833 ;
    wire \c0.FRAME_MATCHER_state_3 ;
    wire \c0.FRAME_MATCHER_state_5 ;
    wire n9;
    wire n21_adj_2487_cascade_;
    wire n63_adj_2418;
    wire n6_adj_2410;
    wire n2061;
    wire \c0.n51_adj_2173 ;
    wire \c0.n10166 ;
    wire \c0.FRAME_MATCHER_i_30 ;
    wire \c0.FRAME_MATCHER_i_31_N_1310_30 ;
    wire \c0.n16696 ;
    wire rand_setpoint_2;
    wire rand_setpoint_3;
    wire \c0.FRAME_MATCHER_state_7 ;
    wire \c0.n16141 ;
    wire rand_setpoint_23;
    wire \c0.n17639_cascade_ ;
    wire rand_setpoint_20;
    wire rand_setpoint_22;
    wire \c0.n17647 ;
    wire rand_setpoint_19;
    wire \c0.n17631_cascade_ ;
    wire rand_setpoint_18;
    wire \c0.n17627_cascade_ ;
    wire rand_setpoint_21;
    wire \c0.n17643 ;
    wire \c0.n18268_cascade_ ;
    wire \c0.tx.n55_cascade_ ;
    wire \c0.n5_adj_2136 ;
    wire rand_setpoint_12;
    wire \c0.n5 ;
    wire \c0.n18172_cascade_ ;
    wire \c0.n17764 ;
    wire \c0.n17676 ;
    wire rand_setpoint_14;
    wire \c0.n17703 ;
    wire \c0.data_out_1_4 ;
    wire \c0.n17675 ;
    wire \c0.n17697 ;
    wire n18271;
    wire n10_adj_2408_cascade_;
    wire \c0.data_out_2_3 ;
    wire data_out_0_5;
    wire data_out_2_2;
    wire n2699_cascade_;
    wire data_out_3_4;
    wire n2699;
    wire data_out_3_2;
    wire \c0.data_in_frame_2_6 ;
    wire \c0.n17713 ;
    wire \c0.n4_adj_2325 ;
    wire \c0.tx2_transmit_N_1996 ;
    wire \c0.byte_transmit_counter2_7 ;
    wire \c0.byte_transmit_counter2_6 ;
    wire \c0.n13284 ;
    wire \c0.n13628 ;
    wire \c0.n13628_cascade_ ;
    wire tx2_active;
    wire \c0.data_in_frame_3_2 ;
    wire data_in_frame_6_2;
    wire \c0.n17475_cascade_ ;
    wire \c0.data_out_frame2_0_5 ;
    wire \c0.n16352 ;
    wire \c0.n24_adj_2340 ;
    wire data_in_frame_6_5;
    wire \c0.n2122 ;
    wire \c0.n17469_cascade_ ;
    wire \c0.data_out_frame2_0_7 ;
    wire data_in_frame_6_1;
    wire \c0.data_in_frame_5_1 ;
    wire \c0.n17114_cascade_ ;
    wire \c0.data_in_frame_5_7 ;
    wire \c0.data_in_frame_1_4 ;
    wire \c0.n17101_cascade_ ;
    wire \c0.n10_adj_2299_cascade_ ;
    wire \c0.n17206 ;
    wire \c0.n10407 ;
    wire data_in_frame_6_0;
    wire \c0.n10407_cascade_ ;
    wire \c0.data_in_frame_1_5 ;
    wire \c0.n17215 ;
    wire \c0.n2128 ;
    wire data_in_frame_6_7;
    wire \c0.data_in_frame_5_0 ;
    wire \c0.n2128_cascade_ ;
    wire \c0.n19_adj_2324 ;
    wire data_in_3_0;
    wire \c0.data_in_frame_0_3 ;
    wire \c0.data_in_frame_0_2 ;
    wire \c0.n2120 ;
    wire \c0.n22_adj_2201_cascade_ ;
    wire \c0.n27_adj_2202 ;
    wire \c0.data_in_frame_0_5 ;
    wire \c0.data_in_frame_0_6 ;
    wire \c0.data_in_frame_2_0 ;
    wire data_in_3_6;
    wire data_in_1_0;
    wire data_in_0_0;
    wire data_in_3_1;
    wire data_in_2_1;
    wire data_in_1_1;
    wire \c0.data_in_frame_3_5 ;
    wire \c0.data_in_frame_2_3 ;
    wire rx_data_3;
    wire data_in_3_3;
    wire \c0.FRAME_MATCHER_state_28 ;
    wire \c0.n50 ;
    wire \c0.n47_cascade_ ;
    wire \c0.n49 ;
    wire \c0.n51 ;
    wire \c0.n56_cascade_ ;
    wire \c0.n45 ;
    wire \c0.n10018_cascade_ ;
    wire n5;
    wire n1_adj_2486;
    wire n9378;
    wire FRAME_MATCHER_state_1;
    wire \c0.n16261 ;
    wire \c0.r_SM_Main_2_N_2034_0_adj_2167 ;
    wire \c0.n10018 ;
    wire n10088;
    wire n17086;
    wire n17063;
    wire n17089;
    wire n17090;
    wire n3_adj_2485;
    wire n6;
    wire n17349;
    wire n3_adj_2485_cascade_;
    wire blink_counter_24;
    wire blink_counter_23;
    wire blink_counter_22;
    wire blink_counter_21;
    wire n10140;
    wire n8;
    wire n4_adj_2417_cascade_;
    wire FRAME_MATCHER_state_31_N_1406_2;
    wire FRAME_MATCHER_state_2;
    wire blink_counter_25;
    wire n17428;
    wire n17427;
    wire LED_c;
    wire n3779;
    wire FRAME_MATCHER_i_31__N_1273;
    wire n6_adj_2488;
    wire data_out_3_0;
    wire n18175;
    wire n10_adj_2409_cascade_;
    wire \c0.n8_adj_2183_cascade_ ;
    wire \c0.n17671 ;
    wire rand_setpoint_4;
    wire data_out_10__7__N_110_cascade_;
    wire rand_setpoint_6;
    wire \c0.data_out_1_2 ;
    wire \c0.n17696 ;
    wire n18073_cascade_;
    wire \c0.tx.n10688_cascade_ ;
    wire r_Tx_Data_1;
    wire rand_setpoint_1;
    wire r_Tx_Data_3;
    wire n18070;
    wire \c0.tx.n10688 ;
    wire n4_adj_2419_cascade_;
    wire n5_adj_2407_cascade_;
    wire n10_adj_2444_cascade_;
    wire n8_adj_2447;
    wire n4_adj_2419;
    wire bfn_12_31_0_;
    wire \c0.n27 ;
    wire \c0.n16066 ;
    wire \c0.n16067 ;
    wire \c0.n25_adj_2386 ;
    wire \c0.n16068 ;
    wire \c0.n16069 ;
    wire \c0.n16070 ;
    wire \c0.n22_adj_2313 ;
    wire \c0.n16071 ;
    wire \c0.n21_adj_2262 ;
    wire \c0.n16072 ;
    wire \c0.n16073 ;
    wire bfn_12_32_0_;
    wire \c0.n16074 ;
    wire \c0.n16075 ;
    wire \c0.n16076 ;
    wire \c0.n16077 ;
    wire \c0.n16078 ;
    wire \c0.n10594 ;
    wire \c0.n16353 ;
    wire \c0.n26_adj_2368 ;
    wire \c0.n16474 ;
    wire \c0.n18_adj_2360 ;
    wire rx_data_0;
    wire \c0.rx.r_Rx_Data_R ;
    wire n10010;
    wire rx_data_5;
    wire \c0.n24_adj_2317 ;
    wire \c0.n22_adj_2319 ;
    wire \c0.n21_adj_2323 ;
    wire \c0.FRAME_MATCHER_i_0 ;
    wire \c0.FRAME_MATCHER_i_2 ;
    wire \c0.n15171_cascade_ ;
    wire \c0.data_in_frame_1_6 ;
    wire \c0.n2124 ;
    wire data_in_frame_6_6;
    wire \c0.n17214 ;
    wire \c0.n28_adj_2374 ;
    wire \c0.n27_adj_2381_cascade_ ;
    wire \c0.n29 ;
    wire \c0.n12491_cascade_ ;
    wire \c0.data_in_frame_0_1 ;
    wire \c0.n10259 ;
    wire \c0.data_in_frame_2_7 ;
    wire rx_data_2;
    wire \c0.n15179 ;
    wire \c0.n17686 ;
    wire \c0.data_out_frame2_0_4 ;
    wire \c0.n17688 ;
    wire \c0.data_out_frame2_0_3 ;
    wire \c0.data_in_frame_3_7 ;
    wire \c0.n2126 ;
    wire \c0.data_in_frame_3_0 ;
    wire \c0.n2138 ;
    wire \c0.data_in_frame_2_1 ;
    wire \c0.data_in_frame_2_2 ;
    wire \c0.n18_adj_2316_cascade_ ;
    wire \c0.data_in_frame_0_7 ;
    wire \c0.n23_adj_2322 ;
    wire \c0.FRAME_MATCHER_state_23 ;
    wire \c0.n13381 ;
    wire \c0.FRAME_MATCHER_state_11 ;
    wire \c0.n8_adj_2333 ;
    wire data_out_frame2_8_2;
    wire \c0.n16 ;
    wire n4_adj_2427;
    wire n4_adj_2416;
    wire r_Bit_Index_1_adj_2436;
    wire r_Bit_Index_2_adj_2435;
    wire r_Bit_Index_0;
    wire \c0.rx.n10158 ;
    wire \c0.FRAME_MATCHER_state_16 ;
    wire \c0.n48 ;
    wire \c0.FRAME_MATCHER_state_30 ;
    wire \c0.n16698 ;
    wire \c0.FRAME_MATCHER_state_27 ;
    wire \c0.n16718 ;
    wire rand_setpoint_0;
    wire n2;
    wire data_out_2_0;
    wire rand_setpoint_7;
    wire data_out_0_0;
    wire rand_setpoint_16;
    wire rand_setpoint_15;
    wire n10_adj_2450;
    wire n10_adj_2411_cascade_;
    wire n5_adj_2407;
    wire \c0.n5_adj_2141 ;
    wire r_Tx_Data_2;
    wire r_Tx_Data_4;
    wire n18196_cascade_;
    wire n18199;
    wire \c0.tx.n31 ;
    wire n17759;
    wire n17664;
    wire \c0.n18166 ;
    wire \c0.n2_adj_2145 ;
    wire \c0.n17701 ;
    wire n18169;
    wire \c0.n453 ;
    wire n4_adj_2414;
    wire \c0.n19 ;
    wire n9524_cascade_;
    wire \c0.n16267_cascade_ ;
    wire \c0.n445 ;
    wire \c0.n23_adj_2314 ;
    wire \c0.n28 ;
    wire n17765;
    wire n17392_cascade_;
    wire n17416;
    wire \c0.n20_adj_2255 ;
    wire \c0.delay_counter_7 ;
    wire \c0.delay_counter_5 ;
    wire \c0.n24_adj_2389_cascade_ ;
    wire n17327;
    wire \c0.delay_counter_1 ;
    wire \c0.delay_counter_9 ;
    wire \c0.n26_adj_2391 ;
    wire \c0.delay_counter_4 ;
    wire \c0.n9453_cascade_ ;
    wire \c0.n24_adj_2342 ;
    wire \c0.delay_counter_12 ;
    wire \c0.n16_adj_2212 ;
    wire \c0.delay_counter_2 ;
    wire \c0.n26 ;
    wire \c0.delay_counter_0 ;
    wire \c0.delay_counter_6 ;
    wire \c0.n22_adj_2390 ;
    wire \c0.delay_counter_10 ;
    wire \c0.n18_adj_2220 ;
    wire \c0.delay_counter_13 ;
    wire \c0.n15_adj_2211 ;
    wire r_Tx_Data_5;
    wire \c0.delay_counter_11 ;
    wire \c0.n9453 ;
    wire \c0.n16267 ;
    wire \c0.n17_adj_2219 ;
    wire \c0.delay_counter_8 ;
    wire \c0.delay_counter_3 ;
    wire \c0.n18_adj_2388 ;
    wire \c0.n17712 ;
    wire \c0.n11867 ;
    wire \c0.byte_transmit_counter2_5 ;
    wire \c0.n4_adj_2147 ;
    wire n13116;
    wire rx_data_6;
    wire rx_data_1;
    wire \c0.n17072 ;
    wire \c0.data_in_frame_3_1 ;
    wire \c0.n17472_cascade_ ;
    wire \c0.data_out_frame2_0_6 ;
    wire rx_data_ready;
    wire data_in_3_2;
    wire data_in_2_2;
    wire \c0.data_in_frame_1_3 ;
    wire \c0.data_in_frame_5_4 ;
    wire \c0.data_in_frame_1_2 ;
    wire \c0.n21_adj_2357 ;
    wire \c0.data_out_frame2_0_0 ;
    wire \c0.n17490 ;
    wire \c0.n15171 ;
    wire rx_data_7;
    wire \c0.n17076 ;
    wire \c0.n26_adj_2174 ;
    wire \c0.n17487_cascade_ ;
    wire \c0.data_out_frame2_0_1 ;
    wire FRAME_MATCHER_state_0;
    wire \c0.n12491 ;
    wire \c0.n17690_cascade_ ;
    wire \c0.data_out_frame2_0_2 ;
    wire \c0.data_in_frame_5_2 ;
    wire \c0.data_in_frame_1_0 ;
    wire \c0.data_in_frame_1_1 ;
    wire \c0.n17102 ;
    wire \c0.n5815 ;
    wire \c0.n4494 ;
    wire \c0.n5817 ;
    wire n31_adj_2415;
    wire \c0.n18202 ;
    wire \c0.FRAME_MATCHER_state_29 ;
    wire \c0.n16658 ;
    wire \c0.FRAME_MATCHER_state_10 ;
    wire \c0.n16710 ;
    wire data_out_frame2_13_4;
    wire data_out_frame2_9_0;
    wire \c0.n17315 ;
    wire \c0.data_in_frame_0_0 ;
    wire \c0.data_in_frame_1_7 ;
    wire \c0.n17213 ;
    wire data_out_frame2_8_5;
    wire data_out_frame2_6_6;
    wire \c0.n10472 ;
    wire \c0.n15821 ;
    wire \c0.FRAME_MATCHER_state_18 ;
    wire \c0.n8_adj_2329 ;
    wire \c0.n8_adj_2385 ;
    wire \c0.n46 ;
    wire FRAME_MATCHER_i_31__N_1272;
    wire n488;
    wire \c0.n13146 ;
    wire n4408;
    wire \c0.n276_cascade_ ;
    wire \c0.n4_adj_2135 ;
    wire \c0.n4_adj_2135_cascade_ ;
    wire \c0.FRAME_MATCHER_state_31 ;
    wire \c0.n16700 ;
    wire \c0.n9334 ;
    wire n44;
    wire \c0.n17069 ;
    wire \c0.FRAME_MATCHER_state_17 ;
    wire \c0.n16704 ;
    wire \c0.n3_adj_2193 ;
    wire n10_adj_2431;
    wire \c0.n6_adj_2221 ;
    wire \c0.n17147 ;
    wire rand_setpoint_8;
    wire \c0.n17653 ;
    wire data_out_8_1;
    wire \c0.n1_adj_2160 ;
    wire \c0.n18184_cascade_ ;
    wire n18187_cascade_;
    wire \c0.data_out_6_6 ;
    wire \c0.n5_adj_2159 ;
    wire rand_setpoint_30;
    wire \c0.n17698 ;
    wire \c0.n17612 ;
    wire \c0.n17626 ;
    wire n25;
    wire n28;
    wire n5_adj_2448_cascade_;
    wire n31_cascade_;
    wire n22;
    wire n9524;
    wire n450;
    wire r_Bit_Index_1;
    wire \c0.tx.r_Bit_Index_0 ;
    wire r_Bit_Index_2;
    wire \c0.tx.n17673_cascade_ ;
    wire \c0.n10326 ;
    wire \c0.n17126 ;
    wire \c0.n17126_cascade_ ;
    wire \c0.n17651 ;
    wire n10705;
    wire n10_adj_2444;
    wire bfn_14_30_0_;
    wire \c0.n16110 ;
    wire \c0.n16111 ;
    wire \c0.n16112 ;
    wire \c0.n16113 ;
    wire byte_transmit_counter_5;
    wire \c0.n16114 ;
    wire byte_transmit_counter_6;
    wire \c0.n16115 ;
    wire byte_transmit_counter_7;
    wire \c0.n16116 ;
    wire \c0.n68_cascade_ ;
    wire tx_transmit_N_1947_7;
    wire \c0.n4650 ;
    wire tx_transmit_N_1947_3;
    wire \c0.n59 ;
    wire \c0.n65 ;
    wire tx_transmit_N_1947_4;
    wire tx_transmit_N_1947_5;
    wire tx_transmit_N_1947_6;
    wire \c0.n17404 ;
    wire tx_transmit_N_1947_1;
    wire tx_transmit_N_1947_0;
    wire \c0.n13662 ;
    wire \c0.n13662_cascade_ ;
    wire tx_transmit_N_1947_2;
    wire \c0.n13726 ;
    wire \c0.n10815 ;
    wire data_out_0_3;
    wire n10_adj_2483;
    wire \c0.data_out_3_6 ;
    wire \c0.FRAME_MATCHER_state_25 ;
    wire \c0.n16690 ;
    wire \c0.FRAME_MATCHER_state_26 ;
    wire \c0.n16702 ;
    wire \c0.FRAME_MATCHER_state_15 ;
    wire \c0.n8_adj_2330 ;
    wire \c0.FRAME_MATCHER_state_21 ;
    wire \c0.n16686 ;
    wire \c0.FRAME_MATCHER_state_24 ;
    wire \c0.n16688 ;
    wire \c0.n15_adj_2177 ;
    wire \c0.n17270 ;
    wire \c0.data_out_7_2 ;
    wire \c0.n10316 ;
    wire \c0.n17201 ;
    wire \c0.n10316_cascade_ ;
    wire \c0.n17177 ;
    wire data_out_8_6;
    wire \c0.data_out_6__1__N_537 ;
    wire \c0.data_out_7_7 ;
    wire rand_setpoint_5;
    wire n2594;
    wire rand_setpoint_13;
    wire \c0.data_out_7_5 ;
    wire r_Tx_Data_7;
    wire \c0.data_out_1_1 ;
    wire data_out_0_1;
    wire n1_adj_2449;
    wire \c0.n12630 ;
    wire \c0.data_out_7_0 ;
    wire \c0.n10395 ;
    wire \c0.n10_adj_2189_cascade_ ;
    wire r_Tx_Data_0;
    wire \c0.n8_adj_2157 ;
    wire n10_adj_2422;
    wire \c0.tx.n77_cascade_ ;
    wire \c0.tx.n12 ;
    wire tx_o;
    wire \c0.tx.n10 ;
    wire byte_transmit_counter_4;
    wire n10_adj_2443;
    wire r_Tx_Data_6;
    wire \c0.tx.n12_adj_2134 ;
    wire \c0.n8_cascade_ ;
    wire n9257;
    wire \c0.n65_adj_2192 ;
    wire \c0.tx.r_SM_Main_0 ;
    wire \c0.tx.n83 ;
    wire n5142_cascade_;
    wire \c0.tx.n6759 ;
    wire \c0.tx.n13702 ;
    wire \c0.tx_active_prev ;
    wire \c0.data_out_5_5 ;
    wire \c0.n5_adj_2163 ;
    wire \c0.n17581_cascade_ ;
    wire n10_adj_2432;
    wire \c0.tx.r_SM_Main_1 ;
    wire \c0.tx.n10613 ;
    wire \c0.n17622 ;
    wire \c0.n18088 ;
    wire \c0.n2_adj_2164_cascade_ ;
    wire n18091;
    wire data_out_3_5;
    wire \c0.data_out_0_6 ;
    wire n4;
    wire r_Rx_Data;
    wire n9999;
    wire rx_data_4;
    wire data_out_1_6;
    wire \c0.n9369 ;
    wire \c0.n276 ;
    wire FRAME_MATCHER_i_31__N_1275;
    wire \c0.FRAME_MATCHER_state_22 ;
    wire \c0.n16714 ;
    wire data_out_1_7;
    wire \c0.n8_adj_2352 ;
    wire \c0.n10179 ;
    wire \c0.n10188 ;
    wire \c0.n17209_cascade_ ;
    wire \c0.data_out_10_2 ;
    wire \c0.n6_adj_2216 ;
    wire \c0.data_out_9_6 ;
    wire \c0.n17200 ;
    wire \c0.data_out_8_0 ;
    wire n8_adj_2445;
    wire n6_adj_2446;
    wire n23;
    wire n32;
    wire n29_cascade_;
    wire n26;
    wire \c0.data_out_5_2 ;
    wire \c0.n10196 ;
    wire \c0.n10196_cascade_ ;
    wire \c0.data_out_10_3 ;
    wire \c0.data_out_6_4 ;
    wire data_out_8_5;
    wire \c0.n10392 ;
    wire bfn_16_28_0_;
    wire \c0.tx.n16117 ;
    wire \c0.tx.r_Clock_Count_2 ;
    wire n10954;
    wire \c0.tx.n16118 ;
    wire \c0.tx.r_Clock_Count_3 ;
    wire n10957;
    wire \c0.tx.n16119 ;
    wire \c0.tx.n16120 ;
    wire \c0.tx.r_Clock_Count_5 ;
    wire n10963;
    wire \c0.tx.n16121 ;
    wire \c0.tx.r_Clock_Count_6 ;
    wire n10966;
    wire \c0.tx.n16122 ;
    wire \c0.tx.n16123 ;
    wire \c0.tx.n16124 ;
    wire \c0.tx.r_Clock_Count_8 ;
    wire \c0.tx.r_SM_Main_2 ;
    wire bfn_16_29_0_;
    wire n10972;
    wire data_out_8_7;
    wire n10951;
    wire \c0.tx.r_Clock_Count_1 ;
    wire n10969;
    wire \c0.tx.r_Clock_Count_7 ;
    wire data_out_3_7;
    wire data_out_2_7;
    wire \c0.data_out_7__3__N_441 ;
    wire \c0.n1 ;
    wire \c0.n17747_cascade_ ;
    wire \c0.n2_adj_2156 ;
    wire \c0.n18220_cascade_ ;
    wire \c0.n17607 ;
    wire byte_transmit_counter_3;
    wire n10_adj_2413;
    wire n18223_cascade_;
    wire byte_transmit_counter_2;
    wire n10;
    wire n10960;
    wire \c0.tx.r_Clock_Count_4 ;
    wire n10994;
    wire n5142;
    wire \c0.tx.r_Clock_Count_0 ;
    wire \c0.n10595 ;
    wire \c0.data_out_6_0 ;
    wire \c0.n17129 ;
    wire \c0.n10447_cascade_ ;
    wire \c0.data_out_6_1 ;
    wire \c0.n10183 ;
    wire \c0.data_out_6_3 ;
    wire \c0.n17222 ;
    wire \c0.data_out_9_7 ;
    wire \c0.n17243 ;
    wire \c0.n17264 ;
    wire \c0.n10_adj_2191_cascade_ ;
    wire byte_transmit_counter_0;
    wire \c0.data_out_10_4 ;
    wire \c0.n8_adj_2198_cascade_ ;
    wire byte_transmit_counter_1;
    wire n10_adj_2430;
    wire \c0.n17209 ;
    wire \c0.n17297 ;
    wire \c0.n17297_cascade_ ;
    wire \c0.data_out_7__2__N_447 ;
    wire \c0.n14_adj_2176 ;
    wire \c0.data_out_7_6 ;
    wire \c0.n12_adj_2180 ;
    wire data_out_10_0;
    wire \c0.data_out_7_3 ;
    wire \c0.data_out_5_3 ;
    wire \c0.n17180 ;
    wire \c0.data_out_9_4 ;
    wire \c0.n17162_cascade_ ;
    wire \c0.data_out_6_2 ;
    wire \c0.n17197 ;
    wire \c0.n10_adj_2196_cascade_ ;
    wire \c0.n17261 ;
    wire \c0.data_out_6_7 ;
    wire \c0.n26_adj_2165 ;
    wire \c0.data_out_6_5 ;
    wire data_out_8_3;
    wire \c0.n10_adj_2166_cascade_ ;
    wire \c0.n10170 ;
    wire \c0.n17252 ;
    wire data_out_10_1;
    wire data_out_8_2;
    wire \c0.data_out_10_5 ;
    wire \c0.data_out_7_1 ;
    wire \c0.data_out_9_0 ;
    wire \c0.n6_adj_2169 ;
    wire \c0.n17162 ;
    wire \c0.n17150_cascade_ ;
    wire \c0.data_out_9_1 ;
    wire \c0.data_out_9_5 ;
    wire \c0.n17110 ;
    wire data_out_8_4;
    wire \c0.data_out_10_7 ;
    wire UART_TRANSMITTER_state_2;
    wire UART_TRANSMITTER_state_0;
    wire rand_setpoint_25;
    wire data_out_5_1;
    wire \c0.r_SM_Main_2_N_2034_0 ;
    wire \c0.tx_active ;
    wire n444;
    wire n10596;
    wire UART_TRANSMITTER_state_1;
    wire data_out_2_5;
    wire data_out_10__7__N_110;
    wire data_out_9__2__N_367;
    wire CLK_c;
    wire data_out_9_2;
    wire \c0.data_out_5_4 ;
    wire \c0.data_out_10_6 ;
    wire \c0.data_out_9_3 ;
    wire \c0.n10204_cascade_ ;
    wire \c0.data_out_7_4 ;
    wire \c0.n10_adj_2172 ;
    wire _gnd_net_;

    defparam LED_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam LED_pad_iopad.PULLUP=1'b0;
    IO_PAD LED_pad_iopad (
            .OE(N__50887),
            .DIN(N__50886),
            .DOUT(N__50885),
            .PACKAGEPIN(LED));
    defparam LED_pad_preio.PIN_TYPE=6'b011001;
    defparam LED_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO LED_pad_preio (
            .PADOEN(N__50887),
            .PADOUT(N__50886),
            .PADIN(N__50885),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__35976),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam USBPU_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam USBPU_pad_iopad.PULLUP=1'b0;
    IO_PAD USBPU_pad_iopad (
            .OE(N__50878),
            .DIN(N__50877),
            .DOUT(N__50876),
            .PACKAGEPIN(USBPU));
    defparam USBPU_pad_preio.PIN_TYPE=6'b011001;
    defparam USBPU_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO USBPU_pad_preio (
            .PADOEN(N__50878),
            .PADOUT(N__50877),
            .PADIN(N__50876),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam rx_input_iopad.IO_STANDARD="SB_LVCMOS";
    defparam rx_input_iopad.PULLUP=1'b1;
    IO_PAD rx_input_iopad (
            .OE(N__50869),
            .DIN(N__50868),
            .DOUT(N__50867),
            .PACKAGEPIN(PIN_2));
    defparam rx_input_preio.PIN_TYPE=6'b000000;
    defparam rx_input_preio.NEG_TRIGGER=1'b0;
    PRE_IO rx_input_preio (
            .PADOEN(N__50869),
            .PADOUT(N__50868),
            .PADIN(N__50867),
            .CLOCKENABLE(VCCG0),
            .DIN0(\c0.rx.r_Rx_Data_R ),
            .DIN1(),
            .DOUT0(GNDG0),
            .DOUT1(GNDG0),
            .INPUTCLK(N__49762),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    defparam tx2_output_iopad.IO_STANDARD="SB_LVCMOS";
    defparam tx2_output_iopad.PULLUP=1'b1;
    IO_PAD tx2_output_iopad (
            .OE(N__50860),
            .DIN(N__50859),
            .DOUT(N__50858),
            .PACKAGEPIN(PIN_3));
    defparam tx2_output_preio.PIN_TYPE=6'b101001;
    defparam tx2_output_preio.NEG_TRIGGER=1'b0;
    PRE_IO tx2_output_preio (
            .PADOEN(N__50860),
            .PADOUT(N__50859),
            .PADIN(N__50858),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__22131),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__17694));
    defparam tx_output_iopad.IO_STANDARD="SB_LVCMOS";
    defparam tx_output_iopad.PULLUP=1'b1;
    IO_PAD tx_output_iopad (
            .OE(N__50851),
            .DIN(N__50850),
            .DOUT(N__50849),
            .PACKAGEPIN(PIN_1));
    defparam tx_output_preio.PIN_TYPE=6'b101001;
    defparam tx_output_preio.NEG_TRIGGER=1'b0;
    PRE_IO tx_output_preio (
            .PADOEN(N__50851),
            .PADOUT(N__50850),
            .PADIN(N__50849),
            .CLOCKENABLE(),
            .DIN0(),
            .DIN1(),
            .DOUT0(N__43887),
            .DOUT1(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(N__25689));
    defparam CLK_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam CLK_pad_iopad.PULLUP=1'b0;
    IO_PAD CLK_pad_iopad (
            .OE(N__50842),
            .DIN(N__50841),
            .DOUT(N__50840),
            .PACKAGEPIN(CLK));
    defparam CLK_pad_preio.PIN_TYPE=6'b000001;
    defparam CLK_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO CLK_pad_preio (
            .PADOEN(N__50842),
            .PADOUT(N__50841),
            .PADIN(N__50840),
            .CLOCKENABLE(),
            .DIN0(CLK_pad_gb_input),
            .DIN1(),
            .DOUT0(),
            .DOUT1(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .OUTPUTCLK(),
            .OUTPUTENABLE());
    InMux I__12827 (
            .O(N__50823),
            .I(N__50820));
    LocalMux I__12826 (
            .O(N__50820),
            .I(N__50813));
    InMux I__12825 (
            .O(N__50819),
            .I(N__50808));
    InMux I__12824 (
            .O(N__50818),
            .I(N__50808));
    InMux I__12823 (
            .O(N__50817),
            .I(N__50805));
    InMux I__12822 (
            .O(N__50816),
            .I(N__50802));
    Span4Mux_v I__12821 (
            .O(N__50813),
            .I(N__50799));
    LocalMux I__12820 (
            .O(N__50808),
            .I(N__50796));
    LocalMux I__12819 (
            .O(N__50805),
            .I(N__50793));
    LocalMux I__12818 (
            .O(N__50802),
            .I(N__50790));
    Odrv4 I__12817 (
            .O(N__50799),
            .I(\c0.r_SM_Main_2_N_2034_0 ));
    Odrv4 I__12816 (
            .O(N__50796),
            .I(\c0.r_SM_Main_2_N_2034_0 ));
    Odrv4 I__12815 (
            .O(N__50793),
            .I(\c0.r_SM_Main_2_N_2034_0 ));
    Odrv4 I__12814 (
            .O(N__50790),
            .I(\c0.r_SM_Main_2_N_2034_0 ));
    CascadeMux I__12813 (
            .O(N__50781),
            .I(N__50777));
    InMux I__12812 (
            .O(N__50780),
            .I(N__50774));
    InMux I__12811 (
            .O(N__50777),
            .I(N__50770));
    LocalMux I__12810 (
            .O(N__50774),
            .I(N__50767));
    InMux I__12809 (
            .O(N__50773),
            .I(N__50764));
    LocalMux I__12808 (
            .O(N__50770),
            .I(N__50755));
    Span4Mux_v I__12807 (
            .O(N__50767),
            .I(N__50755));
    LocalMux I__12806 (
            .O(N__50764),
            .I(N__50755));
    InMux I__12805 (
            .O(N__50763),
            .I(N__50750));
    InMux I__12804 (
            .O(N__50762),
            .I(N__50750));
    Odrv4 I__12803 (
            .O(N__50755),
            .I(\c0.tx_active ));
    LocalMux I__12802 (
            .O(N__50750),
            .I(\c0.tx_active ));
    CascadeMux I__12801 (
            .O(N__50745),
            .I(N__50737));
    CascadeMux I__12800 (
            .O(N__50744),
            .I(N__50734));
    CascadeMux I__12799 (
            .O(N__50743),
            .I(N__50730));
    CascadeMux I__12798 (
            .O(N__50742),
            .I(N__50727));
    CascadeMux I__12797 (
            .O(N__50741),
            .I(N__50724));
    InMux I__12796 (
            .O(N__50740),
            .I(N__50710));
    InMux I__12795 (
            .O(N__50737),
            .I(N__50710));
    InMux I__12794 (
            .O(N__50734),
            .I(N__50710));
    InMux I__12793 (
            .O(N__50733),
            .I(N__50707));
    InMux I__12792 (
            .O(N__50730),
            .I(N__50700));
    InMux I__12791 (
            .O(N__50727),
            .I(N__50700));
    InMux I__12790 (
            .O(N__50724),
            .I(N__50700));
    CascadeMux I__12789 (
            .O(N__50723),
            .I(N__50695));
    CascadeMux I__12788 (
            .O(N__50722),
            .I(N__50692));
    CascadeMux I__12787 (
            .O(N__50721),
            .I(N__50689));
    CascadeMux I__12786 (
            .O(N__50720),
            .I(N__50685));
    InMux I__12785 (
            .O(N__50719),
            .I(N__50681));
    InMux I__12784 (
            .O(N__50718),
            .I(N__50678));
    CascadeMux I__12783 (
            .O(N__50717),
            .I(N__50673));
    LocalMux I__12782 (
            .O(N__50710),
            .I(N__50670));
    LocalMux I__12781 (
            .O(N__50707),
            .I(N__50667));
    LocalMux I__12780 (
            .O(N__50700),
            .I(N__50664));
    InMux I__12779 (
            .O(N__50699),
            .I(N__50657));
    InMux I__12778 (
            .O(N__50698),
            .I(N__50657));
    InMux I__12777 (
            .O(N__50695),
            .I(N__50657));
    InMux I__12776 (
            .O(N__50692),
            .I(N__50654));
    InMux I__12775 (
            .O(N__50689),
            .I(N__50649));
    InMux I__12774 (
            .O(N__50688),
            .I(N__50649));
    InMux I__12773 (
            .O(N__50685),
            .I(N__50646));
    InMux I__12772 (
            .O(N__50684),
            .I(N__50643));
    LocalMux I__12771 (
            .O(N__50681),
            .I(N__50638));
    LocalMux I__12770 (
            .O(N__50678),
            .I(N__50638));
    InMux I__12769 (
            .O(N__50677),
            .I(N__50631));
    InMux I__12768 (
            .O(N__50676),
            .I(N__50631));
    InMux I__12767 (
            .O(N__50673),
            .I(N__50631));
    Span4Mux_s2_v I__12766 (
            .O(N__50670),
            .I(N__50622));
    Span4Mux_v I__12765 (
            .O(N__50667),
            .I(N__50622));
    Span4Mux_h I__12764 (
            .O(N__50664),
            .I(N__50622));
    LocalMux I__12763 (
            .O(N__50657),
            .I(N__50622));
    LocalMux I__12762 (
            .O(N__50654),
            .I(N__50617));
    LocalMux I__12761 (
            .O(N__50649),
            .I(N__50617));
    LocalMux I__12760 (
            .O(N__50646),
            .I(N__50612));
    LocalMux I__12759 (
            .O(N__50643),
            .I(N__50612));
    Span4Mux_v I__12758 (
            .O(N__50638),
            .I(N__50607));
    LocalMux I__12757 (
            .O(N__50631),
            .I(N__50607));
    Span4Mux_h I__12756 (
            .O(N__50622),
            .I(N__50604));
    Span12Mux_h I__12755 (
            .O(N__50617),
            .I(N__50601));
    Span4Mux_h I__12754 (
            .O(N__50612),
            .I(N__50596));
    Span4Mux_h I__12753 (
            .O(N__50607),
            .I(N__50596));
    Odrv4 I__12752 (
            .O(N__50604),
            .I(n444));
    Odrv12 I__12751 (
            .O(N__50601),
            .I(n444));
    Odrv4 I__12750 (
            .O(N__50596),
            .I(n444));
    CEMux I__12749 (
            .O(N__50589),
            .I(N__50584));
    CEMux I__12748 (
            .O(N__50588),
            .I(N__50580));
    CascadeMux I__12747 (
            .O(N__50587),
            .I(N__50577));
    LocalMux I__12746 (
            .O(N__50584),
            .I(N__50571));
    CascadeMux I__12745 (
            .O(N__50583),
            .I(N__50568));
    LocalMux I__12744 (
            .O(N__50580),
            .I(N__50563));
    InMux I__12743 (
            .O(N__50577),
            .I(N__50560));
    CascadeMux I__12742 (
            .O(N__50576),
            .I(N__50557));
    CEMux I__12741 (
            .O(N__50575),
            .I(N__50549));
    CascadeMux I__12740 (
            .O(N__50574),
            .I(N__50543));
    Span4Mux_s3_h I__12739 (
            .O(N__50571),
            .I(N__50538));
    InMux I__12738 (
            .O(N__50568),
            .I(N__50534));
    CEMux I__12737 (
            .O(N__50567),
            .I(N__50530));
    CEMux I__12736 (
            .O(N__50566),
            .I(N__50526));
    Span4Mux_v I__12735 (
            .O(N__50563),
            .I(N__50521));
    LocalMux I__12734 (
            .O(N__50560),
            .I(N__50521));
    InMux I__12733 (
            .O(N__50557),
            .I(N__50518));
    InMux I__12732 (
            .O(N__50556),
            .I(N__50511));
    InMux I__12731 (
            .O(N__50555),
            .I(N__50511));
    InMux I__12730 (
            .O(N__50554),
            .I(N__50511));
    InMux I__12729 (
            .O(N__50553),
            .I(N__50506));
    InMux I__12728 (
            .O(N__50552),
            .I(N__50506));
    LocalMux I__12727 (
            .O(N__50549),
            .I(N__50502));
    CEMux I__12726 (
            .O(N__50548),
            .I(N__50499));
    CascadeMux I__12725 (
            .O(N__50547),
            .I(N__50496));
    CascadeMux I__12724 (
            .O(N__50546),
            .I(N__50493));
    InMux I__12723 (
            .O(N__50543),
            .I(N__50484));
    InMux I__12722 (
            .O(N__50542),
            .I(N__50484));
    InMux I__12721 (
            .O(N__50541),
            .I(N__50484));
    Span4Mux_h I__12720 (
            .O(N__50538),
            .I(N__50481));
    InMux I__12719 (
            .O(N__50537),
            .I(N__50478));
    LocalMux I__12718 (
            .O(N__50534),
            .I(N__50475));
    InMux I__12717 (
            .O(N__50533),
            .I(N__50472));
    LocalMux I__12716 (
            .O(N__50530),
            .I(N__50467));
    CascadeMux I__12715 (
            .O(N__50529),
            .I(N__50464));
    LocalMux I__12714 (
            .O(N__50526),
            .I(N__50457));
    Span4Mux_h I__12713 (
            .O(N__50521),
            .I(N__50457));
    LocalMux I__12712 (
            .O(N__50518),
            .I(N__50457));
    LocalMux I__12711 (
            .O(N__50511),
            .I(N__50452));
    LocalMux I__12710 (
            .O(N__50506),
            .I(N__50452));
    InMux I__12709 (
            .O(N__50505),
            .I(N__50449));
    Span4Mux_v I__12708 (
            .O(N__50502),
            .I(N__50446));
    LocalMux I__12707 (
            .O(N__50499),
            .I(N__50443));
    InMux I__12706 (
            .O(N__50496),
            .I(N__50436));
    InMux I__12705 (
            .O(N__50493),
            .I(N__50436));
    InMux I__12704 (
            .O(N__50492),
            .I(N__50436));
    CEMux I__12703 (
            .O(N__50491),
            .I(N__50433));
    LocalMux I__12702 (
            .O(N__50484),
            .I(N__50430));
    Span4Mux_h I__12701 (
            .O(N__50481),
            .I(N__50427));
    LocalMux I__12700 (
            .O(N__50478),
            .I(N__50424));
    Span4Mux_v I__12699 (
            .O(N__50475),
            .I(N__50419));
    LocalMux I__12698 (
            .O(N__50472),
            .I(N__50419));
    CascadeMux I__12697 (
            .O(N__50471),
            .I(N__50415));
    CascadeMux I__12696 (
            .O(N__50470),
            .I(N__50412));
    Span4Mux_v I__12695 (
            .O(N__50467),
            .I(N__50408));
    InMux I__12694 (
            .O(N__50464),
            .I(N__50405));
    Span4Mux_v I__12693 (
            .O(N__50457),
            .I(N__50398));
    Span4Mux_s1_v I__12692 (
            .O(N__50452),
            .I(N__50398));
    LocalMux I__12691 (
            .O(N__50449),
            .I(N__50398));
    Span4Mux_h I__12690 (
            .O(N__50446),
            .I(N__50391));
    Span4Mux_v I__12689 (
            .O(N__50443),
            .I(N__50391));
    LocalMux I__12688 (
            .O(N__50436),
            .I(N__50391));
    LocalMux I__12687 (
            .O(N__50433),
            .I(N__50387));
    Span12Mux_v I__12686 (
            .O(N__50430),
            .I(N__50384));
    Span4Mux_h I__12685 (
            .O(N__50427),
            .I(N__50377));
    Span4Mux_v I__12684 (
            .O(N__50424),
            .I(N__50377));
    Span4Mux_v I__12683 (
            .O(N__50419),
            .I(N__50377));
    InMux I__12682 (
            .O(N__50418),
            .I(N__50372));
    InMux I__12681 (
            .O(N__50415),
            .I(N__50372));
    InMux I__12680 (
            .O(N__50412),
            .I(N__50369));
    InMux I__12679 (
            .O(N__50411),
            .I(N__50366));
    Span4Mux_v I__12678 (
            .O(N__50408),
            .I(N__50357));
    LocalMux I__12677 (
            .O(N__50405),
            .I(N__50357));
    Span4Mux_h I__12676 (
            .O(N__50398),
            .I(N__50357));
    Span4Mux_s1_v I__12675 (
            .O(N__50391),
            .I(N__50357));
    InMux I__12674 (
            .O(N__50390),
            .I(N__50354));
    Odrv4 I__12673 (
            .O(N__50387),
            .I(n10596));
    Odrv12 I__12672 (
            .O(N__50384),
            .I(n10596));
    Odrv4 I__12671 (
            .O(N__50377),
            .I(n10596));
    LocalMux I__12670 (
            .O(N__50372),
            .I(n10596));
    LocalMux I__12669 (
            .O(N__50369),
            .I(n10596));
    LocalMux I__12668 (
            .O(N__50366),
            .I(n10596));
    Odrv4 I__12667 (
            .O(N__50357),
            .I(n10596));
    LocalMux I__12666 (
            .O(N__50354),
            .I(n10596));
    InMux I__12665 (
            .O(N__50337),
            .I(N__50334));
    LocalMux I__12664 (
            .O(N__50334),
            .I(N__50330));
    CascadeMux I__12663 (
            .O(N__50333),
            .I(N__50325));
    Span4Mux_h I__12662 (
            .O(N__50330),
            .I(N__50311));
    InMux I__12661 (
            .O(N__50329),
            .I(N__50306));
    InMux I__12660 (
            .O(N__50328),
            .I(N__50306));
    InMux I__12659 (
            .O(N__50325),
            .I(N__50301));
    InMux I__12658 (
            .O(N__50324),
            .I(N__50301));
    InMux I__12657 (
            .O(N__50323),
            .I(N__50296));
    InMux I__12656 (
            .O(N__50322),
            .I(N__50296));
    CascadeMux I__12655 (
            .O(N__50321),
            .I(N__50293));
    InMux I__12654 (
            .O(N__50320),
            .I(N__50287));
    InMux I__12653 (
            .O(N__50319),
            .I(N__50284));
    InMux I__12652 (
            .O(N__50318),
            .I(N__50281));
    InMux I__12651 (
            .O(N__50317),
            .I(N__50278));
    InMux I__12650 (
            .O(N__50316),
            .I(N__50272));
    InMux I__12649 (
            .O(N__50315),
            .I(N__50267));
    CascadeMux I__12648 (
            .O(N__50314),
            .I(N__50263));
    Span4Mux_h I__12647 (
            .O(N__50311),
            .I(N__50254));
    LocalMux I__12646 (
            .O(N__50306),
            .I(N__50254));
    LocalMux I__12645 (
            .O(N__50301),
            .I(N__50249));
    LocalMux I__12644 (
            .O(N__50296),
            .I(N__50249));
    InMux I__12643 (
            .O(N__50293),
            .I(N__50245));
    InMux I__12642 (
            .O(N__50292),
            .I(N__50241));
    InMux I__12641 (
            .O(N__50291),
            .I(N__50238));
    InMux I__12640 (
            .O(N__50290),
            .I(N__50233));
    LocalMux I__12639 (
            .O(N__50287),
            .I(N__50230));
    LocalMux I__12638 (
            .O(N__50284),
            .I(N__50227));
    LocalMux I__12637 (
            .O(N__50281),
            .I(N__50222));
    LocalMux I__12636 (
            .O(N__50278),
            .I(N__50222));
    InMux I__12635 (
            .O(N__50277),
            .I(N__50215));
    InMux I__12634 (
            .O(N__50276),
            .I(N__50215));
    InMux I__12633 (
            .O(N__50275),
            .I(N__50215));
    LocalMux I__12632 (
            .O(N__50272),
            .I(N__50212));
    InMux I__12631 (
            .O(N__50271),
            .I(N__50207));
    InMux I__12630 (
            .O(N__50270),
            .I(N__50207));
    LocalMux I__12629 (
            .O(N__50267),
            .I(N__50201));
    InMux I__12628 (
            .O(N__50266),
            .I(N__50198));
    InMux I__12627 (
            .O(N__50263),
            .I(N__50195));
    InMux I__12626 (
            .O(N__50262),
            .I(N__50192));
    InMux I__12625 (
            .O(N__50261),
            .I(N__50187));
    InMux I__12624 (
            .O(N__50260),
            .I(N__50187));
    InMux I__12623 (
            .O(N__50259),
            .I(N__50184));
    Span4Mux_h I__12622 (
            .O(N__50254),
            .I(N__50179));
    Span4Mux_h I__12621 (
            .O(N__50249),
            .I(N__50179));
    InMux I__12620 (
            .O(N__50248),
            .I(N__50176));
    LocalMux I__12619 (
            .O(N__50245),
            .I(N__50173));
    InMux I__12618 (
            .O(N__50244),
            .I(N__50170));
    LocalMux I__12617 (
            .O(N__50241),
            .I(N__50165));
    LocalMux I__12616 (
            .O(N__50238),
            .I(N__50165));
    InMux I__12615 (
            .O(N__50237),
            .I(N__50162));
    InMux I__12614 (
            .O(N__50236),
            .I(N__50159));
    LocalMux I__12613 (
            .O(N__50233),
            .I(N__50147));
    Span4Mux_h I__12612 (
            .O(N__50230),
            .I(N__50138));
    Span4Mux_s1_v I__12611 (
            .O(N__50227),
            .I(N__50138));
    Span4Mux_h I__12610 (
            .O(N__50222),
            .I(N__50138));
    LocalMux I__12609 (
            .O(N__50215),
            .I(N__50138));
    Span4Mux_s3_v I__12608 (
            .O(N__50212),
            .I(N__50130));
    LocalMux I__12607 (
            .O(N__50207),
            .I(N__50130));
    InMux I__12606 (
            .O(N__50206),
            .I(N__50125));
    InMux I__12605 (
            .O(N__50205),
            .I(N__50125));
    InMux I__12604 (
            .O(N__50204),
            .I(N__50122));
    Span4Mux_v I__12603 (
            .O(N__50201),
            .I(N__50119));
    LocalMux I__12602 (
            .O(N__50198),
            .I(N__50116));
    LocalMux I__12601 (
            .O(N__50195),
            .I(N__50111));
    LocalMux I__12600 (
            .O(N__50192),
            .I(N__50111));
    LocalMux I__12599 (
            .O(N__50187),
            .I(N__50108));
    LocalMux I__12598 (
            .O(N__50184),
            .I(N__50105));
    IoSpan4Mux I__12597 (
            .O(N__50179),
            .I(N__50100));
    LocalMux I__12596 (
            .O(N__50176),
            .I(N__50100));
    Span4Mux_v I__12595 (
            .O(N__50173),
            .I(N__50097));
    LocalMux I__12594 (
            .O(N__50170),
            .I(N__50088));
    Span12Mux_v I__12593 (
            .O(N__50165),
            .I(N__50088));
    LocalMux I__12592 (
            .O(N__50162),
            .I(N__50088));
    LocalMux I__12591 (
            .O(N__50159),
            .I(N__50088));
    InMux I__12590 (
            .O(N__50158),
            .I(N__50081));
    InMux I__12589 (
            .O(N__50157),
            .I(N__50081));
    InMux I__12588 (
            .O(N__50156),
            .I(N__50081));
    InMux I__12587 (
            .O(N__50155),
            .I(N__50076));
    InMux I__12586 (
            .O(N__50154),
            .I(N__50076));
    InMux I__12585 (
            .O(N__50153),
            .I(N__50073));
    InMux I__12584 (
            .O(N__50152),
            .I(N__50066));
    InMux I__12583 (
            .O(N__50151),
            .I(N__50066));
    InMux I__12582 (
            .O(N__50150),
            .I(N__50066));
    Span4Mux_v I__12581 (
            .O(N__50147),
            .I(N__50061));
    Span4Mux_v I__12580 (
            .O(N__50138),
            .I(N__50061));
    InMux I__12579 (
            .O(N__50137),
            .I(N__50054));
    InMux I__12578 (
            .O(N__50136),
            .I(N__50054));
    InMux I__12577 (
            .O(N__50135),
            .I(N__50054));
    Span4Mux_h I__12576 (
            .O(N__50130),
            .I(N__50047));
    LocalMux I__12575 (
            .O(N__50125),
            .I(N__50047));
    LocalMux I__12574 (
            .O(N__50122),
            .I(N__50047));
    Span4Mux_h I__12573 (
            .O(N__50119),
            .I(N__50044));
    Span4Mux_h I__12572 (
            .O(N__50116),
            .I(N__50033));
    Span4Mux_h I__12571 (
            .O(N__50111),
            .I(N__50033));
    Span4Mux_h I__12570 (
            .O(N__50108),
            .I(N__50033));
    Span4Mux_h I__12569 (
            .O(N__50105),
            .I(N__50033));
    Span4Mux_s2_v I__12568 (
            .O(N__50100),
            .I(N__50033));
    Sp12to4 I__12567 (
            .O(N__50097),
            .I(N__50028));
    Span12Mux_s5_v I__12566 (
            .O(N__50088),
            .I(N__50028));
    LocalMux I__12565 (
            .O(N__50081),
            .I(UART_TRANSMITTER_state_1));
    LocalMux I__12564 (
            .O(N__50076),
            .I(UART_TRANSMITTER_state_1));
    LocalMux I__12563 (
            .O(N__50073),
            .I(UART_TRANSMITTER_state_1));
    LocalMux I__12562 (
            .O(N__50066),
            .I(UART_TRANSMITTER_state_1));
    Odrv4 I__12561 (
            .O(N__50061),
            .I(UART_TRANSMITTER_state_1));
    LocalMux I__12560 (
            .O(N__50054),
            .I(UART_TRANSMITTER_state_1));
    Odrv4 I__12559 (
            .O(N__50047),
            .I(UART_TRANSMITTER_state_1));
    Odrv4 I__12558 (
            .O(N__50044),
            .I(UART_TRANSMITTER_state_1));
    Odrv4 I__12557 (
            .O(N__50033),
            .I(UART_TRANSMITTER_state_1));
    Odrv12 I__12556 (
            .O(N__50028),
            .I(UART_TRANSMITTER_state_1));
    InMux I__12555 (
            .O(N__50007),
            .I(N__50004));
    LocalMux I__12554 (
            .O(N__50004),
            .I(N__50000));
    InMux I__12553 (
            .O(N__50003),
            .I(N__49997));
    Span4Mux_s1_v I__12552 (
            .O(N__50000),
            .I(N__49994));
    LocalMux I__12551 (
            .O(N__49997),
            .I(data_out_2_5));
    Odrv4 I__12550 (
            .O(N__49994),
            .I(data_out_2_5));
    CEMux I__12549 (
            .O(N__49989),
            .I(N__49985));
    CEMux I__12548 (
            .O(N__49988),
            .I(N__49981));
    LocalMux I__12547 (
            .O(N__49985),
            .I(N__49974));
    CEMux I__12546 (
            .O(N__49984),
            .I(N__49971));
    LocalMux I__12545 (
            .O(N__49981),
            .I(N__49967));
    CEMux I__12544 (
            .O(N__49980),
            .I(N__49964));
    CEMux I__12543 (
            .O(N__49979),
            .I(N__49959));
    InMux I__12542 (
            .O(N__49978),
            .I(N__49956));
    InMux I__12541 (
            .O(N__49977),
            .I(N__49953));
    Span4Mux_v I__12540 (
            .O(N__49974),
            .I(N__49950));
    LocalMux I__12539 (
            .O(N__49971),
            .I(N__49947));
    CEMux I__12538 (
            .O(N__49970),
            .I(N__49944));
    Span4Mux_v I__12537 (
            .O(N__49967),
            .I(N__49939));
    LocalMux I__12536 (
            .O(N__49964),
            .I(N__49939));
    CascadeMux I__12535 (
            .O(N__49963),
            .I(N__49936));
    CascadeMux I__12534 (
            .O(N__49962),
            .I(N__49931));
    LocalMux I__12533 (
            .O(N__49959),
            .I(N__49924));
    LocalMux I__12532 (
            .O(N__49956),
            .I(N__49924));
    LocalMux I__12531 (
            .O(N__49953),
            .I(N__49921));
    Span4Mux_h I__12530 (
            .O(N__49950),
            .I(N__49916));
    Span4Mux_h I__12529 (
            .O(N__49947),
            .I(N__49916));
    LocalMux I__12528 (
            .O(N__49944),
            .I(N__49913));
    Span4Mux_h I__12527 (
            .O(N__49939),
            .I(N__49910));
    InMux I__12526 (
            .O(N__49936),
            .I(N__49907));
    InMux I__12525 (
            .O(N__49935),
            .I(N__49902));
    InMux I__12524 (
            .O(N__49934),
            .I(N__49902));
    InMux I__12523 (
            .O(N__49931),
            .I(N__49897));
    InMux I__12522 (
            .O(N__49930),
            .I(N__49897));
    InMux I__12521 (
            .O(N__49929),
            .I(N__49894));
    Span4Mux_h I__12520 (
            .O(N__49924),
            .I(N__49889));
    Span4Mux_v I__12519 (
            .O(N__49921),
            .I(N__49889));
    Span4Mux_h I__12518 (
            .O(N__49916),
            .I(N__49886));
    Span4Mux_h I__12517 (
            .O(N__49913),
            .I(N__49881));
    Span4Mux_h I__12516 (
            .O(N__49910),
            .I(N__49881));
    LocalMux I__12515 (
            .O(N__49907),
            .I(data_out_10__7__N_110));
    LocalMux I__12514 (
            .O(N__49902),
            .I(data_out_10__7__N_110));
    LocalMux I__12513 (
            .O(N__49897),
            .I(data_out_10__7__N_110));
    LocalMux I__12512 (
            .O(N__49894),
            .I(data_out_10__7__N_110));
    Odrv4 I__12511 (
            .O(N__49889),
            .I(data_out_10__7__N_110));
    Odrv4 I__12510 (
            .O(N__49886),
            .I(data_out_10__7__N_110));
    Odrv4 I__12509 (
            .O(N__49881),
            .I(data_out_10__7__N_110));
    InMux I__12508 (
            .O(N__49866),
            .I(N__49862));
    InMux I__12507 (
            .O(N__49865),
            .I(N__49859));
    LocalMux I__12506 (
            .O(N__49862),
            .I(N__49854));
    LocalMux I__12505 (
            .O(N__49859),
            .I(N__49854));
    Odrv4 I__12504 (
            .O(N__49854),
            .I(data_out_9__2__N_367));
    ClkMux I__12503 (
            .O(N__49851),
            .I(N__49176));
    ClkMux I__12502 (
            .O(N__49850),
            .I(N__49176));
    ClkMux I__12501 (
            .O(N__49849),
            .I(N__49176));
    ClkMux I__12500 (
            .O(N__49848),
            .I(N__49176));
    ClkMux I__12499 (
            .O(N__49847),
            .I(N__49176));
    ClkMux I__12498 (
            .O(N__49846),
            .I(N__49176));
    ClkMux I__12497 (
            .O(N__49845),
            .I(N__49176));
    ClkMux I__12496 (
            .O(N__49844),
            .I(N__49176));
    ClkMux I__12495 (
            .O(N__49843),
            .I(N__49176));
    ClkMux I__12494 (
            .O(N__49842),
            .I(N__49176));
    ClkMux I__12493 (
            .O(N__49841),
            .I(N__49176));
    ClkMux I__12492 (
            .O(N__49840),
            .I(N__49176));
    ClkMux I__12491 (
            .O(N__49839),
            .I(N__49176));
    ClkMux I__12490 (
            .O(N__49838),
            .I(N__49176));
    ClkMux I__12489 (
            .O(N__49837),
            .I(N__49176));
    ClkMux I__12488 (
            .O(N__49836),
            .I(N__49176));
    ClkMux I__12487 (
            .O(N__49835),
            .I(N__49176));
    ClkMux I__12486 (
            .O(N__49834),
            .I(N__49176));
    ClkMux I__12485 (
            .O(N__49833),
            .I(N__49176));
    ClkMux I__12484 (
            .O(N__49832),
            .I(N__49176));
    ClkMux I__12483 (
            .O(N__49831),
            .I(N__49176));
    ClkMux I__12482 (
            .O(N__49830),
            .I(N__49176));
    ClkMux I__12481 (
            .O(N__49829),
            .I(N__49176));
    ClkMux I__12480 (
            .O(N__49828),
            .I(N__49176));
    ClkMux I__12479 (
            .O(N__49827),
            .I(N__49176));
    ClkMux I__12478 (
            .O(N__49826),
            .I(N__49176));
    ClkMux I__12477 (
            .O(N__49825),
            .I(N__49176));
    ClkMux I__12476 (
            .O(N__49824),
            .I(N__49176));
    ClkMux I__12475 (
            .O(N__49823),
            .I(N__49176));
    ClkMux I__12474 (
            .O(N__49822),
            .I(N__49176));
    ClkMux I__12473 (
            .O(N__49821),
            .I(N__49176));
    ClkMux I__12472 (
            .O(N__49820),
            .I(N__49176));
    ClkMux I__12471 (
            .O(N__49819),
            .I(N__49176));
    ClkMux I__12470 (
            .O(N__49818),
            .I(N__49176));
    ClkMux I__12469 (
            .O(N__49817),
            .I(N__49176));
    ClkMux I__12468 (
            .O(N__49816),
            .I(N__49176));
    ClkMux I__12467 (
            .O(N__49815),
            .I(N__49176));
    ClkMux I__12466 (
            .O(N__49814),
            .I(N__49176));
    ClkMux I__12465 (
            .O(N__49813),
            .I(N__49176));
    ClkMux I__12464 (
            .O(N__49812),
            .I(N__49176));
    ClkMux I__12463 (
            .O(N__49811),
            .I(N__49176));
    ClkMux I__12462 (
            .O(N__49810),
            .I(N__49176));
    ClkMux I__12461 (
            .O(N__49809),
            .I(N__49176));
    ClkMux I__12460 (
            .O(N__49808),
            .I(N__49176));
    ClkMux I__12459 (
            .O(N__49807),
            .I(N__49176));
    ClkMux I__12458 (
            .O(N__49806),
            .I(N__49176));
    ClkMux I__12457 (
            .O(N__49805),
            .I(N__49176));
    ClkMux I__12456 (
            .O(N__49804),
            .I(N__49176));
    ClkMux I__12455 (
            .O(N__49803),
            .I(N__49176));
    ClkMux I__12454 (
            .O(N__49802),
            .I(N__49176));
    ClkMux I__12453 (
            .O(N__49801),
            .I(N__49176));
    ClkMux I__12452 (
            .O(N__49800),
            .I(N__49176));
    ClkMux I__12451 (
            .O(N__49799),
            .I(N__49176));
    ClkMux I__12450 (
            .O(N__49798),
            .I(N__49176));
    ClkMux I__12449 (
            .O(N__49797),
            .I(N__49176));
    ClkMux I__12448 (
            .O(N__49796),
            .I(N__49176));
    ClkMux I__12447 (
            .O(N__49795),
            .I(N__49176));
    ClkMux I__12446 (
            .O(N__49794),
            .I(N__49176));
    ClkMux I__12445 (
            .O(N__49793),
            .I(N__49176));
    ClkMux I__12444 (
            .O(N__49792),
            .I(N__49176));
    ClkMux I__12443 (
            .O(N__49791),
            .I(N__49176));
    ClkMux I__12442 (
            .O(N__49790),
            .I(N__49176));
    ClkMux I__12441 (
            .O(N__49789),
            .I(N__49176));
    ClkMux I__12440 (
            .O(N__49788),
            .I(N__49176));
    ClkMux I__12439 (
            .O(N__49787),
            .I(N__49176));
    ClkMux I__12438 (
            .O(N__49786),
            .I(N__49176));
    ClkMux I__12437 (
            .O(N__49785),
            .I(N__49176));
    ClkMux I__12436 (
            .O(N__49784),
            .I(N__49176));
    ClkMux I__12435 (
            .O(N__49783),
            .I(N__49176));
    ClkMux I__12434 (
            .O(N__49782),
            .I(N__49176));
    ClkMux I__12433 (
            .O(N__49781),
            .I(N__49176));
    ClkMux I__12432 (
            .O(N__49780),
            .I(N__49176));
    ClkMux I__12431 (
            .O(N__49779),
            .I(N__49176));
    ClkMux I__12430 (
            .O(N__49778),
            .I(N__49176));
    ClkMux I__12429 (
            .O(N__49777),
            .I(N__49176));
    ClkMux I__12428 (
            .O(N__49776),
            .I(N__49176));
    ClkMux I__12427 (
            .O(N__49775),
            .I(N__49176));
    ClkMux I__12426 (
            .O(N__49774),
            .I(N__49176));
    ClkMux I__12425 (
            .O(N__49773),
            .I(N__49176));
    ClkMux I__12424 (
            .O(N__49772),
            .I(N__49176));
    ClkMux I__12423 (
            .O(N__49771),
            .I(N__49176));
    ClkMux I__12422 (
            .O(N__49770),
            .I(N__49176));
    ClkMux I__12421 (
            .O(N__49769),
            .I(N__49176));
    ClkMux I__12420 (
            .O(N__49768),
            .I(N__49176));
    ClkMux I__12419 (
            .O(N__49767),
            .I(N__49176));
    ClkMux I__12418 (
            .O(N__49766),
            .I(N__49176));
    ClkMux I__12417 (
            .O(N__49765),
            .I(N__49176));
    ClkMux I__12416 (
            .O(N__49764),
            .I(N__49176));
    ClkMux I__12415 (
            .O(N__49763),
            .I(N__49176));
    ClkMux I__12414 (
            .O(N__49762),
            .I(N__49176));
    ClkMux I__12413 (
            .O(N__49761),
            .I(N__49176));
    ClkMux I__12412 (
            .O(N__49760),
            .I(N__49176));
    ClkMux I__12411 (
            .O(N__49759),
            .I(N__49176));
    ClkMux I__12410 (
            .O(N__49758),
            .I(N__49176));
    ClkMux I__12409 (
            .O(N__49757),
            .I(N__49176));
    ClkMux I__12408 (
            .O(N__49756),
            .I(N__49176));
    ClkMux I__12407 (
            .O(N__49755),
            .I(N__49176));
    ClkMux I__12406 (
            .O(N__49754),
            .I(N__49176));
    ClkMux I__12405 (
            .O(N__49753),
            .I(N__49176));
    ClkMux I__12404 (
            .O(N__49752),
            .I(N__49176));
    ClkMux I__12403 (
            .O(N__49751),
            .I(N__49176));
    ClkMux I__12402 (
            .O(N__49750),
            .I(N__49176));
    ClkMux I__12401 (
            .O(N__49749),
            .I(N__49176));
    ClkMux I__12400 (
            .O(N__49748),
            .I(N__49176));
    ClkMux I__12399 (
            .O(N__49747),
            .I(N__49176));
    ClkMux I__12398 (
            .O(N__49746),
            .I(N__49176));
    ClkMux I__12397 (
            .O(N__49745),
            .I(N__49176));
    ClkMux I__12396 (
            .O(N__49744),
            .I(N__49176));
    ClkMux I__12395 (
            .O(N__49743),
            .I(N__49176));
    ClkMux I__12394 (
            .O(N__49742),
            .I(N__49176));
    ClkMux I__12393 (
            .O(N__49741),
            .I(N__49176));
    ClkMux I__12392 (
            .O(N__49740),
            .I(N__49176));
    ClkMux I__12391 (
            .O(N__49739),
            .I(N__49176));
    ClkMux I__12390 (
            .O(N__49738),
            .I(N__49176));
    ClkMux I__12389 (
            .O(N__49737),
            .I(N__49176));
    ClkMux I__12388 (
            .O(N__49736),
            .I(N__49176));
    ClkMux I__12387 (
            .O(N__49735),
            .I(N__49176));
    ClkMux I__12386 (
            .O(N__49734),
            .I(N__49176));
    ClkMux I__12385 (
            .O(N__49733),
            .I(N__49176));
    ClkMux I__12384 (
            .O(N__49732),
            .I(N__49176));
    ClkMux I__12383 (
            .O(N__49731),
            .I(N__49176));
    ClkMux I__12382 (
            .O(N__49730),
            .I(N__49176));
    ClkMux I__12381 (
            .O(N__49729),
            .I(N__49176));
    ClkMux I__12380 (
            .O(N__49728),
            .I(N__49176));
    ClkMux I__12379 (
            .O(N__49727),
            .I(N__49176));
    ClkMux I__12378 (
            .O(N__49726),
            .I(N__49176));
    ClkMux I__12377 (
            .O(N__49725),
            .I(N__49176));
    ClkMux I__12376 (
            .O(N__49724),
            .I(N__49176));
    ClkMux I__12375 (
            .O(N__49723),
            .I(N__49176));
    ClkMux I__12374 (
            .O(N__49722),
            .I(N__49176));
    ClkMux I__12373 (
            .O(N__49721),
            .I(N__49176));
    ClkMux I__12372 (
            .O(N__49720),
            .I(N__49176));
    ClkMux I__12371 (
            .O(N__49719),
            .I(N__49176));
    ClkMux I__12370 (
            .O(N__49718),
            .I(N__49176));
    ClkMux I__12369 (
            .O(N__49717),
            .I(N__49176));
    ClkMux I__12368 (
            .O(N__49716),
            .I(N__49176));
    ClkMux I__12367 (
            .O(N__49715),
            .I(N__49176));
    ClkMux I__12366 (
            .O(N__49714),
            .I(N__49176));
    ClkMux I__12365 (
            .O(N__49713),
            .I(N__49176));
    ClkMux I__12364 (
            .O(N__49712),
            .I(N__49176));
    ClkMux I__12363 (
            .O(N__49711),
            .I(N__49176));
    ClkMux I__12362 (
            .O(N__49710),
            .I(N__49176));
    ClkMux I__12361 (
            .O(N__49709),
            .I(N__49176));
    ClkMux I__12360 (
            .O(N__49708),
            .I(N__49176));
    ClkMux I__12359 (
            .O(N__49707),
            .I(N__49176));
    ClkMux I__12358 (
            .O(N__49706),
            .I(N__49176));
    ClkMux I__12357 (
            .O(N__49705),
            .I(N__49176));
    ClkMux I__12356 (
            .O(N__49704),
            .I(N__49176));
    ClkMux I__12355 (
            .O(N__49703),
            .I(N__49176));
    ClkMux I__12354 (
            .O(N__49702),
            .I(N__49176));
    ClkMux I__12353 (
            .O(N__49701),
            .I(N__49176));
    ClkMux I__12352 (
            .O(N__49700),
            .I(N__49176));
    ClkMux I__12351 (
            .O(N__49699),
            .I(N__49176));
    ClkMux I__12350 (
            .O(N__49698),
            .I(N__49176));
    ClkMux I__12349 (
            .O(N__49697),
            .I(N__49176));
    ClkMux I__12348 (
            .O(N__49696),
            .I(N__49176));
    ClkMux I__12347 (
            .O(N__49695),
            .I(N__49176));
    ClkMux I__12346 (
            .O(N__49694),
            .I(N__49176));
    ClkMux I__12345 (
            .O(N__49693),
            .I(N__49176));
    ClkMux I__12344 (
            .O(N__49692),
            .I(N__49176));
    ClkMux I__12343 (
            .O(N__49691),
            .I(N__49176));
    ClkMux I__12342 (
            .O(N__49690),
            .I(N__49176));
    ClkMux I__12341 (
            .O(N__49689),
            .I(N__49176));
    ClkMux I__12340 (
            .O(N__49688),
            .I(N__49176));
    ClkMux I__12339 (
            .O(N__49687),
            .I(N__49176));
    ClkMux I__12338 (
            .O(N__49686),
            .I(N__49176));
    ClkMux I__12337 (
            .O(N__49685),
            .I(N__49176));
    ClkMux I__12336 (
            .O(N__49684),
            .I(N__49176));
    ClkMux I__12335 (
            .O(N__49683),
            .I(N__49176));
    ClkMux I__12334 (
            .O(N__49682),
            .I(N__49176));
    ClkMux I__12333 (
            .O(N__49681),
            .I(N__49176));
    ClkMux I__12332 (
            .O(N__49680),
            .I(N__49176));
    ClkMux I__12331 (
            .O(N__49679),
            .I(N__49176));
    ClkMux I__12330 (
            .O(N__49678),
            .I(N__49176));
    ClkMux I__12329 (
            .O(N__49677),
            .I(N__49176));
    ClkMux I__12328 (
            .O(N__49676),
            .I(N__49176));
    ClkMux I__12327 (
            .O(N__49675),
            .I(N__49176));
    ClkMux I__12326 (
            .O(N__49674),
            .I(N__49176));
    ClkMux I__12325 (
            .O(N__49673),
            .I(N__49176));
    ClkMux I__12324 (
            .O(N__49672),
            .I(N__49176));
    ClkMux I__12323 (
            .O(N__49671),
            .I(N__49176));
    ClkMux I__12322 (
            .O(N__49670),
            .I(N__49176));
    ClkMux I__12321 (
            .O(N__49669),
            .I(N__49176));
    ClkMux I__12320 (
            .O(N__49668),
            .I(N__49176));
    ClkMux I__12319 (
            .O(N__49667),
            .I(N__49176));
    ClkMux I__12318 (
            .O(N__49666),
            .I(N__49176));
    ClkMux I__12317 (
            .O(N__49665),
            .I(N__49176));
    ClkMux I__12316 (
            .O(N__49664),
            .I(N__49176));
    ClkMux I__12315 (
            .O(N__49663),
            .I(N__49176));
    ClkMux I__12314 (
            .O(N__49662),
            .I(N__49176));
    ClkMux I__12313 (
            .O(N__49661),
            .I(N__49176));
    ClkMux I__12312 (
            .O(N__49660),
            .I(N__49176));
    ClkMux I__12311 (
            .O(N__49659),
            .I(N__49176));
    ClkMux I__12310 (
            .O(N__49658),
            .I(N__49176));
    ClkMux I__12309 (
            .O(N__49657),
            .I(N__49176));
    ClkMux I__12308 (
            .O(N__49656),
            .I(N__49176));
    ClkMux I__12307 (
            .O(N__49655),
            .I(N__49176));
    ClkMux I__12306 (
            .O(N__49654),
            .I(N__49176));
    ClkMux I__12305 (
            .O(N__49653),
            .I(N__49176));
    ClkMux I__12304 (
            .O(N__49652),
            .I(N__49176));
    ClkMux I__12303 (
            .O(N__49651),
            .I(N__49176));
    ClkMux I__12302 (
            .O(N__49650),
            .I(N__49176));
    ClkMux I__12301 (
            .O(N__49649),
            .I(N__49176));
    ClkMux I__12300 (
            .O(N__49648),
            .I(N__49176));
    ClkMux I__12299 (
            .O(N__49647),
            .I(N__49176));
    ClkMux I__12298 (
            .O(N__49646),
            .I(N__49176));
    ClkMux I__12297 (
            .O(N__49645),
            .I(N__49176));
    ClkMux I__12296 (
            .O(N__49644),
            .I(N__49176));
    ClkMux I__12295 (
            .O(N__49643),
            .I(N__49176));
    ClkMux I__12294 (
            .O(N__49642),
            .I(N__49176));
    ClkMux I__12293 (
            .O(N__49641),
            .I(N__49176));
    ClkMux I__12292 (
            .O(N__49640),
            .I(N__49176));
    ClkMux I__12291 (
            .O(N__49639),
            .I(N__49176));
    ClkMux I__12290 (
            .O(N__49638),
            .I(N__49176));
    ClkMux I__12289 (
            .O(N__49637),
            .I(N__49176));
    ClkMux I__12288 (
            .O(N__49636),
            .I(N__49176));
    ClkMux I__12287 (
            .O(N__49635),
            .I(N__49176));
    ClkMux I__12286 (
            .O(N__49634),
            .I(N__49176));
    ClkMux I__12285 (
            .O(N__49633),
            .I(N__49176));
    ClkMux I__12284 (
            .O(N__49632),
            .I(N__49176));
    ClkMux I__12283 (
            .O(N__49631),
            .I(N__49176));
    ClkMux I__12282 (
            .O(N__49630),
            .I(N__49176));
    ClkMux I__12281 (
            .O(N__49629),
            .I(N__49176));
    ClkMux I__12280 (
            .O(N__49628),
            .I(N__49176));
    ClkMux I__12279 (
            .O(N__49627),
            .I(N__49176));
    GlobalMux I__12278 (
            .O(N__49176),
            .I(N__49173));
    gio2CtrlBuf I__12277 (
            .O(N__49173),
            .I(CLK_c));
    InMux I__12276 (
            .O(N__49170),
            .I(N__49165));
    InMux I__12275 (
            .O(N__49169),
            .I(N__49162));
    InMux I__12274 (
            .O(N__49168),
            .I(N__49158));
    LocalMux I__12273 (
            .O(N__49165),
            .I(N__49155));
    LocalMux I__12272 (
            .O(N__49162),
            .I(N__49152));
    CascadeMux I__12271 (
            .O(N__49161),
            .I(N__49148));
    LocalMux I__12270 (
            .O(N__49158),
            .I(N__49144));
    Span4Mux_v I__12269 (
            .O(N__49155),
            .I(N__49141));
    Span4Mux_v I__12268 (
            .O(N__49152),
            .I(N__49138));
    InMux I__12267 (
            .O(N__49151),
            .I(N__49135));
    InMux I__12266 (
            .O(N__49148),
            .I(N__49132));
    InMux I__12265 (
            .O(N__49147),
            .I(N__49129));
    Span4Mux_v I__12264 (
            .O(N__49144),
            .I(N__49122));
    Span4Mux_h I__12263 (
            .O(N__49141),
            .I(N__49122));
    Span4Mux_h I__12262 (
            .O(N__49138),
            .I(N__49122));
    LocalMux I__12261 (
            .O(N__49135),
            .I(data_out_9_2));
    LocalMux I__12260 (
            .O(N__49132),
            .I(data_out_9_2));
    LocalMux I__12259 (
            .O(N__49129),
            .I(data_out_9_2));
    Odrv4 I__12258 (
            .O(N__49122),
            .I(data_out_9_2));
    InMux I__12257 (
            .O(N__49113),
            .I(N__49106));
    InMux I__12256 (
            .O(N__49112),
            .I(N__49103));
    InMux I__12255 (
            .O(N__49111),
            .I(N__49100));
    InMux I__12254 (
            .O(N__49110),
            .I(N__49094));
    InMux I__12253 (
            .O(N__49109),
            .I(N__49094));
    LocalMux I__12252 (
            .O(N__49106),
            .I(N__49091));
    LocalMux I__12251 (
            .O(N__49103),
            .I(N__49088));
    LocalMux I__12250 (
            .O(N__49100),
            .I(N__49085));
    InMux I__12249 (
            .O(N__49099),
            .I(N__49081));
    LocalMux I__12248 (
            .O(N__49094),
            .I(N__49078));
    Span4Mux_v I__12247 (
            .O(N__49091),
            .I(N__49075));
    Span4Mux_v I__12246 (
            .O(N__49088),
            .I(N__49072));
    Span4Mux_v I__12245 (
            .O(N__49085),
            .I(N__49069));
    InMux I__12244 (
            .O(N__49084),
            .I(N__49066));
    LocalMux I__12243 (
            .O(N__49081),
            .I(N__49060));
    Span4Mux_h I__12242 (
            .O(N__49078),
            .I(N__49060));
    Sp12to4 I__12241 (
            .O(N__49075),
            .I(N__49051));
    Sp12to4 I__12240 (
            .O(N__49072),
            .I(N__49051));
    Sp12to4 I__12239 (
            .O(N__49069),
            .I(N__49051));
    LocalMux I__12238 (
            .O(N__49066),
            .I(N__49051));
    InMux I__12237 (
            .O(N__49065),
            .I(N__49048));
    Odrv4 I__12236 (
            .O(N__49060),
            .I(\c0.data_out_5_4 ));
    Odrv12 I__12235 (
            .O(N__49051),
            .I(\c0.data_out_5_4 ));
    LocalMux I__12234 (
            .O(N__49048),
            .I(\c0.data_out_5_4 ));
    InMux I__12233 (
            .O(N__49041),
            .I(N__49037));
    CascadeMux I__12232 (
            .O(N__49040),
            .I(N__49034));
    LocalMux I__12231 (
            .O(N__49037),
            .I(N__49030));
    InMux I__12230 (
            .O(N__49034),
            .I(N__49025));
    InMux I__12229 (
            .O(N__49033),
            .I(N__49025));
    Span4Mux_v I__12228 (
            .O(N__49030),
            .I(N__49022));
    LocalMux I__12227 (
            .O(N__49025),
            .I(N__49019));
    Odrv4 I__12226 (
            .O(N__49022),
            .I(\c0.data_out_10_6 ));
    Odrv4 I__12225 (
            .O(N__49019),
            .I(\c0.data_out_10_6 ));
    InMux I__12224 (
            .O(N__49014),
            .I(N__49010));
    InMux I__12223 (
            .O(N__49013),
            .I(N__49007));
    LocalMux I__12222 (
            .O(N__49010),
            .I(N__49000));
    LocalMux I__12221 (
            .O(N__49007),
            .I(N__49000));
    InMux I__12220 (
            .O(N__49006),
            .I(N__48997));
    InMux I__12219 (
            .O(N__49005),
            .I(N__48994));
    Span4Mux_v I__12218 (
            .O(N__49000),
            .I(N__48991));
    LocalMux I__12217 (
            .O(N__48997),
            .I(N__48988));
    LocalMux I__12216 (
            .O(N__48994),
            .I(\c0.data_out_9_3 ));
    Odrv4 I__12215 (
            .O(N__48991),
            .I(\c0.data_out_9_3 ));
    Odrv4 I__12214 (
            .O(N__48988),
            .I(\c0.data_out_9_3 ));
    CascadeMux I__12213 (
            .O(N__48981),
            .I(\c0.n10204_cascade_ ));
    InMux I__12212 (
            .O(N__48978),
            .I(N__48975));
    LocalMux I__12211 (
            .O(N__48975),
            .I(N__48972));
    Span4Mux_v I__12210 (
            .O(N__48972),
            .I(N__48968));
    InMux I__12209 (
            .O(N__48971),
            .I(N__48965));
    Sp12to4 I__12208 (
            .O(N__48968),
            .I(N__48958));
    LocalMux I__12207 (
            .O(N__48965),
            .I(N__48958));
    InMux I__12206 (
            .O(N__48964),
            .I(N__48953));
    InMux I__12205 (
            .O(N__48963),
            .I(N__48953));
    Odrv12 I__12204 (
            .O(N__48958),
            .I(\c0.data_out_7_4 ));
    LocalMux I__12203 (
            .O(N__48953),
            .I(\c0.data_out_7_4 ));
    CascadeMux I__12202 (
            .O(N__48948),
            .I(N__48945));
    InMux I__12201 (
            .O(N__48945),
            .I(N__48942));
    LocalMux I__12200 (
            .O(N__48942),
            .I(N__48939));
    Span4Mux_v I__12199 (
            .O(N__48939),
            .I(N__48936));
    Odrv4 I__12198 (
            .O(N__48936),
            .I(\c0.n10_adj_2172 ));
    InMux I__12197 (
            .O(N__48933),
            .I(N__48930));
    LocalMux I__12196 (
            .O(N__48930),
            .I(N__48927));
    Span4Mux_h I__12195 (
            .O(N__48927),
            .I(N__48922));
    InMux I__12194 (
            .O(N__48926),
            .I(N__48919));
    InMux I__12193 (
            .O(N__48925),
            .I(N__48916));
    Span4Mux_h I__12192 (
            .O(N__48922),
            .I(N__48913));
    LocalMux I__12191 (
            .O(N__48919),
            .I(N__48908));
    LocalMux I__12190 (
            .O(N__48916),
            .I(N__48908));
    Odrv4 I__12189 (
            .O(N__48913),
            .I(\c0.data_out_6_7 ));
    Odrv12 I__12188 (
            .O(N__48908),
            .I(\c0.data_out_6_7 ));
    InMux I__12187 (
            .O(N__48903),
            .I(N__48900));
    LocalMux I__12186 (
            .O(N__48900),
            .I(N__48897));
    Span4Mux_h I__12185 (
            .O(N__48897),
            .I(N__48893));
    InMux I__12184 (
            .O(N__48896),
            .I(N__48890));
    Odrv4 I__12183 (
            .O(N__48893),
            .I(\c0.n26_adj_2165 ));
    LocalMux I__12182 (
            .O(N__48890),
            .I(\c0.n26_adj_2165 ));
    InMux I__12181 (
            .O(N__48885),
            .I(N__48880));
    InMux I__12180 (
            .O(N__48884),
            .I(N__48877));
    InMux I__12179 (
            .O(N__48883),
            .I(N__48874));
    LocalMux I__12178 (
            .O(N__48880),
            .I(N__48871));
    LocalMux I__12177 (
            .O(N__48877),
            .I(N__48868));
    LocalMux I__12176 (
            .O(N__48874),
            .I(N__48865));
    Span4Mux_v I__12175 (
            .O(N__48871),
            .I(N__48861));
    Span4Mux_h I__12174 (
            .O(N__48868),
            .I(N__48858));
    Span4Mux_h I__12173 (
            .O(N__48865),
            .I(N__48855));
    InMux I__12172 (
            .O(N__48864),
            .I(N__48852));
    Span4Mux_h I__12171 (
            .O(N__48861),
            .I(N__48849));
    Span4Mux_h I__12170 (
            .O(N__48858),
            .I(N__48844));
    Span4Mux_v I__12169 (
            .O(N__48855),
            .I(N__48844));
    LocalMux I__12168 (
            .O(N__48852),
            .I(N__48841));
    Odrv4 I__12167 (
            .O(N__48849),
            .I(\c0.data_out_6_5 ));
    Odrv4 I__12166 (
            .O(N__48844),
            .I(\c0.data_out_6_5 ));
    Odrv4 I__12165 (
            .O(N__48841),
            .I(\c0.data_out_6_5 ));
    InMux I__12164 (
            .O(N__48834),
            .I(N__48831));
    LocalMux I__12163 (
            .O(N__48831),
            .I(N__48828));
    Span4Mux_v I__12162 (
            .O(N__48828),
            .I(N__48822));
    InMux I__12161 (
            .O(N__48827),
            .I(N__48819));
    InMux I__12160 (
            .O(N__48826),
            .I(N__48816));
    InMux I__12159 (
            .O(N__48825),
            .I(N__48812));
    Sp12to4 I__12158 (
            .O(N__48822),
            .I(N__48805));
    LocalMux I__12157 (
            .O(N__48819),
            .I(N__48805));
    LocalMux I__12156 (
            .O(N__48816),
            .I(N__48805));
    InMux I__12155 (
            .O(N__48815),
            .I(N__48802));
    LocalMux I__12154 (
            .O(N__48812),
            .I(data_out_8_3));
    Odrv12 I__12153 (
            .O(N__48805),
            .I(data_out_8_3));
    LocalMux I__12152 (
            .O(N__48802),
            .I(data_out_8_3));
    CascadeMux I__12151 (
            .O(N__48795),
            .I(\c0.n10_adj_2166_cascade_ ));
    CascadeMux I__12150 (
            .O(N__48792),
            .I(N__48788));
    InMux I__12149 (
            .O(N__48791),
            .I(N__48785));
    InMux I__12148 (
            .O(N__48788),
            .I(N__48782));
    LocalMux I__12147 (
            .O(N__48785),
            .I(N__48779));
    LocalMux I__12146 (
            .O(N__48782),
            .I(\c0.n10170 ));
    Odrv4 I__12145 (
            .O(N__48779),
            .I(\c0.n10170 ));
    InMux I__12144 (
            .O(N__48774),
            .I(N__48771));
    LocalMux I__12143 (
            .O(N__48771),
            .I(N__48767));
    InMux I__12142 (
            .O(N__48770),
            .I(N__48764));
    Odrv12 I__12141 (
            .O(N__48767),
            .I(\c0.n17252 ));
    LocalMux I__12140 (
            .O(N__48764),
            .I(\c0.n17252 ));
    CascadeMux I__12139 (
            .O(N__48759),
            .I(N__48756));
    InMux I__12138 (
            .O(N__48756),
            .I(N__48753));
    LocalMux I__12137 (
            .O(N__48753),
            .I(N__48750));
    Span4Mux_v I__12136 (
            .O(N__48750),
            .I(N__48747));
    Span4Mux_h I__12135 (
            .O(N__48747),
            .I(N__48742));
    InMux I__12134 (
            .O(N__48746),
            .I(N__48737));
    InMux I__12133 (
            .O(N__48745),
            .I(N__48737));
    Odrv4 I__12132 (
            .O(N__48742),
            .I(data_out_10_1));
    LocalMux I__12131 (
            .O(N__48737),
            .I(data_out_10_1));
    InMux I__12130 (
            .O(N__48732),
            .I(N__48729));
    LocalMux I__12129 (
            .O(N__48729),
            .I(N__48725));
    InMux I__12128 (
            .O(N__48728),
            .I(N__48722));
    Span4Mux_h I__12127 (
            .O(N__48725),
            .I(N__48719));
    LocalMux I__12126 (
            .O(N__48722),
            .I(N__48714));
    Span4Mux_h I__12125 (
            .O(N__48719),
            .I(N__48710));
    InMux I__12124 (
            .O(N__48718),
            .I(N__48707));
    InMux I__12123 (
            .O(N__48717),
            .I(N__48704));
    Span4Mux_h I__12122 (
            .O(N__48714),
            .I(N__48701));
    InMux I__12121 (
            .O(N__48713),
            .I(N__48698));
    Odrv4 I__12120 (
            .O(N__48710),
            .I(data_out_8_2));
    LocalMux I__12119 (
            .O(N__48707),
            .I(data_out_8_2));
    LocalMux I__12118 (
            .O(N__48704),
            .I(data_out_8_2));
    Odrv4 I__12117 (
            .O(N__48701),
            .I(data_out_8_2));
    LocalMux I__12116 (
            .O(N__48698),
            .I(data_out_8_2));
    CascadeMux I__12115 (
            .O(N__48687),
            .I(N__48684));
    InMux I__12114 (
            .O(N__48684),
            .I(N__48680));
    InMux I__12113 (
            .O(N__48683),
            .I(N__48677));
    LocalMux I__12112 (
            .O(N__48680),
            .I(N__48674));
    LocalMux I__12111 (
            .O(N__48677),
            .I(N__48668));
    Span4Mux_s3_v I__12110 (
            .O(N__48674),
            .I(N__48668));
    InMux I__12109 (
            .O(N__48673),
            .I(N__48665));
    Odrv4 I__12108 (
            .O(N__48668),
            .I(\c0.data_out_10_5 ));
    LocalMux I__12107 (
            .O(N__48665),
            .I(\c0.data_out_10_5 ));
    InMux I__12106 (
            .O(N__48660),
            .I(N__48656));
    InMux I__12105 (
            .O(N__48659),
            .I(N__48653));
    LocalMux I__12104 (
            .O(N__48656),
            .I(N__48647));
    LocalMux I__12103 (
            .O(N__48653),
            .I(N__48647));
    InMux I__12102 (
            .O(N__48652),
            .I(N__48644));
    Span4Mux_v I__12101 (
            .O(N__48647),
            .I(N__48641));
    LocalMux I__12100 (
            .O(N__48644),
            .I(N__48638));
    Span4Mux_h I__12099 (
            .O(N__48641),
            .I(N__48635));
    Span4Mux_h I__12098 (
            .O(N__48638),
            .I(N__48632));
    Span4Mux_h I__12097 (
            .O(N__48635),
            .I(N__48629));
    Span4Mux_h I__12096 (
            .O(N__48632),
            .I(N__48626));
    Odrv4 I__12095 (
            .O(N__48629),
            .I(\c0.data_out_7_1 ));
    Odrv4 I__12094 (
            .O(N__48626),
            .I(\c0.data_out_7_1 ));
    InMux I__12093 (
            .O(N__48621),
            .I(N__48617));
    CascadeMux I__12092 (
            .O(N__48620),
            .I(N__48611));
    LocalMux I__12091 (
            .O(N__48617),
            .I(N__48608));
    InMux I__12090 (
            .O(N__48616),
            .I(N__48603));
    InMux I__12089 (
            .O(N__48615),
            .I(N__48603));
    InMux I__12088 (
            .O(N__48614),
            .I(N__48598));
    InMux I__12087 (
            .O(N__48611),
            .I(N__48598));
    Odrv4 I__12086 (
            .O(N__48608),
            .I(\c0.data_out_9_0 ));
    LocalMux I__12085 (
            .O(N__48603),
            .I(\c0.data_out_9_0 ));
    LocalMux I__12084 (
            .O(N__48598),
            .I(\c0.data_out_9_0 ));
    InMux I__12083 (
            .O(N__48591),
            .I(N__48588));
    LocalMux I__12082 (
            .O(N__48588),
            .I(N__48585));
    Odrv4 I__12081 (
            .O(N__48585),
            .I(\c0.n6_adj_2169 ));
    InMux I__12080 (
            .O(N__48582),
            .I(N__48579));
    LocalMux I__12079 (
            .O(N__48579),
            .I(\c0.n17162 ));
    CascadeMux I__12078 (
            .O(N__48576),
            .I(\c0.n17150_cascade_ ));
    InMux I__12077 (
            .O(N__48573),
            .I(N__48567));
    InMux I__12076 (
            .O(N__48572),
            .I(N__48561));
    InMux I__12075 (
            .O(N__48571),
            .I(N__48561));
    InMux I__12074 (
            .O(N__48570),
            .I(N__48558));
    LocalMux I__12073 (
            .O(N__48567),
            .I(N__48555));
    InMux I__12072 (
            .O(N__48566),
            .I(N__48552));
    LocalMux I__12071 (
            .O(N__48561),
            .I(N__48549));
    LocalMux I__12070 (
            .O(N__48558),
            .I(N__48546));
    Span4Mux_h I__12069 (
            .O(N__48555),
            .I(N__48543));
    LocalMux I__12068 (
            .O(N__48552),
            .I(\c0.data_out_9_1 ));
    Odrv4 I__12067 (
            .O(N__48549),
            .I(\c0.data_out_9_1 ));
    Odrv4 I__12066 (
            .O(N__48546),
            .I(\c0.data_out_9_1 ));
    Odrv4 I__12065 (
            .O(N__48543),
            .I(\c0.data_out_9_1 ));
    InMux I__12064 (
            .O(N__48534),
            .I(N__48529));
    InMux I__12063 (
            .O(N__48533),
            .I(N__48526));
    InMux I__12062 (
            .O(N__48532),
            .I(N__48523));
    LocalMux I__12061 (
            .O(N__48529),
            .I(N__48518));
    LocalMux I__12060 (
            .O(N__48526),
            .I(N__48518));
    LocalMux I__12059 (
            .O(N__48523),
            .I(N__48513));
    Span4Mux_h I__12058 (
            .O(N__48518),
            .I(N__48513));
    Odrv4 I__12057 (
            .O(N__48513),
            .I(\c0.data_out_9_5 ));
    InMux I__12056 (
            .O(N__48510),
            .I(N__48507));
    LocalMux I__12055 (
            .O(N__48507),
            .I(N__48504));
    Span4Mux_h I__12054 (
            .O(N__48504),
            .I(N__48501));
    Span4Mux_v I__12053 (
            .O(N__48501),
            .I(N__48497));
    InMux I__12052 (
            .O(N__48500),
            .I(N__48494));
    Sp12to4 I__12051 (
            .O(N__48497),
            .I(N__48489));
    LocalMux I__12050 (
            .O(N__48494),
            .I(N__48489));
    Span12Mux_h I__12049 (
            .O(N__48489),
            .I(N__48486));
    Odrv12 I__12048 (
            .O(N__48486),
            .I(\c0.n17110 ));
    InMux I__12047 (
            .O(N__48483),
            .I(N__48477));
    InMux I__12046 (
            .O(N__48482),
            .I(N__48477));
    LocalMux I__12045 (
            .O(N__48477),
            .I(N__48474));
    Sp12to4 I__12044 (
            .O(N__48474),
            .I(N__48469));
    InMux I__12043 (
            .O(N__48473),
            .I(N__48466));
    InMux I__12042 (
            .O(N__48472),
            .I(N__48462));
    Span12Mux_s5_v I__12041 (
            .O(N__48469),
            .I(N__48457));
    LocalMux I__12040 (
            .O(N__48466),
            .I(N__48457));
    InMux I__12039 (
            .O(N__48465),
            .I(N__48454));
    LocalMux I__12038 (
            .O(N__48462),
            .I(data_out_8_4));
    Odrv12 I__12037 (
            .O(N__48457),
            .I(data_out_8_4));
    LocalMux I__12036 (
            .O(N__48454),
            .I(data_out_8_4));
    InMux I__12035 (
            .O(N__48447),
            .I(N__48443));
    InMux I__12034 (
            .O(N__48446),
            .I(N__48440));
    LocalMux I__12033 (
            .O(N__48443),
            .I(N__48437));
    LocalMux I__12032 (
            .O(N__48440),
            .I(N__48434));
    Span4Mux_h I__12031 (
            .O(N__48437),
            .I(N__48431));
    Odrv4 I__12030 (
            .O(N__48434),
            .I(\c0.data_out_10_7 ));
    Odrv4 I__12029 (
            .O(N__48431),
            .I(\c0.data_out_10_7 ));
    InMux I__12028 (
            .O(N__48426),
            .I(N__48422));
    InMux I__12027 (
            .O(N__48425),
            .I(N__48413));
    LocalMux I__12026 (
            .O(N__48422),
            .I(N__48406));
    InMux I__12025 (
            .O(N__48421),
            .I(N__48401));
    InMux I__12024 (
            .O(N__48420),
            .I(N__48396));
    InMux I__12023 (
            .O(N__48419),
            .I(N__48396));
    CascadeMux I__12022 (
            .O(N__48418),
            .I(N__48393));
    CascadeMux I__12021 (
            .O(N__48417),
            .I(N__48389));
    InMux I__12020 (
            .O(N__48416),
            .I(N__48385));
    LocalMux I__12019 (
            .O(N__48413),
            .I(N__48376));
    InMux I__12018 (
            .O(N__48412),
            .I(N__48373));
    CascadeMux I__12017 (
            .O(N__48411),
            .I(N__48368));
    CascadeMux I__12016 (
            .O(N__48410),
            .I(N__48365));
    InMux I__12015 (
            .O(N__48409),
            .I(N__48362));
    Span4Mux_h I__12014 (
            .O(N__48406),
            .I(N__48359));
    InMux I__12013 (
            .O(N__48405),
            .I(N__48356));
    CascadeMux I__12012 (
            .O(N__48404),
            .I(N__48353));
    LocalMux I__12011 (
            .O(N__48401),
            .I(N__48348));
    LocalMux I__12010 (
            .O(N__48396),
            .I(N__48348));
    InMux I__12009 (
            .O(N__48393),
            .I(N__48343));
    InMux I__12008 (
            .O(N__48392),
            .I(N__48343));
    InMux I__12007 (
            .O(N__48389),
            .I(N__48340));
    InMux I__12006 (
            .O(N__48388),
            .I(N__48337));
    LocalMux I__12005 (
            .O(N__48385),
            .I(N__48334));
    InMux I__12004 (
            .O(N__48384),
            .I(N__48331));
    InMux I__12003 (
            .O(N__48383),
            .I(N__48328));
    InMux I__12002 (
            .O(N__48382),
            .I(N__48325));
    InMux I__12001 (
            .O(N__48381),
            .I(N__48322));
    InMux I__12000 (
            .O(N__48380),
            .I(N__48319));
    CascadeMux I__11999 (
            .O(N__48379),
            .I(N__48316));
    Span4Mux_v I__11998 (
            .O(N__48376),
            .I(N__48310));
    LocalMux I__11997 (
            .O(N__48373),
            .I(N__48307));
    InMux I__11996 (
            .O(N__48372),
            .I(N__48304));
    CascadeMux I__11995 (
            .O(N__48371),
            .I(N__48299));
    InMux I__11994 (
            .O(N__48368),
            .I(N__48295));
    InMux I__11993 (
            .O(N__48365),
            .I(N__48292));
    LocalMux I__11992 (
            .O(N__48362),
            .I(N__48285));
    Span4Mux_h I__11991 (
            .O(N__48359),
            .I(N__48285));
    LocalMux I__11990 (
            .O(N__48356),
            .I(N__48285));
    InMux I__11989 (
            .O(N__48353),
            .I(N__48282));
    Span4Mux_h I__11988 (
            .O(N__48348),
            .I(N__48279));
    LocalMux I__11987 (
            .O(N__48343),
            .I(N__48273));
    LocalMux I__11986 (
            .O(N__48340),
            .I(N__48264));
    LocalMux I__11985 (
            .O(N__48337),
            .I(N__48264));
    Span4Mux_h I__11984 (
            .O(N__48334),
            .I(N__48264));
    LocalMux I__11983 (
            .O(N__48331),
            .I(N__48264));
    LocalMux I__11982 (
            .O(N__48328),
            .I(N__48259));
    LocalMux I__11981 (
            .O(N__48325),
            .I(N__48259));
    LocalMux I__11980 (
            .O(N__48322),
            .I(N__48254));
    LocalMux I__11979 (
            .O(N__48319),
            .I(N__48254));
    InMux I__11978 (
            .O(N__48316),
            .I(N__48247));
    InMux I__11977 (
            .O(N__48315),
            .I(N__48247));
    InMux I__11976 (
            .O(N__48314),
            .I(N__48247));
    InMux I__11975 (
            .O(N__48313),
            .I(N__48244));
    Span4Mux_h I__11974 (
            .O(N__48310),
            .I(N__48241));
    Span4Mux_v I__11973 (
            .O(N__48307),
            .I(N__48236));
    LocalMux I__11972 (
            .O(N__48304),
            .I(N__48236));
    InMux I__11971 (
            .O(N__48303),
            .I(N__48233));
    InMux I__11970 (
            .O(N__48302),
            .I(N__48230));
    InMux I__11969 (
            .O(N__48299),
            .I(N__48225));
    InMux I__11968 (
            .O(N__48298),
            .I(N__48225));
    LocalMux I__11967 (
            .O(N__48295),
            .I(N__48220));
    LocalMux I__11966 (
            .O(N__48292),
            .I(N__48220));
    Span4Mux_v I__11965 (
            .O(N__48285),
            .I(N__48217));
    LocalMux I__11964 (
            .O(N__48282),
            .I(N__48212));
    Span4Mux_h I__11963 (
            .O(N__48279),
            .I(N__48212));
    InMux I__11962 (
            .O(N__48278),
            .I(N__48205));
    InMux I__11961 (
            .O(N__48277),
            .I(N__48205));
    InMux I__11960 (
            .O(N__48276),
            .I(N__48205));
    Span4Mux_h I__11959 (
            .O(N__48273),
            .I(N__48198));
    Span4Mux_v I__11958 (
            .O(N__48264),
            .I(N__48198));
    Span4Mux_v I__11957 (
            .O(N__48259),
            .I(N__48198));
    Span4Mux_h I__11956 (
            .O(N__48254),
            .I(N__48187));
    LocalMux I__11955 (
            .O(N__48247),
            .I(N__48187));
    LocalMux I__11954 (
            .O(N__48244),
            .I(N__48187));
    Span4Mux_v I__11953 (
            .O(N__48241),
            .I(N__48187));
    Span4Mux_h I__11952 (
            .O(N__48236),
            .I(N__48187));
    LocalMux I__11951 (
            .O(N__48233),
            .I(UART_TRANSMITTER_state_2));
    LocalMux I__11950 (
            .O(N__48230),
            .I(UART_TRANSMITTER_state_2));
    LocalMux I__11949 (
            .O(N__48225),
            .I(UART_TRANSMITTER_state_2));
    Odrv12 I__11948 (
            .O(N__48220),
            .I(UART_TRANSMITTER_state_2));
    Odrv4 I__11947 (
            .O(N__48217),
            .I(UART_TRANSMITTER_state_2));
    Odrv4 I__11946 (
            .O(N__48212),
            .I(UART_TRANSMITTER_state_2));
    LocalMux I__11945 (
            .O(N__48205),
            .I(UART_TRANSMITTER_state_2));
    Odrv4 I__11944 (
            .O(N__48198),
            .I(UART_TRANSMITTER_state_2));
    Odrv4 I__11943 (
            .O(N__48187),
            .I(UART_TRANSMITTER_state_2));
    InMux I__11942 (
            .O(N__48168),
            .I(N__48161));
    InMux I__11941 (
            .O(N__48167),
            .I(N__48158));
    InMux I__11940 (
            .O(N__48166),
            .I(N__48145));
    InMux I__11939 (
            .O(N__48165),
            .I(N__48145));
    InMux I__11938 (
            .O(N__48164),
            .I(N__48141));
    LocalMux I__11937 (
            .O(N__48161),
            .I(N__48138));
    LocalMux I__11936 (
            .O(N__48158),
            .I(N__48135));
    CascadeMux I__11935 (
            .O(N__48157),
            .I(N__48124));
    InMux I__11934 (
            .O(N__48156),
            .I(N__48118));
    CascadeMux I__11933 (
            .O(N__48155),
            .I(N__48115));
    InMux I__11932 (
            .O(N__48154),
            .I(N__48101));
    InMux I__11931 (
            .O(N__48153),
            .I(N__48101));
    InMux I__11930 (
            .O(N__48152),
            .I(N__48101));
    InMux I__11929 (
            .O(N__48151),
            .I(N__48101));
    InMux I__11928 (
            .O(N__48150),
            .I(N__48096));
    LocalMux I__11927 (
            .O(N__48145),
            .I(N__48093));
    CascadeMux I__11926 (
            .O(N__48144),
            .I(N__48090));
    LocalMux I__11925 (
            .O(N__48141),
            .I(N__48085));
    Span4Mux_v I__11924 (
            .O(N__48138),
            .I(N__48082));
    Span4Mux_v I__11923 (
            .O(N__48135),
            .I(N__48079));
    InMux I__11922 (
            .O(N__48134),
            .I(N__48076));
    InMux I__11921 (
            .O(N__48133),
            .I(N__48073));
    InMux I__11920 (
            .O(N__48132),
            .I(N__48066));
    InMux I__11919 (
            .O(N__48131),
            .I(N__48066));
    InMux I__11918 (
            .O(N__48130),
            .I(N__48066));
    InMux I__11917 (
            .O(N__48129),
            .I(N__48059));
    InMux I__11916 (
            .O(N__48128),
            .I(N__48059));
    InMux I__11915 (
            .O(N__48127),
            .I(N__48059));
    InMux I__11914 (
            .O(N__48124),
            .I(N__48050));
    InMux I__11913 (
            .O(N__48123),
            .I(N__48050));
    InMux I__11912 (
            .O(N__48122),
            .I(N__48050));
    InMux I__11911 (
            .O(N__48121),
            .I(N__48050));
    LocalMux I__11910 (
            .O(N__48118),
            .I(N__48047));
    InMux I__11909 (
            .O(N__48115),
            .I(N__48042));
    InMux I__11908 (
            .O(N__48114),
            .I(N__48042));
    InMux I__11907 (
            .O(N__48113),
            .I(N__48039));
    InMux I__11906 (
            .O(N__48112),
            .I(N__48036));
    InMux I__11905 (
            .O(N__48111),
            .I(N__48033));
    InMux I__11904 (
            .O(N__48110),
            .I(N__48029));
    LocalMux I__11903 (
            .O(N__48101),
            .I(N__48026));
    CascadeMux I__11902 (
            .O(N__48100),
            .I(N__48023));
    CascadeMux I__11901 (
            .O(N__48099),
            .I(N__48017));
    LocalMux I__11900 (
            .O(N__48096),
            .I(N__48014));
    Span12Mux_s8_v I__11899 (
            .O(N__48093),
            .I(N__48011));
    InMux I__11898 (
            .O(N__48090),
            .I(N__48008));
    InMux I__11897 (
            .O(N__48089),
            .I(N__48003));
    InMux I__11896 (
            .O(N__48088),
            .I(N__48003));
    Span4Mux_h I__11895 (
            .O(N__48085),
            .I(N__47996));
    Span4Mux_h I__11894 (
            .O(N__48082),
            .I(N__47996));
    Span4Mux_h I__11893 (
            .O(N__48079),
            .I(N__47996));
    LocalMux I__11892 (
            .O(N__48076),
            .I(N__47993));
    LocalMux I__11891 (
            .O(N__48073),
            .I(N__47990));
    LocalMux I__11890 (
            .O(N__48066),
            .I(N__47987));
    LocalMux I__11889 (
            .O(N__48059),
            .I(N__47978));
    LocalMux I__11888 (
            .O(N__48050),
            .I(N__47978));
    Span4Mux_h I__11887 (
            .O(N__48047),
            .I(N__47978));
    LocalMux I__11886 (
            .O(N__48042),
            .I(N__47978));
    LocalMux I__11885 (
            .O(N__48039),
            .I(N__47971));
    LocalMux I__11884 (
            .O(N__48036),
            .I(N__47971));
    LocalMux I__11883 (
            .O(N__48033),
            .I(N__47971));
    InMux I__11882 (
            .O(N__48032),
            .I(N__47968));
    LocalMux I__11881 (
            .O(N__48029),
            .I(N__47965));
    Span4Mux_h I__11880 (
            .O(N__48026),
            .I(N__47962));
    InMux I__11879 (
            .O(N__48023),
            .I(N__47959));
    InMux I__11878 (
            .O(N__48022),
            .I(N__47956));
    InMux I__11877 (
            .O(N__48021),
            .I(N__47953));
    InMux I__11876 (
            .O(N__48020),
            .I(N__47948));
    InMux I__11875 (
            .O(N__48017),
            .I(N__47948));
    Sp12to4 I__11874 (
            .O(N__48014),
            .I(N__47941));
    Span12Mux_h I__11873 (
            .O(N__48011),
            .I(N__47941));
    LocalMux I__11872 (
            .O(N__48008),
            .I(N__47941));
    LocalMux I__11871 (
            .O(N__48003),
            .I(N__47938));
    Span4Mux_v I__11870 (
            .O(N__47996),
            .I(N__47935));
    Span4Mux_h I__11869 (
            .O(N__47993),
            .I(N__47924));
    Span4Mux_s2_v I__11868 (
            .O(N__47990),
            .I(N__47924));
    Span4Mux_h I__11867 (
            .O(N__47987),
            .I(N__47924));
    Span4Mux_v I__11866 (
            .O(N__47978),
            .I(N__47924));
    Span4Mux_s2_v I__11865 (
            .O(N__47971),
            .I(N__47924));
    LocalMux I__11864 (
            .O(N__47968),
            .I(UART_TRANSMITTER_state_0));
    Odrv4 I__11863 (
            .O(N__47965),
            .I(UART_TRANSMITTER_state_0));
    Odrv4 I__11862 (
            .O(N__47962),
            .I(UART_TRANSMITTER_state_0));
    LocalMux I__11861 (
            .O(N__47959),
            .I(UART_TRANSMITTER_state_0));
    LocalMux I__11860 (
            .O(N__47956),
            .I(UART_TRANSMITTER_state_0));
    LocalMux I__11859 (
            .O(N__47953),
            .I(UART_TRANSMITTER_state_0));
    LocalMux I__11858 (
            .O(N__47948),
            .I(UART_TRANSMITTER_state_0));
    Odrv12 I__11857 (
            .O(N__47941),
            .I(UART_TRANSMITTER_state_0));
    Odrv12 I__11856 (
            .O(N__47938),
            .I(UART_TRANSMITTER_state_0));
    Odrv4 I__11855 (
            .O(N__47935),
            .I(UART_TRANSMITTER_state_0));
    Odrv4 I__11854 (
            .O(N__47924),
            .I(UART_TRANSMITTER_state_0));
    CascadeMux I__11853 (
            .O(N__47901),
            .I(N__47898));
    InMux I__11852 (
            .O(N__47898),
            .I(N__47895));
    LocalMux I__11851 (
            .O(N__47895),
            .I(N__47891));
    CascadeMux I__11850 (
            .O(N__47894),
            .I(N__47888));
    Span12Mux_s4_v I__11849 (
            .O(N__47891),
            .I(N__47885));
    InMux I__11848 (
            .O(N__47888),
            .I(N__47882));
    Odrv12 I__11847 (
            .O(N__47885),
            .I(rand_setpoint_25));
    LocalMux I__11846 (
            .O(N__47882),
            .I(rand_setpoint_25));
    InMux I__11845 (
            .O(N__47877),
            .I(N__47866));
    InMux I__11844 (
            .O(N__47876),
            .I(N__47866));
    InMux I__11843 (
            .O(N__47875),
            .I(N__47866));
    InMux I__11842 (
            .O(N__47874),
            .I(N__47861));
    InMux I__11841 (
            .O(N__47873),
            .I(N__47861));
    LocalMux I__11840 (
            .O(N__47866),
            .I(N__47858));
    LocalMux I__11839 (
            .O(N__47861),
            .I(N__47853));
    Span4Mux_h I__11838 (
            .O(N__47858),
            .I(N__47853));
    Span4Mux_h I__11837 (
            .O(N__47853),
            .I(N__47850));
    Odrv4 I__11836 (
            .O(N__47850),
            .I(data_out_5_1));
    CascadeMux I__11835 (
            .O(N__47847),
            .I(N__47843));
    InMux I__11834 (
            .O(N__47846),
            .I(N__47835));
    InMux I__11833 (
            .O(N__47843),
            .I(N__47822));
    InMux I__11832 (
            .O(N__47842),
            .I(N__47814));
    InMux I__11831 (
            .O(N__47841),
            .I(N__47806));
    InMux I__11830 (
            .O(N__47840),
            .I(N__47806));
    InMux I__11829 (
            .O(N__47839),
            .I(N__47797));
    InMux I__11828 (
            .O(N__47838),
            .I(N__47797));
    LocalMux I__11827 (
            .O(N__47835),
            .I(N__47788));
    InMux I__11826 (
            .O(N__47834),
            .I(N__47782));
    InMux I__11825 (
            .O(N__47833),
            .I(N__47782));
    InMux I__11824 (
            .O(N__47832),
            .I(N__47777));
    InMux I__11823 (
            .O(N__47831),
            .I(N__47777));
    InMux I__11822 (
            .O(N__47830),
            .I(N__47772));
    InMux I__11821 (
            .O(N__47829),
            .I(N__47772));
    InMux I__11820 (
            .O(N__47828),
            .I(N__47769));
    InMux I__11819 (
            .O(N__47827),
            .I(N__47764));
    InMux I__11818 (
            .O(N__47826),
            .I(N__47764));
    CascadeMux I__11817 (
            .O(N__47825),
            .I(N__47761));
    LocalMux I__11816 (
            .O(N__47822),
            .I(N__47758));
    InMux I__11815 (
            .O(N__47821),
            .I(N__47755));
    InMux I__11814 (
            .O(N__47820),
            .I(N__47752));
    InMux I__11813 (
            .O(N__47819),
            .I(N__47749));
    InMux I__11812 (
            .O(N__47818),
            .I(N__47744));
    InMux I__11811 (
            .O(N__47817),
            .I(N__47744));
    LocalMux I__11810 (
            .O(N__47814),
            .I(N__47741));
    InMux I__11809 (
            .O(N__47813),
            .I(N__47733));
    InMux I__11808 (
            .O(N__47812),
            .I(N__47733));
    InMux I__11807 (
            .O(N__47811),
            .I(N__47733));
    LocalMux I__11806 (
            .O(N__47806),
            .I(N__47730));
    InMux I__11805 (
            .O(N__47805),
            .I(N__47723));
    InMux I__11804 (
            .O(N__47804),
            .I(N__47723));
    InMux I__11803 (
            .O(N__47803),
            .I(N__47723));
    InMux I__11802 (
            .O(N__47802),
            .I(N__47720));
    LocalMux I__11801 (
            .O(N__47797),
            .I(N__47717));
    InMux I__11800 (
            .O(N__47796),
            .I(N__47714));
    InMux I__11799 (
            .O(N__47795),
            .I(N__47709));
    InMux I__11798 (
            .O(N__47794),
            .I(N__47709));
    InMux I__11797 (
            .O(N__47793),
            .I(N__47704));
    InMux I__11796 (
            .O(N__47792),
            .I(N__47704));
    InMux I__11795 (
            .O(N__47791),
            .I(N__47701));
    Span4Mux_h I__11794 (
            .O(N__47788),
            .I(N__47697));
    InMux I__11793 (
            .O(N__47787),
            .I(N__47694));
    LocalMux I__11792 (
            .O(N__47782),
            .I(N__47689));
    LocalMux I__11791 (
            .O(N__47777),
            .I(N__47689));
    LocalMux I__11790 (
            .O(N__47772),
            .I(N__47686));
    LocalMux I__11789 (
            .O(N__47769),
            .I(N__47681));
    LocalMux I__11788 (
            .O(N__47764),
            .I(N__47681));
    InMux I__11787 (
            .O(N__47761),
            .I(N__47678));
    Span4Mux_h I__11786 (
            .O(N__47758),
            .I(N__47662));
    LocalMux I__11785 (
            .O(N__47755),
            .I(N__47662));
    LocalMux I__11784 (
            .O(N__47752),
            .I(N__47662));
    LocalMux I__11783 (
            .O(N__47749),
            .I(N__47657));
    LocalMux I__11782 (
            .O(N__47744),
            .I(N__47657));
    Span4Mux_v I__11781 (
            .O(N__47741),
            .I(N__47654));
    InMux I__11780 (
            .O(N__47740),
            .I(N__47650));
    LocalMux I__11779 (
            .O(N__47733),
            .I(N__47637));
    Span4Mux_h I__11778 (
            .O(N__47730),
            .I(N__47637));
    LocalMux I__11777 (
            .O(N__47723),
            .I(N__47637));
    LocalMux I__11776 (
            .O(N__47720),
            .I(N__47637));
    Span4Mux_v I__11775 (
            .O(N__47717),
            .I(N__47637));
    LocalMux I__11774 (
            .O(N__47714),
            .I(N__47637));
    LocalMux I__11773 (
            .O(N__47709),
            .I(N__47630));
    LocalMux I__11772 (
            .O(N__47704),
            .I(N__47630));
    LocalMux I__11771 (
            .O(N__47701),
            .I(N__47630));
    InMux I__11770 (
            .O(N__47700),
            .I(N__47627));
    Span4Mux_v I__11769 (
            .O(N__47697),
            .I(N__47622));
    LocalMux I__11768 (
            .O(N__47694),
            .I(N__47622));
    Span4Mux_v I__11767 (
            .O(N__47689),
            .I(N__47613));
    Span4Mux_h I__11766 (
            .O(N__47686),
            .I(N__47613));
    Span4Mux_s2_v I__11765 (
            .O(N__47681),
            .I(N__47613));
    LocalMux I__11764 (
            .O(N__47678),
            .I(N__47613));
    InMux I__11763 (
            .O(N__47677),
            .I(N__47608));
    InMux I__11762 (
            .O(N__47676),
            .I(N__47608));
    InMux I__11761 (
            .O(N__47675),
            .I(N__47599));
    InMux I__11760 (
            .O(N__47674),
            .I(N__47599));
    InMux I__11759 (
            .O(N__47673),
            .I(N__47599));
    InMux I__11758 (
            .O(N__47672),
            .I(N__47599));
    InMux I__11757 (
            .O(N__47671),
            .I(N__47596));
    InMux I__11756 (
            .O(N__47670),
            .I(N__47591));
    InMux I__11755 (
            .O(N__47669),
            .I(N__47591));
    Span4Mux_v I__11754 (
            .O(N__47662),
            .I(N__47586));
    Span4Mux_s3_v I__11753 (
            .O(N__47657),
            .I(N__47586));
    Span4Mux_h I__11752 (
            .O(N__47654),
            .I(N__47583));
    InMux I__11751 (
            .O(N__47653),
            .I(N__47580));
    LocalMux I__11750 (
            .O(N__47650),
            .I(N__47575));
    Span4Mux_h I__11749 (
            .O(N__47637),
            .I(N__47575));
    Span4Mux_h I__11748 (
            .O(N__47630),
            .I(N__47566));
    LocalMux I__11747 (
            .O(N__47627),
            .I(N__47566));
    Span4Mux_v I__11746 (
            .O(N__47622),
            .I(N__47566));
    Span4Mux_h I__11745 (
            .O(N__47613),
            .I(N__47566));
    LocalMux I__11744 (
            .O(N__47608),
            .I(byte_transmit_counter_0));
    LocalMux I__11743 (
            .O(N__47599),
            .I(byte_transmit_counter_0));
    LocalMux I__11742 (
            .O(N__47596),
            .I(byte_transmit_counter_0));
    LocalMux I__11741 (
            .O(N__47591),
            .I(byte_transmit_counter_0));
    Odrv4 I__11740 (
            .O(N__47586),
            .I(byte_transmit_counter_0));
    Odrv4 I__11739 (
            .O(N__47583),
            .I(byte_transmit_counter_0));
    LocalMux I__11738 (
            .O(N__47580),
            .I(byte_transmit_counter_0));
    Odrv4 I__11737 (
            .O(N__47575),
            .I(byte_transmit_counter_0));
    Odrv4 I__11736 (
            .O(N__47566),
            .I(byte_transmit_counter_0));
    InMux I__11735 (
            .O(N__47547),
            .I(N__47543));
    InMux I__11734 (
            .O(N__47546),
            .I(N__47540));
    LocalMux I__11733 (
            .O(N__47543),
            .I(N__47537));
    LocalMux I__11732 (
            .O(N__47540),
            .I(N__47533));
    Span4Mux_h I__11731 (
            .O(N__47537),
            .I(N__47530));
    InMux I__11730 (
            .O(N__47536),
            .I(N__47527));
    Span4Mux_h I__11729 (
            .O(N__47533),
            .I(N__47524));
    Odrv4 I__11728 (
            .O(N__47530),
            .I(\c0.data_out_10_4 ));
    LocalMux I__11727 (
            .O(N__47527),
            .I(\c0.data_out_10_4 ));
    Odrv4 I__11726 (
            .O(N__47524),
            .I(\c0.data_out_10_4 ));
    CascadeMux I__11725 (
            .O(N__47517),
            .I(\c0.n8_adj_2198_cascade_ ));
    InMux I__11724 (
            .O(N__47514),
            .I(N__47510));
    InMux I__11723 (
            .O(N__47513),
            .I(N__47504));
    LocalMux I__11722 (
            .O(N__47510),
            .I(N__47501));
    InMux I__11721 (
            .O(N__47509),
            .I(N__47498));
    InMux I__11720 (
            .O(N__47508),
            .I(N__47489));
    InMux I__11719 (
            .O(N__47507),
            .I(N__47489));
    LocalMux I__11718 (
            .O(N__47504),
            .I(N__47478));
    Span4Mux_v I__11717 (
            .O(N__47501),
            .I(N__47473));
    LocalMux I__11716 (
            .O(N__47498),
            .I(N__47473));
    InMux I__11715 (
            .O(N__47497),
            .I(N__47470));
    InMux I__11714 (
            .O(N__47496),
            .I(N__47465));
    InMux I__11713 (
            .O(N__47495),
            .I(N__47465));
    InMux I__11712 (
            .O(N__47494),
            .I(N__47462));
    LocalMux I__11711 (
            .O(N__47489),
            .I(N__47459));
    InMux I__11710 (
            .O(N__47488),
            .I(N__47455));
    InMux I__11709 (
            .O(N__47487),
            .I(N__47451));
    InMux I__11708 (
            .O(N__47486),
            .I(N__47448));
    InMux I__11707 (
            .O(N__47485),
            .I(N__47445));
    InMux I__11706 (
            .O(N__47484),
            .I(N__47442));
    InMux I__11705 (
            .O(N__47483),
            .I(N__47439));
    InMux I__11704 (
            .O(N__47482),
            .I(N__47435));
    InMux I__11703 (
            .O(N__47481),
            .I(N__47432));
    Span4Mux_v I__11702 (
            .O(N__47478),
            .I(N__47428));
    Span4Mux_h I__11701 (
            .O(N__47473),
            .I(N__47423));
    LocalMux I__11700 (
            .O(N__47470),
            .I(N__47423));
    LocalMux I__11699 (
            .O(N__47465),
            .I(N__47416));
    LocalMux I__11698 (
            .O(N__47462),
            .I(N__47416));
    Span4Mux_s2_v I__11697 (
            .O(N__47459),
            .I(N__47416));
    InMux I__11696 (
            .O(N__47458),
            .I(N__47413));
    LocalMux I__11695 (
            .O(N__47455),
            .I(N__47410));
    InMux I__11694 (
            .O(N__47454),
            .I(N__47407));
    LocalMux I__11693 (
            .O(N__47451),
            .I(N__47404));
    LocalMux I__11692 (
            .O(N__47448),
            .I(N__47395));
    LocalMux I__11691 (
            .O(N__47445),
            .I(N__47395));
    LocalMux I__11690 (
            .O(N__47442),
            .I(N__47395));
    LocalMux I__11689 (
            .O(N__47439),
            .I(N__47395));
    InMux I__11688 (
            .O(N__47438),
            .I(N__47392));
    LocalMux I__11687 (
            .O(N__47435),
            .I(N__47387));
    LocalMux I__11686 (
            .O(N__47432),
            .I(N__47387));
    InMux I__11685 (
            .O(N__47431),
            .I(N__47384));
    Span4Mux_h I__11684 (
            .O(N__47428),
            .I(N__47379));
    Span4Mux_v I__11683 (
            .O(N__47423),
            .I(N__47379));
    Span4Mux_v I__11682 (
            .O(N__47416),
            .I(N__47376));
    LocalMux I__11681 (
            .O(N__47413),
            .I(N__47365));
    Span4Mux_v I__11680 (
            .O(N__47410),
            .I(N__47365));
    LocalMux I__11679 (
            .O(N__47407),
            .I(N__47365));
    Span4Mux_h I__11678 (
            .O(N__47404),
            .I(N__47365));
    Span4Mux_v I__11677 (
            .O(N__47395),
            .I(N__47365));
    LocalMux I__11676 (
            .O(N__47392),
            .I(byte_transmit_counter_1));
    Odrv12 I__11675 (
            .O(N__47387),
            .I(byte_transmit_counter_1));
    LocalMux I__11674 (
            .O(N__47384),
            .I(byte_transmit_counter_1));
    Odrv4 I__11673 (
            .O(N__47379),
            .I(byte_transmit_counter_1));
    Odrv4 I__11672 (
            .O(N__47376),
            .I(byte_transmit_counter_1));
    Odrv4 I__11671 (
            .O(N__47365),
            .I(byte_transmit_counter_1));
    CascadeMux I__11670 (
            .O(N__47352),
            .I(N__47349));
    InMux I__11669 (
            .O(N__47349),
            .I(N__47346));
    LocalMux I__11668 (
            .O(N__47346),
            .I(N__47343));
    Span12Mux_h I__11667 (
            .O(N__47343),
            .I(N__47340));
    Odrv12 I__11666 (
            .O(N__47340),
            .I(n10_adj_2430));
    InMux I__11665 (
            .O(N__47337),
            .I(N__47334));
    LocalMux I__11664 (
            .O(N__47334),
            .I(\c0.n17209 ));
    InMux I__11663 (
            .O(N__47331),
            .I(N__47328));
    LocalMux I__11662 (
            .O(N__47328),
            .I(\c0.n17297 ));
    CascadeMux I__11661 (
            .O(N__47325),
            .I(\c0.n17297_cascade_ ));
    InMux I__11660 (
            .O(N__47322),
            .I(N__47317));
    InMux I__11659 (
            .O(N__47321),
            .I(N__47314));
    InMux I__11658 (
            .O(N__47320),
            .I(N__47310));
    LocalMux I__11657 (
            .O(N__47317),
            .I(N__47307));
    LocalMux I__11656 (
            .O(N__47314),
            .I(N__47304));
    InMux I__11655 (
            .O(N__47313),
            .I(N__47301));
    LocalMux I__11654 (
            .O(N__47310),
            .I(N__47297));
    Span4Mux_h I__11653 (
            .O(N__47307),
            .I(N__47294));
    Span4Mux_h I__11652 (
            .O(N__47304),
            .I(N__47289));
    LocalMux I__11651 (
            .O(N__47301),
            .I(N__47289));
    InMux I__11650 (
            .O(N__47300),
            .I(N__47286));
    Odrv4 I__11649 (
            .O(N__47297),
            .I(\c0.data_out_7__2__N_447 ));
    Odrv4 I__11648 (
            .O(N__47294),
            .I(\c0.data_out_7__2__N_447 ));
    Odrv4 I__11647 (
            .O(N__47289),
            .I(\c0.data_out_7__2__N_447 ));
    LocalMux I__11646 (
            .O(N__47286),
            .I(\c0.data_out_7__2__N_447 ));
    InMux I__11645 (
            .O(N__47277),
            .I(N__47274));
    LocalMux I__11644 (
            .O(N__47274),
            .I(N__47271));
    Span4Mux_h I__11643 (
            .O(N__47271),
            .I(N__47268));
    Odrv4 I__11642 (
            .O(N__47268),
            .I(\c0.n14_adj_2176 ));
    InMux I__11641 (
            .O(N__47265),
            .I(N__47260));
    InMux I__11640 (
            .O(N__47264),
            .I(N__47257));
    InMux I__11639 (
            .O(N__47263),
            .I(N__47253));
    LocalMux I__11638 (
            .O(N__47260),
            .I(N__47250));
    LocalMux I__11637 (
            .O(N__47257),
            .I(N__47247));
    InMux I__11636 (
            .O(N__47256),
            .I(N__47244));
    LocalMux I__11635 (
            .O(N__47253),
            .I(N__47241));
    Span4Mux_v I__11634 (
            .O(N__47250),
            .I(N__47234));
    Span4Mux_h I__11633 (
            .O(N__47247),
            .I(N__47234));
    LocalMux I__11632 (
            .O(N__47244),
            .I(N__47234));
    Span4Mux_h I__11631 (
            .O(N__47241),
            .I(N__47231));
    Span4Mux_v I__11630 (
            .O(N__47234),
            .I(N__47227));
    Span4Mux_h I__11629 (
            .O(N__47231),
            .I(N__47224));
    InMux I__11628 (
            .O(N__47230),
            .I(N__47221));
    Span4Mux_s2_v I__11627 (
            .O(N__47227),
            .I(N__47218));
    Odrv4 I__11626 (
            .O(N__47224),
            .I(\c0.data_out_7_6 ));
    LocalMux I__11625 (
            .O(N__47221),
            .I(\c0.data_out_7_6 ));
    Odrv4 I__11624 (
            .O(N__47218),
            .I(\c0.data_out_7_6 ));
    CascadeMux I__11623 (
            .O(N__47211),
            .I(N__47208));
    InMux I__11622 (
            .O(N__47208),
            .I(N__47205));
    LocalMux I__11621 (
            .O(N__47205),
            .I(N__47202));
    Odrv4 I__11620 (
            .O(N__47202),
            .I(\c0.n12_adj_2180 ));
    CascadeMux I__11619 (
            .O(N__47199),
            .I(N__47196));
    InMux I__11618 (
            .O(N__47196),
            .I(N__47191));
    CascadeMux I__11617 (
            .O(N__47195),
            .I(N__47188));
    CascadeMux I__11616 (
            .O(N__47194),
            .I(N__47185));
    LocalMux I__11615 (
            .O(N__47191),
            .I(N__47182));
    InMux I__11614 (
            .O(N__47188),
            .I(N__47179));
    InMux I__11613 (
            .O(N__47185),
            .I(N__47176));
    Span4Mux_v I__11612 (
            .O(N__47182),
            .I(N__47173));
    LocalMux I__11611 (
            .O(N__47179),
            .I(N__47168));
    LocalMux I__11610 (
            .O(N__47176),
            .I(N__47168));
    Odrv4 I__11609 (
            .O(N__47173),
            .I(data_out_10_0));
    Odrv4 I__11608 (
            .O(N__47168),
            .I(data_out_10_0));
    InMux I__11607 (
            .O(N__47163),
            .I(N__47157));
    InMux I__11606 (
            .O(N__47162),
            .I(N__47157));
    LocalMux I__11605 (
            .O(N__47157),
            .I(N__47153));
    InMux I__11604 (
            .O(N__47156),
            .I(N__47150));
    Span12Mux_h I__11603 (
            .O(N__47153),
            .I(N__47147));
    LocalMux I__11602 (
            .O(N__47150),
            .I(N__47144));
    Span12Mux_h I__11601 (
            .O(N__47147),
            .I(N__47141));
    Span12Mux_v I__11600 (
            .O(N__47144),
            .I(N__47138));
    Odrv12 I__11599 (
            .O(N__47141),
            .I(\c0.data_out_7_3 ));
    Odrv12 I__11598 (
            .O(N__47138),
            .I(\c0.data_out_7_3 ));
    InMux I__11597 (
            .O(N__47133),
            .I(N__47128));
    InMux I__11596 (
            .O(N__47132),
            .I(N__47125));
    InMux I__11595 (
            .O(N__47131),
            .I(N__47121));
    LocalMux I__11594 (
            .O(N__47128),
            .I(N__47116));
    LocalMux I__11593 (
            .O(N__47125),
            .I(N__47113));
    InMux I__11592 (
            .O(N__47124),
            .I(N__47110));
    LocalMux I__11591 (
            .O(N__47121),
            .I(N__47107));
    InMux I__11590 (
            .O(N__47120),
            .I(N__47103));
    InMux I__11589 (
            .O(N__47119),
            .I(N__47100));
    Span4Mux_v I__11588 (
            .O(N__47116),
            .I(N__47097));
    Span4Mux_v I__11587 (
            .O(N__47113),
            .I(N__47092));
    LocalMux I__11586 (
            .O(N__47110),
            .I(N__47092));
    Span4Mux_v I__11585 (
            .O(N__47107),
            .I(N__47089));
    InMux I__11584 (
            .O(N__47106),
            .I(N__47086));
    LocalMux I__11583 (
            .O(N__47103),
            .I(N__47082));
    LocalMux I__11582 (
            .O(N__47100),
            .I(N__47075));
    Span4Mux_h I__11581 (
            .O(N__47097),
            .I(N__47075));
    Span4Mux_h I__11580 (
            .O(N__47092),
            .I(N__47075));
    Sp12to4 I__11579 (
            .O(N__47089),
            .I(N__47070));
    LocalMux I__11578 (
            .O(N__47086),
            .I(N__47070));
    InMux I__11577 (
            .O(N__47085),
            .I(N__47067));
    Odrv4 I__11576 (
            .O(N__47082),
            .I(\c0.data_out_5_3 ));
    Odrv4 I__11575 (
            .O(N__47075),
            .I(\c0.data_out_5_3 ));
    Odrv12 I__11574 (
            .O(N__47070),
            .I(\c0.data_out_5_3 ));
    LocalMux I__11573 (
            .O(N__47067),
            .I(\c0.data_out_5_3 ));
    InMux I__11572 (
            .O(N__47058),
            .I(N__47055));
    LocalMux I__11571 (
            .O(N__47055),
            .I(N__47052));
    Odrv4 I__11570 (
            .O(N__47052),
            .I(\c0.n17180 ));
    InMux I__11569 (
            .O(N__47049),
            .I(N__47045));
    InMux I__11568 (
            .O(N__47048),
            .I(N__47042));
    LocalMux I__11567 (
            .O(N__47045),
            .I(N__47039));
    LocalMux I__11566 (
            .O(N__47042),
            .I(N__47035));
    Span4Mux_h I__11565 (
            .O(N__47039),
            .I(N__47032));
    InMux I__11564 (
            .O(N__47038),
            .I(N__47029));
    Span4Mux_h I__11563 (
            .O(N__47035),
            .I(N__47026));
    Odrv4 I__11562 (
            .O(N__47032),
            .I(\c0.data_out_9_4 ));
    LocalMux I__11561 (
            .O(N__47029),
            .I(\c0.data_out_9_4 ));
    Odrv4 I__11560 (
            .O(N__47026),
            .I(\c0.data_out_9_4 ));
    CascadeMux I__11559 (
            .O(N__47019),
            .I(\c0.n17162_cascade_ ));
    InMux I__11558 (
            .O(N__47016),
            .I(N__47010));
    InMux I__11557 (
            .O(N__47015),
            .I(N__47007));
    InMux I__11556 (
            .O(N__47014),
            .I(N__47004));
    InMux I__11555 (
            .O(N__47013),
            .I(N__47001));
    LocalMux I__11554 (
            .O(N__47010),
            .I(N__46998));
    LocalMux I__11553 (
            .O(N__47007),
            .I(N__46994));
    LocalMux I__11552 (
            .O(N__47004),
            .I(N__46991));
    LocalMux I__11551 (
            .O(N__47001),
            .I(N__46986));
    Span4Mux_v I__11550 (
            .O(N__46998),
            .I(N__46986));
    InMux I__11549 (
            .O(N__46997),
            .I(N__46983));
    Span12Mux_v I__11548 (
            .O(N__46994),
            .I(N__46980));
    Span4Mux_v I__11547 (
            .O(N__46991),
            .I(N__46977));
    Span4Mux_h I__11546 (
            .O(N__46986),
            .I(N__46972));
    LocalMux I__11545 (
            .O(N__46983),
            .I(N__46972));
    Odrv12 I__11544 (
            .O(N__46980),
            .I(\c0.data_out_6_2 ));
    Odrv4 I__11543 (
            .O(N__46977),
            .I(\c0.data_out_6_2 ));
    Odrv4 I__11542 (
            .O(N__46972),
            .I(\c0.data_out_6_2 ));
    CascadeMux I__11541 (
            .O(N__46965),
            .I(N__46962));
    InMux I__11540 (
            .O(N__46962),
            .I(N__46959));
    LocalMux I__11539 (
            .O(N__46959),
            .I(N__46955));
    InMux I__11538 (
            .O(N__46958),
            .I(N__46952));
    Odrv4 I__11537 (
            .O(N__46955),
            .I(\c0.n17197 ));
    LocalMux I__11536 (
            .O(N__46952),
            .I(\c0.n17197 ));
    CascadeMux I__11535 (
            .O(N__46947),
            .I(\c0.n10_adj_2196_cascade_ ));
    InMux I__11534 (
            .O(N__46944),
            .I(N__46938));
    InMux I__11533 (
            .O(N__46943),
            .I(N__46938));
    LocalMux I__11532 (
            .O(N__46938),
            .I(\c0.n17261 ));
    CEMux I__11531 (
            .O(N__46935),
            .I(N__46930));
    CEMux I__11530 (
            .O(N__46934),
            .I(N__46927));
    CEMux I__11529 (
            .O(N__46933),
            .I(N__46924));
    LocalMux I__11528 (
            .O(N__46930),
            .I(N__46919));
    LocalMux I__11527 (
            .O(N__46927),
            .I(N__46915));
    LocalMux I__11526 (
            .O(N__46924),
            .I(N__46912));
    CEMux I__11525 (
            .O(N__46923),
            .I(N__46909));
    InMux I__11524 (
            .O(N__46922),
            .I(N__46906));
    Span4Mux_s3_h I__11523 (
            .O(N__46919),
            .I(N__46902));
    InMux I__11522 (
            .O(N__46918),
            .I(N__46899));
    Span4Mux_h I__11521 (
            .O(N__46915),
            .I(N__46895));
    Span4Mux_v I__11520 (
            .O(N__46912),
            .I(N__46890));
    LocalMux I__11519 (
            .O(N__46909),
            .I(N__46890));
    LocalMux I__11518 (
            .O(N__46906),
            .I(N__46887));
    InMux I__11517 (
            .O(N__46905),
            .I(N__46884));
    Span4Mux_h I__11516 (
            .O(N__46902),
            .I(N__46881));
    LocalMux I__11515 (
            .O(N__46899),
            .I(N__46878));
    InMux I__11514 (
            .O(N__46898),
            .I(N__46875));
    Span4Mux_v I__11513 (
            .O(N__46895),
            .I(N__46870));
    Span4Mux_h I__11512 (
            .O(N__46890),
            .I(N__46870));
    Span4Mux_v I__11511 (
            .O(N__46887),
            .I(N__46867));
    LocalMux I__11510 (
            .O(N__46884),
            .I(N__46864));
    Span4Mux_h I__11509 (
            .O(N__46881),
            .I(N__46859));
    Span4Mux_v I__11508 (
            .O(N__46878),
            .I(N__46859));
    LocalMux I__11507 (
            .O(N__46875),
            .I(N__46856));
    Span4Mux_h I__11506 (
            .O(N__46870),
            .I(N__46853));
    Span4Mux_h I__11505 (
            .O(N__46867),
            .I(N__46850));
    Span12Mux_h I__11504 (
            .O(N__46864),
            .I(N__46847));
    Span4Mux_h I__11503 (
            .O(N__46859),
            .I(N__46842));
    Span4Mux_v I__11502 (
            .O(N__46856),
            .I(N__46842));
    Odrv4 I__11501 (
            .O(N__46853),
            .I(\c0.n10595 ));
    Odrv4 I__11500 (
            .O(N__46850),
            .I(\c0.n10595 ));
    Odrv12 I__11499 (
            .O(N__46847),
            .I(\c0.n10595 ));
    Odrv4 I__11498 (
            .O(N__46842),
            .I(\c0.n10595 ));
    InMux I__11497 (
            .O(N__46833),
            .I(N__46829));
    CascadeMux I__11496 (
            .O(N__46832),
            .I(N__46826));
    LocalMux I__11495 (
            .O(N__46829),
            .I(N__46821));
    InMux I__11494 (
            .O(N__46826),
            .I(N__46818));
    InMux I__11493 (
            .O(N__46825),
            .I(N__46814));
    InMux I__11492 (
            .O(N__46824),
            .I(N__46811));
    Span4Mux_v I__11491 (
            .O(N__46821),
            .I(N__46806));
    LocalMux I__11490 (
            .O(N__46818),
            .I(N__46806));
    InMux I__11489 (
            .O(N__46817),
            .I(N__46803));
    LocalMux I__11488 (
            .O(N__46814),
            .I(N__46798));
    LocalMux I__11487 (
            .O(N__46811),
            .I(N__46798));
    Span4Mux_h I__11486 (
            .O(N__46806),
            .I(N__46795));
    LocalMux I__11485 (
            .O(N__46803),
            .I(\c0.data_out_6_0 ));
    Odrv12 I__11484 (
            .O(N__46798),
            .I(\c0.data_out_6_0 ));
    Odrv4 I__11483 (
            .O(N__46795),
            .I(\c0.data_out_6_0 ));
    InMux I__11482 (
            .O(N__46788),
            .I(N__46785));
    LocalMux I__11481 (
            .O(N__46785),
            .I(N__46781));
    InMux I__11480 (
            .O(N__46784),
            .I(N__46778));
    Odrv4 I__11479 (
            .O(N__46781),
            .I(\c0.n17129 ));
    LocalMux I__11478 (
            .O(N__46778),
            .I(\c0.n17129 ));
    CascadeMux I__11477 (
            .O(N__46773),
            .I(\c0.n10447_cascade_ ));
    InMux I__11476 (
            .O(N__46770),
            .I(N__46767));
    LocalMux I__11475 (
            .O(N__46767),
            .I(N__46763));
    InMux I__11474 (
            .O(N__46766),
            .I(N__46760));
    Span4Mux_v I__11473 (
            .O(N__46763),
            .I(N__46754));
    LocalMux I__11472 (
            .O(N__46760),
            .I(N__46754));
    InMux I__11471 (
            .O(N__46759),
            .I(N__46751));
    Span4Mux_h I__11470 (
            .O(N__46754),
            .I(N__46747));
    LocalMux I__11469 (
            .O(N__46751),
            .I(N__46744));
    InMux I__11468 (
            .O(N__46750),
            .I(N__46741));
    Odrv4 I__11467 (
            .O(N__46747),
            .I(\c0.data_out_6_1 ));
    Odrv4 I__11466 (
            .O(N__46744),
            .I(\c0.data_out_6_1 ));
    LocalMux I__11465 (
            .O(N__46741),
            .I(\c0.data_out_6_1 ));
    CascadeMux I__11464 (
            .O(N__46734),
            .I(N__46731));
    InMux I__11463 (
            .O(N__46731),
            .I(N__46728));
    LocalMux I__11462 (
            .O(N__46728),
            .I(N__46723));
    InMux I__11461 (
            .O(N__46727),
            .I(N__46720));
    InMux I__11460 (
            .O(N__46726),
            .I(N__46717));
    Span4Mux_h I__11459 (
            .O(N__46723),
            .I(N__46714));
    LocalMux I__11458 (
            .O(N__46720),
            .I(N__46711));
    LocalMux I__11457 (
            .O(N__46717),
            .I(\c0.n10183 ));
    Odrv4 I__11456 (
            .O(N__46714),
            .I(\c0.n10183 ));
    Odrv12 I__11455 (
            .O(N__46711),
            .I(\c0.n10183 ));
    InMux I__11454 (
            .O(N__46704),
            .I(N__46700));
    InMux I__11453 (
            .O(N__46703),
            .I(N__46697));
    LocalMux I__11452 (
            .O(N__46700),
            .I(N__46690));
    LocalMux I__11451 (
            .O(N__46697),
            .I(N__46690));
    InMux I__11450 (
            .O(N__46696),
            .I(N__46687));
    InMux I__11449 (
            .O(N__46695),
            .I(N__46684));
    Span4Mux_v I__11448 (
            .O(N__46690),
            .I(N__46681));
    LocalMux I__11447 (
            .O(N__46687),
            .I(N__46678));
    LocalMux I__11446 (
            .O(N__46684),
            .I(N__46675));
    Span4Mux_h I__11445 (
            .O(N__46681),
            .I(N__46670));
    Span4Mux_v I__11444 (
            .O(N__46678),
            .I(N__46670));
    Span4Mux_h I__11443 (
            .O(N__46675),
            .I(N__46667));
    Odrv4 I__11442 (
            .O(N__46670),
            .I(\c0.data_out_6_3 ));
    Odrv4 I__11441 (
            .O(N__46667),
            .I(\c0.data_out_6_3 ));
    CascadeMux I__11440 (
            .O(N__46662),
            .I(N__46659));
    InMux I__11439 (
            .O(N__46659),
            .I(N__46655));
    InMux I__11438 (
            .O(N__46658),
            .I(N__46652));
    LocalMux I__11437 (
            .O(N__46655),
            .I(\c0.n17222 ));
    LocalMux I__11436 (
            .O(N__46652),
            .I(\c0.n17222 ));
    CascadeMux I__11435 (
            .O(N__46647),
            .I(N__46643));
    CascadeMux I__11434 (
            .O(N__46646),
            .I(N__46640));
    InMux I__11433 (
            .O(N__46643),
            .I(N__46637));
    InMux I__11432 (
            .O(N__46640),
            .I(N__46634));
    LocalMux I__11431 (
            .O(N__46637),
            .I(N__46631));
    LocalMux I__11430 (
            .O(N__46634),
            .I(N__46628));
    Span4Mux_v I__11429 (
            .O(N__46631),
            .I(N__46623));
    Span4Mux_h I__11428 (
            .O(N__46628),
            .I(N__46620));
    InMux I__11427 (
            .O(N__46627),
            .I(N__46617));
    InMux I__11426 (
            .O(N__46626),
            .I(N__46614));
    Span4Mux_h I__11425 (
            .O(N__46623),
            .I(N__46611));
    Sp12to4 I__11424 (
            .O(N__46620),
            .I(N__46606));
    LocalMux I__11423 (
            .O(N__46617),
            .I(N__46606));
    LocalMux I__11422 (
            .O(N__46614),
            .I(\c0.data_out_9_7 ));
    Odrv4 I__11421 (
            .O(N__46611),
            .I(\c0.data_out_9_7 ));
    Odrv12 I__11420 (
            .O(N__46606),
            .I(\c0.data_out_9_7 ));
    CascadeMux I__11419 (
            .O(N__46599),
            .I(N__46596));
    InMux I__11418 (
            .O(N__46596),
            .I(N__46593));
    LocalMux I__11417 (
            .O(N__46593),
            .I(N__46590));
    Span4Mux_h I__11416 (
            .O(N__46590),
            .I(N__46586));
    InMux I__11415 (
            .O(N__46589),
            .I(N__46583));
    Odrv4 I__11414 (
            .O(N__46586),
            .I(\c0.n17243 ));
    LocalMux I__11413 (
            .O(N__46583),
            .I(\c0.n17243 ));
    InMux I__11412 (
            .O(N__46578),
            .I(N__46575));
    LocalMux I__11411 (
            .O(N__46575),
            .I(N__46571));
    InMux I__11410 (
            .O(N__46574),
            .I(N__46568));
    Span4Mux_h I__11409 (
            .O(N__46571),
            .I(N__46565));
    LocalMux I__11408 (
            .O(N__46568),
            .I(N__46562));
    Span4Mux_h I__11407 (
            .O(N__46565),
            .I(N__46559));
    Odrv12 I__11406 (
            .O(N__46562),
            .I(\c0.n17264 ));
    Odrv4 I__11405 (
            .O(N__46559),
            .I(\c0.n17264 ));
    CascadeMux I__11404 (
            .O(N__46554),
            .I(\c0.n10_adj_2191_cascade_ ));
    InMux I__11403 (
            .O(N__46551),
            .I(N__46548));
    LocalMux I__11402 (
            .O(N__46548),
            .I(N__46543));
    InMux I__11401 (
            .O(N__46547),
            .I(N__46540));
    InMux I__11400 (
            .O(N__46546),
            .I(N__46537));
    Odrv4 I__11399 (
            .O(N__46543),
            .I(\c0.tx.r_Clock_Count_7 ));
    LocalMux I__11398 (
            .O(N__46540),
            .I(\c0.tx.r_Clock_Count_7 ));
    LocalMux I__11397 (
            .O(N__46537),
            .I(\c0.tx.r_Clock_Count_7 ));
    InMux I__11396 (
            .O(N__46530),
            .I(N__46526));
    InMux I__11395 (
            .O(N__46529),
            .I(N__46523));
    LocalMux I__11394 (
            .O(N__46526),
            .I(data_out_3_7));
    LocalMux I__11393 (
            .O(N__46523),
            .I(data_out_3_7));
    InMux I__11392 (
            .O(N__46518),
            .I(N__46512));
    InMux I__11391 (
            .O(N__46517),
            .I(N__46512));
    LocalMux I__11390 (
            .O(N__46512),
            .I(data_out_2_7));
    InMux I__11389 (
            .O(N__46509),
            .I(N__46503));
    InMux I__11388 (
            .O(N__46508),
            .I(N__46500));
    InMux I__11387 (
            .O(N__46507),
            .I(N__46497));
    InMux I__11386 (
            .O(N__46506),
            .I(N__46494));
    LocalMux I__11385 (
            .O(N__46503),
            .I(N__46491));
    LocalMux I__11384 (
            .O(N__46500),
            .I(N__46488));
    LocalMux I__11383 (
            .O(N__46497),
            .I(N__46483));
    LocalMux I__11382 (
            .O(N__46494),
            .I(N__46483));
    Span4Mux_v I__11381 (
            .O(N__46491),
            .I(N__46480));
    Span4Mux_v I__11380 (
            .O(N__46488),
            .I(N__46477));
    Span12Mux_h I__11379 (
            .O(N__46483),
            .I(N__46473));
    Span4Mux_h I__11378 (
            .O(N__46480),
            .I(N__46470));
    Span4Mux_h I__11377 (
            .O(N__46477),
            .I(N__46467));
    InMux I__11376 (
            .O(N__46476),
            .I(N__46464));
    Span12Mux_h I__11375 (
            .O(N__46473),
            .I(N__46461));
    Sp12to4 I__11374 (
            .O(N__46470),
            .I(N__46456));
    Sp12to4 I__11373 (
            .O(N__46467),
            .I(N__46456));
    LocalMux I__11372 (
            .O(N__46464),
            .I(\c0.data_out_7__3__N_441 ));
    Odrv12 I__11371 (
            .O(N__46461),
            .I(\c0.data_out_7__3__N_441 ));
    Odrv12 I__11370 (
            .O(N__46456),
            .I(\c0.data_out_7__3__N_441 ));
    InMux I__11369 (
            .O(N__46449),
            .I(N__46446));
    LocalMux I__11368 (
            .O(N__46446),
            .I(N__46443));
    Span4Mux_v I__11367 (
            .O(N__46443),
            .I(N__46440));
    Odrv4 I__11366 (
            .O(N__46440),
            .I(\c0.n1 ));
    CascadeMux I__11365 (
            .O(N__46437),
            .I(\c0.n17747_cascade_ ));
    InMux I__11364 (
            .O(N__46434),
            .I(N__46431));
    LocalMux I__11363 (
            .O(N__46431),
            .I(\c0.n2_adj_2156 ));
    CascadeMux I__11362 (
            .O(N__46428),
            .I(\c0.n18220_cascade_ ));
    InMux I__11361 (
            .O(N__46425),
            .I(N__46422));
    LocalMux I__11360 (
            .O(N__46422),
            .I(N__46419));
    Odrv12 I__11359 (
            .O(N__46419),
            .I(\c0.n17607 ));
    InMux I__11358 (
            .O(N__46416),
            .I(N__46410));
    InMux I__11357 (
            .O(N__46415),
            .I(N__46407));
    InMux I__11356 (
            .O(N__46414),
            .I(N__46404));
    InMux I__11355 (
            .O(N__46413),
            .I(N__46397));
    LocalMux I__11354 (
            .O(N__46410),
            .I(N__46392));
    LocalMux I__11353 (
            .O(N__46407),
            .I(N__46392));
    LocalMux I__11352 (
            .O(N__46404),
            .I(N__46389));
    InMux I__11351 (
            .O(N__46403),
            .I(N__46386));
    InMux I__11350 (
            .O(N__46402),
            .I(N__46383));
    InMux I__11349 (
            .O(N__46401),
            .I(N__46380));
    InMux I__11348 (
            .O(N__46400),
            .I(N__46376));
    LocalMux I__11347 (
            .O(N__46397),
            .I(N__46372));
    Span4Mux_v I__11346 (
            .O(N__46392),
            .I(N__46369));
    Span4Mux_s2_v I__11345 (
            .O(N__46389),
            .I(N__46360));
    LocalMux I__11344 (
            .O(N__46386),
            .I(N__46360));
    LocalMux I__11343 (
            .O(N__46383),
            .I(N__46360));
    LocalMux I__11342 (
            .O(N__46380),
            .I(N__46360));
    InMux I__11341 (
            .O(N__46379),
            .I(N__46357));
    LocalMux I__11340 (
            .O(N__46376),
            .I(N__46354));
    InMux I__11339 (
            .O(N__46375),
            .I(N__46351));
    Span4Mux_v I__11338 (
            .O(N__46372),
            .I(N__46346));
    Span4Mux_h I__11337 (
            .O(N__46369),
            .I(N__46346));
    Span4Mux_v I__11336 (
            .O(N__46360),
            .I(N__46343));
    LocalMux I__11335 (
            .O(N__46357),
            .I(byte_transmit_counter_3));
    Odrv12 I__11334 (
            .O(N__46354),
            .I(byte_transmit_counter_3));
    LocalMux I__11333 (
            .O(N__46351),
            .I(byte_transmit_counter_3));
    Odrv4 I__11332 (
            .O(N__46346),
            .I(byte_transmit_counter_3));
    Odrv4 I__11331 (
            .O(N__46343),
            .I(byte_transmit_counter_3));
    InMux I__11330 (
            .O(N__46332),
            .I(N__46329));
    LocalMux I__11329 (
            .O(N__46329),
            .I(n10_adj_2413));
    CascadeMux I__11328 (
            .O(N__46326),
            .I(n18223_cascade_));
    InMux I__11327 (
            .O(N__46323),
            .I(N__46316));
    InMux I__11326 (
            .O(N__46322),
            .I(N__46316));
    InMux I__11325 (
            .O(N__46321),
            .I(N__46310));
    LocalMux I__11324 (
            .O(N__46316),
            .I(N__46307));
    InMux I__11323 (
            .O(N__46315),
            .I(N__46300));
    InMux I__11322 (
            .O(N__46314),
            .I(N__46300));
    InMux I__11321 (
            .O(N__46313),
            .I(N__46300));
    LocalMux I__11320 (
            .O(N__46310),
            .I(N__46285));
    Span4Mux_h I__11319 (
            .O(N__46307),
            .I(N__46280));
    LocalMux I__11318 (
            .O(N__46300),
            .I(N__46280));
    InMux I__11317 (
            .O(N__46299),
            .I(N__46277));
    InMux I__11316 (
            .O(N__46298),
            .I(N__46274));
    InMux I__11315 (
            .O(N__46297),
            .I(N__46267));
    InMux I__11314 (
            .O(N__46296),
            .I(N__46267));
    InMux I__11313 (
            .O(N__46295),
            .I(N__46267));
    InMux I__11312 (
            .O(N__46294),
            .I(N__46262));
    InMux I__11311 (
            .O(N__46293),
            .I(N__46262));
    InMux I__11310 (
            .O(N__46292),
            .I(N__46259));
    InMux I__11309 (
            .O(N__46291),
            .I(N__46256));
    InMux I__11308 (
            .O(N__46290),
            .I(N__46247));
    InMux I__11307 (
            .O(N__46289),
            .I(N__46244));
    InMux I__11306 (
            .O(N__46288),
            .I(N__46241));
    Span4Mux_s1_v I__11305 (
            .O(N__46285),
            .I(N__46234));
    Span4Mux_v I__11304 (
            .O(N__46280),
            .I(N__46234));
    LocalMux I__11303 (
            .O(N__46277),
            .I(N__46234));
    LocalMux I__11302 (
            .O(N__46274),
            .I(N__46227));
    LocalMux I__11301 (
            .O(N__46267),
            .I(N__46227));
    LocalMux I__11300 (
            .O(N__46262),
            .I(N__46227));
    LocalMux I__11299 (
            .O(N__46259),
            .I(N__46222));
    LocalMux I__11298 (
            .O(N__46256),
            .I(N__46222));
    InMux I__11297 (
            .O(N__46255),
            .I(N__46219));
    InMux I__11296 (
            .O(N__46254),
            .I(N__46216));
    InMux I__11295 (
            .O(N__46253),
            .I(N__46211));
    InMux I__11294 (
            .O(N__46252),
            .I(N__46211));
    InMux I__11293 (
            .O(N__46251),
            .I(N__46206));
    InMux I__11292 (
            .O(N__46250),
            .I(N__46206));
    LocalMux I__11291 (
            .O(N__46247),
            .I(N__46201));
    LocalMux I__11290 (
            .O(N__46244),
            .I(N__46201));
    LocalMux I__11289 (
            .O(N__46241),
            .I(N__46196));
    Span4Mux_h I__11288 (
            .O(N__46234),
            .I(N__46196));
    Span4Mux_v I__11287 (
            .O(N__46227),
            .I(N__46191));
    Span4Mux_s3_v I__11286 (
            .O(N__46222),
            .I(N__46191));
    LocalMux I__11285 (
            .O(N__46219),
            .I(byte_transmit_counter_2));
    LocalMux I__11284 (
            .O(N__46216),
            .I(byte_transmit_counter_2));
    LocalMux I__11283 (
            .O(N__46211),
            .I(byte_transmit_counter_2));
    LocalMux I__11282 (
            .O(N__46206),
            .I(byte_transmit_counter_2));
    Odrv4 I__11281 (
            .O(N__46201),
            .I(byte_transmit_counter_2));
    Odrv4 I__11280 (
            .O(N__46196),
            .I(byte_transmit_counter_2));
    Odrv4 I__11279 (
            .O(N__46191),
            .I(byte_transmit_counter_2));
    InMux I__11278 (
            .O(N__46176),
            .I(N__46173));
    LocalMux I__11277 (
            .O(N__46173),
            .I(N__46170));
    Span4Mux_h I__11276 (
            .O(N__46170),
            .I(N__46167));
    Odrv4 I__11275 (
            .O(N__46167),
            .I(n10));
    InMux I__11274 (
            .O(N__46164),
            .I(N__46161));
    LocalMux I__11273 (
            .O(N__46161),
            .I(N__46158));
    Odrv4 I__11272 (
            .O(N__46158),
            .I(n10960));
    InMux I__11271 (
            .O(N__46155),
            .I(N__46150));
    InMux I__11270 (
            .O(N__46154),
            .I(N__46147));
    InMux I__11269 (
            .O(N__46153),
            .I(N__46144));
    LocalMux I__11268 (
            .O(N__46150),
            .I(N__46137));
    LocalMux I__11267 (
            .O(N__46147),
            .I(N__46137));
    LocalMux I__11266 (
            .O(N__46144),
            .I(N__46137));
    Odrv4 I__11265 (
            .O(N__46137),
            .I(\c0.tx.r_Clock_Count_4 ));
    InMux I__11264 (
            .O(N__46134),
            .I(N__46131));
    LocalMux I__11263 (
            .O(N__46131),
            .I(N__46128));
    Odrv12 I__11262 (
            .O(N__46128),
            .I(n10994));
    InMux I__11261 (
            .O(N__46125),
            .I(N__46112));
    InMux I__11260 (
            .O(N__46124),
            .I(N__46112));
    InMux I__11259 (
            .O(N__46123),
            .I(N__46112));
    InMux I__11258 (
            .O(N__46122),
            .I(N__46106));
    InMux I__11257 (
            .O(N__46121),
            .I(N__46106));
    InMux I__11256 (
            .O(N__46120),
            .I(N__46101));
    InMux I__11255 (
            .O(N__46119),
            .I(N__46101));
    LocalMux I__11254 (
            .O(N__46112),
            .I(N__46098));
    InMux I__11253 (
            .O(N__46111),
            .I(N__46095));
    LocalMux I__11252 (
            .O(N__46106),
            .I(n5142));
    LocalMux I__11251 (
            .O(N__46101),
            .I(n5142));
    Odrv4 I__11250 (
            .O(N__46098),
            .I(n5142));
    LocalMux I__11249 (
            .O(N__46095),
            .I(n5142));
    InMux I__11248 (
            .O(N__46086),
            .I(N__46081));
    InMux I__11247 (
            .O(N__46085),
            .I(N__46078));
    InMux I__11246 (
            .O(N__46084),
            .I(N__46075));
    LocalMux I__11245 (
            .O(N__46081),
            .I(N__46070));
    LocalMux I__11244 (
            .O(N__46078),
            .I(N__46070));
    LocalMux I__11243 (
            .O(N__46075),
            .I(N__46067));
    Span4Mux_h I__11242 (
            .O(N__46070),
            .I(N__46062));
    Span4Mux_h I__11241 (
            .O(N__46067),
            .I(N__46062));
    Odrv4 I__11240 (
            .O(N__46062),
            .I(\c0.tx.r_Clock_Count_0 ));
    InMux I__11239 (
            .O(N__46059),
            .I(\c0.tx.n16120 ));
    InMux I__11238 (
            .O(N__46056),
            .I(N__46052));
    InMux I__11237 (
            .O(N__46055),
            .I(N__46048));
    LocalMux I__11236 (
            .O(N__46052),
            .I(N__46045));
    InMux I__11235 (
            .O(N__46051),
            .I(N__46042));
    LocalMux I__11234 (
            .O(N__46048),
            .I(\c0.tx.r_Clock_Count_5 ));
    Odrv4 I__11233 (
            .O(N__46045),
            .I(\c0.tx.r_Clock_Count_5 ));
    LocalMux I__11232 (
            .O(N__46042),
            .I(\c0.tx.r_Clock_Count_5 ));
    CascadeMux I__11231 (
            .O(N__46035),
            .I(N__46032));
    InMux I__11230 (
            .O(N__46032),
            .I(N__46029));
    LocalMux I__11229 (
            .O(N__46029),
            .I(n10963));
    InMux I__11228 (
            .O(N__46026),
            .I(\c0.tx.n16121 ));
    InMux I__11227 (
            .O(N__46023),
            .I(N__46018));
    InMux I__11226 (
            .O(N__46022),
            .I(N__46015));
    InMux I__11225 (
            .O(N__46021),
            .I(N__46012));
    LocalMux I__11224 (
            .O(N__46018),
            .I(\c0.tx.r_Clock_Count_6 ));
    LocalMux I__11223 (
            .O(N__46015),
            .I(\c0.tx.r_Clock_Count_6 ));
    LocalMux I__11222 (
            .O(N__46012),
            .I(\c0.tx.r_Clock_Count_6 ));
    InMux I__11221 (
            .O(N__46005),
            .I(N__46002));
    LocalMux I__11220 (
            .O(N__46002),
            .I(N__45999));
    Odrv4 I__11219 (
            .O(N__45999),
            .I(n10966));
    InMux I__11218 (
            .O(N__45996),
            .I(\c0.tx.n16122 ));
    InMux I__11217 (
            .O(N__45993),
            .I(\c0.tx.n16123 ));
    InMux I__11216 (
            .O(N__45990),
            .I(N__45987));
    LocalMux I__11215 (
            .O(N__45987),
            .I(N__45982));
    InMux I__11214 (
            .O(N__45986),
            .I(N__45979));
    InMux I__11213 (
            .O(N__45985),
            .I(N__45976));
    Span4Mux_h I__11212 (
            .O(N__45982),
            .I(N__45973));
    LocalMux I__11211 (
            .O(N__45979),
            .I(\c0.tx.r_Clock_Count_8 ));
    LocalMux I__11210 (
            .O(N__45976),
            .I(\c0.tx.r_Clock_Count_8 ));
    Odrv4 I__11209 (
            .O(N__45973),
            .I(\c0.tx.r_Clock_Count_8 ));
    CascadeMux I__11208 (
            .O(N__45966),
            .I(N__45955));
    CascadeMux I__11207 (
            .O(N__45965),
            .I(N__45952));
    CascadeMux I__11206 (
            .O(N__45964),
            .I(N__45949));
    CascadeMux I__11205 (
            .O(N__45963),
            .I(N__45946));
    CascadeMux I__11204 (
            .O(N__45962),
            .I(N__45942));
    CascadeMux I__11203 (
            .O(N__45961),
            .I(N__45937));
    CascadeMux I__11202 (
            .O(N__45960),
            .I(N__45934));
    CascadeMux I__11201 (
            .O(N__45959),
            .I(N__45931));
    CascadeMux I__11200 (
            .O(N__45958),
            .I(N__45928));
    InMux I__11199 (
            .O(N__45955),
            .I(N__45915));
    InMux I__11198 (
            .O(N__45952),
            .I(N__45915));
    InMux I__11197 (
            .O(N__45949),
            .I(N__45915));
    InMux I__11196 (
            .O(N__45946),
            .I(N__45915));
    InMux I__11195 (
            .O(N__45945),
            .I(N__45912));
    InMux I__11194 (
            .O(N__45942),
            .I(N__45909));
    InMux I__11193 (
            .O(N__45941),
            .I(N__45904));
    InMux I__11192 (
            .O(N__45940),
            .I(N__45904));
    InMux I__11191 (
            .O(N__45937),
            .I(N__45895));
    InMux I__11190 (
            .O(N__45934),
            .I(N__45895));
    InMux I__11189 (
            .O(N__45931),
            .I(N__45895));
    InMux I__11188 (
            .O(N__45928),
            .I(N__45895));
    InMux I__11187 (
            .O(N__45927),
            .I(N__45891));
    InMux I__11186 (
            .O(N__45926),
            .I(N__45884));
    InMux I__11185 (
            .O(N__45925),
            .I(N__45884));
    InMux I__11184 (
            .O(N__45924),
            .I(N__45884));
    LocalMux I__11183 (
            .O(N__45915),
            .I(N__45881));
    LocalMux I__11182 (
            .O(N__45912),
            .I(N__45872));
    LocalMux I__11181 (
            .O(N__45909),
            .I(N__45872));
    LocalMux I__11180 (
            .O(N__45904),
            .I(N__45872));
    LocalMux I__11179 (
            .O(N__45895),
            .I(N__45872));
    InMux I__11178 (
            .O(N__45894),
            .I(N__45869));
    LocalMux I__11177 (
            .O(N__45891),
            .I(N__45866));
    LocalMux I__11176 (
            .O(N__45884),
            .I(N__45859));
    Span4Mux_v I__11175 (
            .O(N__45881),
            .I(N__45859));
    Span4Mux_v I__11174 (
            .O(N__45872),
            .I(N__45859));
    LocalMux I__11173 (
            .O(N__45869),
            .I(\c0.tx.r_SM_Main_2 ));
    Odrv4 I__11172 (
            .O(N__45866),
            .I(\c0.tx.r_SM_Main_2 ));
    Odrv4 I__11171 (
            .O(N__45859),
            .I(\c0.tx.r_SM_Main_2 ));
    InMux I__11170 (
            .O(N__45852),
            .I(bfn_16_29_0_));
    InMux I__11169 (
            .O(N__45849),
            .I(N__45846));
    LocalMux I__11168 (
            .O(N__45846),
            .I(n10972));
    CascadeMux I__11167 (
            .O(N__45843),
            .I(N__45840));
    InMux I__11166 (
            .O(N__45840),
            .I(N__45833));
    InMux I__11165 (
            .O(N__45839),
            .I(N__45830));
    InMux I__11164 (
            .O(N__45838),
            .I(N__45827));
    CascadeMux I__11163 (
            .O(N__45837),
            .I(N__45824));
    InMux I__11162 (
            .O(N__45836),
            .I(N__45821));
    LocalMux I__11161 (
            .O(N__45833),
            .I(N__45818));
    LocalMux I__11160 (
            .O(N__45830),
            .I(N__45813));
    LocalMux I__11159 (
            .O(N__45827),
            .I(N__45813));
    InMux I__11158 (
            .O(N__45824),
            .I(N__45810));
    LocalMux I__11157 (
            .O(N__45821),
            .I(N__45807));
    Span4Mux_h I__11156 (
            .O(N__45818),
            .I(N__45802));
    Span4Mux_h I__11155 (
            .O(N__45813),
            .I(N__45802));
    LocalMux I__11154 (
            .O(N__45810),
            .I(N__45797));
    Span4Mux_h I__11153 (
            .O(N__45807),
            .I(N__45797));
    Odrv4 I__11152 (
            .O(N__45802),
            .I(data_out_8_7));
    Odrv4 I__11151 (
            .O(N__45797),
            .I(data_out_8_7));
    InMux I__11150 (
            .O(N__45792),
            .I(N__45789));
    LocalMux I__11149 (
            .O(N__45789),
            .I(n10951));
    InMux I__11148 (
            .O(N__45786),
            .I(N__45781));
    InMux I__11147 (
            .O(N__45785),
            .I(N__45778));
    InMux I__11146 (
            .O(N__45784),
            .I(N__45775));
    LocalMux I__11145 (
            .O(N__45781),
            .I(\c0.tx.r_Clock_Count_1 ));
    LocalMux I__11144 (
            .O(N__45778),
            .I(\c0.tx.r_Clock_Count_1 ));
    LocalMux I__11143 (
            .O(N__45775),
            .I(\c0.tx.r_Clock_Count_1 ));
    InMux I__11142 (
            .O(N__45768),
            .I(N__45765));
    LocalMux I__11141 (
            .O(N__45765),
            .I(N__45762));
    Odrv4 I__11140 (
            .O(N__45762),
            .I(n10969));
    InMux I__11139 (
            .O(N__45759),
            .I(N__45756));
    LocalMux I__11138 (
            .O(N__45756),
            .I(n32));
    CascadeMux I__11137 (
            .O(N__45753),
            .I(n29_cascade_));
    InMux I__11136 (
            .O(N__45750),
            .I(N__45747));
    LocalMux I__11135 (
            .O(N__45747),
            .I(n26));
    InMux I__11134 (
            .O(N__45744),
            .I(N__45740));
    InMux I__11133 (
            .O(N__45743),
            .I(N__45737));
    LocalMux I__11132 (
            .O(N__45740),
            .I(N__45734));
    LocalMux I__11131 (
            .O(N__45737),
            .I(N__45729));
    Span4Mux_h I__11130 (
            .O(N__45734),
            .I(N__45724));
    InMux I__11129 (
            .O(N__45733),
            .I(N__45719));
    InMux I__11128 (
            .O(N__45732),
            .I(N__45719));
    Span12Mux_h I__11127 (
            .O(N__45729),
            .I(N__45716));
    InMux I__11126 (
            .O(N__45728),
            .I(N__45711));
    InMux I__11125 (
            .O(N__45727),
            .I(N__45711));
    Span4Mux_h I__11124 (
            .O(N__45724),
            .I(N__45708));
    LocalMux I__11123 (
            .O(N__45719),
            .I(N__45705));
    Odrv12 I__11122 (
            .O(N__45716),
            .I(\c0.data_out_5_2 ));
    LocalMux I__11121 (
            .O(N__45711),
            .I(\c0.data_out_5_2 ));
    Odrv4 I__11120 (
            .O(N__45708),
            .I(\c0.data_out_5_2 ));
    Odrv4 I__11119 (
            .O(N__45705),
            .I(\c0.data_out_5_2 ));
    CascadeMux I__11118 (
            .O(N__45696),
            .I(N__45693));
    InMux I__11117 (
            .O(N__45693),
            .I(N__45690));
    LocalMux I__11116 (
            .O(N__45690),
            .I(N__45687));
    Span4Mux_h I__11115 (
            .O(N__45687),
            .I(N__45684));
    Odrv4 I__11114 (
            .O(N__45684),
            .I(\c0.n10196 ));
    CascadeMux I__11113 (
            .O(N__45681),
            .I(\c0.n10196_cascade_ ));
    InMux I__11112 (
            .O(N__45678),
            .I(N__45675));
    LocalMux I__11111 (
            .O(N__45675),
            .I(N__45672));
    Span4Mux_v I__11110 (
            .O(N__45672),
            .I(N__45667));
    InMux I__11109 (
            .O(N__45671),
            .I(N__45662));
    InMux I__11108 (
            .O(N__45670),
            .I(N__45662));
    Odrv4 I__11107 (
            .O(N__45667),
            .I(\c0.data_out_10_3 ));
    LocalMux I__11106 (
            .O(N__45662),
            .I(\c0.data_out_10_3 ));
    InMux I__11105 (
            .O(N__45657),
            .I(N__45653));
    InMux I__11104 (
            .O(N__45656),
            .I(N__45650));
    LocalMux I__11103 (
            .O(N__45653),
            .I(N__45647));
    LocalMux I__11102 (
            .O(N__45650),
            .I(N__45643));
    Span4Mux_h I__11101 (
            .O(N__45647),
            .I(N__45640));
    InMux I__11100 (
            .O(N__45646),
            .I(N__45637));
    Span4Mux_h I__11099 (
            .O(N__45643),
            .I(N__45634));
    Span4Mux_v I__11098 (
            .O(N__45640),
            .I(N__45631));
    LocalMux I__11097 (
            .O(N__45637),
            .I(N__45626));
    Span4Mux_h I__11096 (
            .O(N__45634),
            .I(N__45626));
    Odrv4 I__11095 (
            .O(N__45631),
            .I(\c0.data_out_6_4 ));
    Odrv4 I__11094 (
            .O(N__45626),
            .I(\c0.data_out_6_4 ));
    InMux I__11093 (
            .O(N__45621),
            .I(N__45617));
    InMux I__11092 (
            .O(N__45620),
            .I(N__45611));
    LocalMux I__11091 (
            .O(N__45617),
            .I(N__45608));
    InMux I__11090 (
            .O(N__45616),
            .I(N__45605));
    InMux I__11089 (
            .O(N__45615),
            .I(N__45600));
    InMux I__11088 (
            .O(N__45614),
            .I(N__45600));
    LocalMux I__11087 (
            .O(N__45611),
            .I(data_out_8_5));
    Odrv4 I__11086 (
            .O(N__45608),
            .I(data_out_8_5));
    LocalMux I__11085 (
            .O(N__45605),
            .I(data_out_8_5));
    LocalMux I__11084 (
            .O(N__45600),
            .I(data_out_8_5));
    InMux I__11083 (
            .O(N__45591),
            .I(N__45587));
    InMux I__11082 (
            .O(N__45590),
            .I(N__45584));
    LocalMux I__11081 (
            .O(N__45587),
            .I(N__45579));
    LocalMux I__11080 (
            .O(N__45584),
            .I(N__45579));
    Odrv12 I__11079 (
            .O(N__45579),
            .I(\c0.n10392 ));
    InMux I__11078 (
            .O(N__45576),
            .I(bfn_16_28_0_));
    InMux I__11077 (
            .O(N__45573),
            .I(\c0.tx.n16117 ));
    InMux I__11076 (
            .O(N__45570),
            .I(N__45565));
    InMux I__11075 (
            .O(N__45569),
            .I(N__45562));
    InMux I__11074 (
            .O(N__45568),
            .I(N__45559));
    LocalMux I__11073 (
            .O(N__45565),
            .I(\c0.tx.r_Clock_Count_2 ));
    LocalMux I__11072 (
            .O(N__45562),
            .I(\c0.tx.r_Clock_Count_2 ));
    LocalMux I__11071 (
            .O(N__45559),
            .I(\c0.tx.r_Clock_Count_2 ));
    InMux I__11070 (
            .O(N__45552),
            .I(N__45549));
    LocalMux I__11069 (
            .O(N__45549),
            .I(n10954));
    InMux I__11068 (
            .O(N__45546),
            .I(\c0.tx.n16118 ));
    CascadeMux I__11067 (
            .O(N__45543),
            .I(N__45538));
    InMux I__11066 (
            .O(N__45542),
            .I(N__45535));
    InMux I__11065 (
            .O(N__45541),
            .I(N__45532));
    InMux I__11064 (
            .O(N__45538),
            .I(N__45529));
    LocalMux I__11063 (
            .O(N__45535),
            .I(\c0.tx.r_Clock_Count_3 ));
    LocalMux I__11062 (
            .O(N__45532),
            .I(\c0.tx.r_Clock_Count_3 ));
    LocalMux I__11061 (
            .O(N__45529),
            .I(\c0.tx.r_Clock_Count_3 ));
    InMux I__11060 (
            .O(N__45522),
            .I(N__45519));
    LocalMux I__11059 (
            .O(N__45519),
            .I(n10957));
    InMux I__11058 (
            .O(N__45516),
            .I(\c0.tx.n16119 ));
    CascadeMux I__11057 (
            .O(N__45513),
            .I(N__45510));
    InMux I__11056 (
            .O(N__45510),
            .I(N__45506));
    InMux I__11055 (
            .O(N__45509),
            .I(N__45503));
    LocalMux I__11054 (
            .O(N__45506),
            .I(N__45500));
    LocalMux I__11053 (
            .O(N__45503),
            .I(\c0.n10179 ));
    Odrv12 I__11052 (
            .O(N__45500),
            .I(\c0.n10179 ));
    InMux I__11051 (
            .O(N__45495),
            .I(N__45491));
    InMux I__11050 (
            .O(N__45494),
            .I(N__45488));
    LocalMux I__11049 (
            .O(N__45491),
            .I(N__45485));
    LocalMux I__11048 (
            .O(N__45488),
            .I(N__45482));
    Span4Mux_h I__11047 (
            .O(N__45485),
            .I(N__45479));
    Span4Mux_h I__11046 (
            .O(N__45482),
            .I(N__45476));
    Span4Mux_h I__11045 (
            .O(N__45479),
            .I(N__45473));
    Odrv4 I__11044 (
            .O(N__45476),
            .I(\c0.n10188 ));
    Odrv4 I__11043 (
            .O(N__45473),
            .I(\c0.n10188 ));
    CascadeMux I__11042 (
            .O(N__45468),
            .I(\c0.n17209_cascade_ ));
    InMux I__11041 (
            .O(N__45465),
            .I(N__45460));
    CascadeMux I__11040 (
            .O(N__45464),
            .I(N__45457));
    InMux I__11039 (
            .O(N__45463),
            .I(N__45454));
    LocalMux I__11038 (
            .O(N__45460),
            .I(N__45451));
    InMux I__11037 (
            .O(N__45457),
            .I(N__45448));
    LocalMux I__11036 (
            .O(N__45454),
            .I(\c0.data_out_10_2 ));
    Odrv12 I__11035 (
            .O(N__45451),
            .I(\c0.data_out_10_2 ));
    LocalMux I__11034 (
            .O(N__45448),
            .I(\c0.data_out_10_2 ));
    InMux I__11033 (
            .O(N__45441),
            .I(N__45438));
    LocalMux I__11032 (
            .O(N__45438),
            .I(\c0.n6_adj_2216 ));
    InMux I__11031 (
            .O(N__45435),
            .I(N__45430));
    InMux I__11030 (
            .O(N__45434),
            .I(N__45425));
    InMux I__11029 (
            .O(N__45433),
            .I(N__45425));
    LocalMux I__11028 (
            .O(N__45430),
            .I(\c0.data_out_9_6 ));
    LocalMux I__11027 (
            .O(N__45425),
            .I(\c0.data_out_9_6 ));
    InMux I__11026 (
            .O(N__45420),
            .I(N__45417));
    LocalMux I__11025 (
            .O(N__45417),
            .I(\c0.n17200 ));
    InMux I__11024 (
            .O(N__45414),
            .I(N__45410));
    InMux I__11023 (
            .O(N__45413),
            .I(N__45407));
    LocalMux I__11022 (
            .O(N__45410),
            .I(N__45402));
    LocalMux I__11021 (
            .O(N__45407),
            .I(N__45399));
    InMux I__11020 (
            .O(N__45406),
            .I(N__45393));
    InMux I__11019 (
            .O(N__45405),
            .I(N__45393));
    Span4Mux_h I__11018 (
            .O(N__45402),
            .I(N__45388));
    Span4Mux_v I__11017 (
            .O(N__45399),
            .I(N__45388));
    InMux I__11016 (
            .O(N__45398),
            .I(N__45385));
    LocalMux I__11015 (
            .O(N__45393),
            .I(\c0.data_out_8_0 ));
    Odrv4 I__11014 (
            .O(N__45388),
            .I(\c0.data_out_8_0 ));
    LocalMux I__11013 (
            .O(N__45385),
            .I(\c0.data_out_8_0 ));
    InMux I__11012 (
            .O(N__45378),
            .I(N__45375));
    LocalMux I__11011 (
            .O(N__45375),
            .I(n8_adj_2445));
    InMux I__11010 (
            .O(N__45372),
            .I(N__45369));
    LocalMux I__11009 (
            .O(N__45369),
            .I(n6_adj_2446));
    InMux I__11008 (
            .O(N__45366),
            .I(N__45363));
    LocalMux I__11007 (
            .O(N__45363),
            .I(N__45360));
    Span4Mux_h I__11006 (
            .O(N__45360),
            .I(N__45357));
    Odrv4 I__11005 (
            .O(N__45357),
            .I(n23));
    InMux I__11004 (
            .O(N__45354),
            .I(N__45351));
    LocalMux I__11003 (
            .O(N__45351),
            .I(N__45348));
    Span4Mux_s1_v I__11002 (
            .O(N__45348),
            .I(N__45345));
    Span4Mux_h I__11001 (
            .O(N__45345),
            .I(N__45342));
    Odrv4 I__11000 (
            .O(N__45342),
            .I(\c0.n17622 ));
    InMux I__10999 (
            .O(N__45339),
            .I(N__45336));
    LocalMux I__10998 (
            .O(N__45336),
            .I(\c0.n18088 ));
    CascadeMux I__10997 (
            .O(N__45333),
            .I(\c0.n2_adj_2164_cascade_ ));
    InMux I__10996 (
            .O(N__45330),
            .I(N__45327));
    LocalMux I__10995 (
            .O(N__45327),
            .I(n18091));
    InMux I__10994 (
            .O(N__45324),
            .I(N__45318));
    InMux I__10993 (
            .O(N__45323),
            .I(N__45318));
    LocalMux I__10992 (
            .O(N__45318),
            .I(data_out_3_5));
    InMux I__10991 (
            .O(N__45315),
            .I(N__45312));
    LocalMux I__10990 (
            .O(N__45312),
            .I(N__45309));
    Sp12to4 I__10989 (
            .O(N__45309),
            .I(N__45305));
    InMux I__10988 (
            .O(N__45308),
            .I(N__45302));
    Span12Mux_v I__10987 (
            .O(N__45305),
            .I(N__45299));
    LocalMux I__10986 (
            .O(N__45302),
            .I(\c0.data_out_0_6 ));
    Odrv12 I__10985 (
            .O(N__45299),
            .I(\c0.data_out_0_6 ));
    CascadeMux I__10984 (
            .O(N__45294),
            .I(N__45290));
    InMux I__10983 (
            .O(N__45293),
            .I(N__45287));
    InMux I__10982 (
            .O(N__45290),
            .I(N__45284));
    LocalMux I__10981 (
            .O(N__45287),
            .I(N__45281));
    LocalMux I__10980 (
            .O(N__45284),
            .I(N__45278));
    Span4Mux_v I__10979 (
            .O(N__45281),
            .I(N__45275));
    Span4Mux_v I__10978 (
            .O(N__45278),
            .I(N__45272));
    Odrv4 I__10977 (
            .O(N__45275),
            .I(n4));
    Odrv4 I__10976 (
            .O(N__45272),
            .I(n4));
    InMux I__10975 (
            .O(N__45267),
            .I(N__45264));
    LocalMux I__10974 (
            .O(N__45264),
            .I(N__45255));
    InMux I__10973 (
            .O(N__45263),
            .I(N__45252));
    InMux I__10972 (
            .O(N__45262),
            .I(N__45247));
    InMux I__10971 (
            .O(N__45261),
            .I(N__45247));
    InMux I__10970 (
            .O(N__45260),
            .I(N__45244));
    InMux I__10969 (
            .O(N__45259),
            .I(N__45241));
    InMux I__10968 (
            .O(N__45258),
            .I(N__45238));
    Span4Mux_s1_v I__10967 (
            .O(N__45255),
            .I(N__45235));
    LocalMux I__10966 (
            .O(N__45252),
            .I(N__45230));
    LocalMux I__10965 (
            .O(N__45247),
            .I(N__45230));
    LocalMux I__10964 (
            .O(N__45244),
            .I(N__45227));
    LocalMux I__10963 (
            .O(N__45241),
            .I(N__45224));
    LocalMux I__10962 (
            .O(N__45238),
            .I(N__45221));
    Sp12to4 I__10961 (
            .O(N__45235),
            .I(N__45211));
    Span12Mux_s2_v I__10960 (
            .O(N__45230),
            .I(N__45211));
    Span4Mux_h I__10959 (
            .O(N__45227),
            .I(N__45208));
    Span4Mux_v I__10958 (
            .O(N__45224),
            .I(N__45203));
    Span4Mux_v I__10957 (
            .O(N__45221),
            .I(N__45203));
    InMux I__10956 (
            .O(N__45220),
            .I(N__45200));
    InMux I__10955 (
            .O(N__45219),
            .I(N__45191));
    InMux I__10954 (
            .O(N__45218),
            .I(N__45191));
    InMux I__10953 (
            .O(N__45217),
            .I(N__45191));
    InMux I__10952 (
            .O(N__45216),
            .I(N__45191));
    Span12Mux_v I__10951 (
            .O(N__45211),
            .I(N__45188));
    Odrv4 I__10950 (
            .O(N__45208),
            .I(r_Rx_Data));
    Odrv4 I__10949 (
            .O(N__45203),
            .I(r_Rx_Data));
    LocalMux I__10948 (
            .O(N__45200),
            .I(r_Rx_Data));
    LocalMux I__10947 (
            .O(N__45191),
            .I(r_Rx_Data));
    Odrv12 I__10946 (
            .O(N__45188),
            .I(r_Rx_Data));
    InMux I__10945 (
            .O(N__45177),
            .I(N__45172));
    InMux I__10944 (
            .O(N__45176),
            .I(N__45169));
    InMux I__10943 (
            .O(N__45175),
            .I(N__45166));
    LocalMux I__10942 (
            .O(N__45172),
            .I(N__45163));
    LocalMux I__10941 (
            .O(N__45169),
            .I(N__45160));
    LocalMux I__10940 (
            .O(N__45166),
            .I(N__45157));
    Span4Mux_v I__10939 (
            .O(N__45163),
            .I(N__45153));
    Span4Mux_h I__10938 (
            .O(N__45160),
            .I(N__45150));
    Span4Mux_v I__10937 (
            .O(N__45157),
            .I(N__45147));
    InMux I__10936 (
            .O(N__45156),
            .I(N__45144));
    Odrv4 I__10935 (
            .O(N__45153),
            .I(n9999));
    Odrv4 I__10934 (
            .O(N__45150),
            .I(n9999));
    Odrv4 I__10933 (
            .O(N__45147),
            .I(n9999));
    LocalMux I__10932 (
            .O(N__45144),
            .I(n9999));
    InMux I__10931 (
            .O(N__45135),
            .I(N__45127));
    InMux I__10930 (
            .O(N__45134),
            .I(N__45124));
    CascadeMux I__10929 (
            .O(N__45133),
            .I(N__45121));
    InMux I__10928 (
            .O(N__45132),
            .I(N__45113));
    InMux I__10927 (
            .O(N__45131),
            .I(N__45113));
    InMux I__10926 (
            .O(N__45130),
            .I(N__45113));
    LocalMux I__10925 (
            .O(N__45127),
            .I(N__45110));
    LocalMux I__10924 (
            .O(N__45124),
            .I(N__45107));
    InMux I__10923 (
            .O(N__45121),
            .I(N__45104));
    InMux I__10922 (
            .O(N__45120),
            .I(N__45101));
    LocalMux I__10921 (
            .O(N__45113),
            .I(N__45098));
    Span4Mux_h I__10920 (
            .O(N__45110),
            .I(N__45094));
    Span4Mux_v I__10919 (
            .O(N__45107),
            .I(N__45089));
    LocalMux I__10918 (
            .O(N__45104),
            .I(N__45089));
    LocalMux I__10917 (
            .O(N__45101),
            .I(N__45086));
    Span4Mux_h I__10916 (
            .O(N__45098),
            .I(N__45083));
    CascadeMux I__10915 (
            .O(N__45097),
            .I(N__45080));
    Span4Mux_h I__10914 (
            .O(N__45094),
            .I(N__45077));
    Span4Mux_h I__10913 (
            .O(N__45089),
            .I(N__45074));
    Span12Mux_h I__10912 (
            .O(N__45086),
            .I(N__45071));
    Span4Mux_h I__10911 (
            .O(N__45083),
            .I(N__45068));
    InMux I__10910 (
            .O(N__45080),
            .I(N__45065));
    Odrv4 I__10909 (
            .O(N__45077),
            .I(rx_data_4));
    Odrv4 I__10908 (
            .O(N__45074),
            .I(rx_data_4));
    Odrv12 I__10907 (
            .O(N__45071),
            .I(rx_data_4));
    Odrv4 I__10906 (
            .O(N__45068),
            .I(rx_data_4));
    LocalMux I__10905 (
            .O(N__45065),
            .I(rx_data_4));
    InMux I__10904 (
            .O(N__45054),
            .I(N__45051));
    LocalMux I__10903 (
            .O(N__45051),
            .I(N__45047));
    InMux I__10902 (
            .O(N__45050),
            .I(N__45044));
    Span4Mux_h I__10901 (
            .O(N__45047),
            .I(N__45041));
    LocalMux I__10900 (
            .O(N__45044),
            .I(data_out_1_6));
    Odrv4 I__10899 (
            .O(N__45041),
            .I(data_out_1_6));
    InMux I__10898 (
            .O(N__45036),
            .I(N__45033));
    LocalMux I__10897 (
            .O(N__45033),
            .I(N__45025));
    InMux I__10896 (
            .O(N__45032),
            .I(N__45022));
    InMux I__10895 (
            .O(N__45031),
            .I(N__45014));
    InMux I__10894 (
            .O(N__45030),
            .I(N__45011));
    InMux I__10893 (
            .O(N__45029),
            .I(N__45008));
    InMux I__10892 (
            .O(N__45028),
            .I(N__45005));
    Span4Mux_s2_v I__10891 (
            .O(N__45025),
            .I(N__45002));
    LocalMux I__10890 (
            .O(N__45022),
            .I(N__44999));
    InMux I__10889 (
            .O(N__45021),
            .I(N__44996));
    InMux I__10888 (
            .O(N__45020),
            .I(N__44993));
    InMux I__10887 (
            .O(N__45019),
            .I(N__44987));
    InMux I__10886 (
            .O(N__45018),
            .I(N__44983));
    CascadeMux I__10885 (
            .O(N__45017),
            .I(N__44979));
    LocalMux I__10884 (
            .O(N__45014),
            .I(N__44972));
    LocalMux I__10883 (
            .O(N__45011),
            .I(N__44967));
    LocalMux I__10882 (
            .O(N__45008),
            .I(N__44967));
    LocalMux I__10881 (
            .O(N__45005),
            .I(N__44964));
    Span4Mux_h I__10880 (
            .O(N__45002),
            .I(N__44955));
    Span4Mux_s2_v I__10879 (
            .O(N__44999),
            .I(N__44955));
    LocalMux I__10878 (
            .O(N__44996),
            .I(N__44955));
    LocalMux I__10877 (
            .O(N__44993),
            .I(N__44955));
    InMux I__10876 (
            .O(N__44992),
            .I(N__44952));
    InMux I__10875 (
            .O(N__44991),
            .I(N__44949));
    InMux I__10874 (
            .O(N__44990),
            .I(N__44946));
    LocalMux I__10873 (
            .O(N__44987),
            .I(N__44942));
    InMux I__10872 (
            .O(N__44986),
            .I(N__44939));
    LocalMux I__10871 (
            .O(N__44983),
            .I(N__44936));
    InMux I__10870 (
            .O(N__44982),
            .I(N__44933));
    InMux I__10869 (
            .O(N__44979),
            .I(N__44928));
    InMux I__10868 (
            .O(N__44978),
            .I(N__44925));
    InMux I__10867 (
            .O(N__44977),
            .I(N__44922));
    InMux I__10866 (
            .O(N__44976),
            .I(N__44919));
    InMux I__10865 (
            .O(N__44975),
            .I(N__44916));
    Span4Mux_v I__10864 (
            .O(N__44972),
            .I(N__44912));
    Span4Mux_v I__10863 (
            .O(N__44967),
            .I(N__44907));
    Span4Mux_v I__10862 (
            .O(N__44964),
            .I(N__44907));
    Span4Mux_v I__10861 (
            .O(N__44955),
            .I(N__44898));
    LocalMux I__10860 (
            .O(N__44952),
            .I(N__44898));
    LocalMux I__10859 (
            .O(N__44949),
            .I(N__44898));
    LocalMux I__10858 (
            .O(N__44946),
            .I(N__44898));
    InMux I__10857 (
            .O(N__44945),
            .I(N__44895));
    Span4Mux_v I__10856 (
            .O(N__44942),
            .I(N__44892));
    LocalMux I__10855 (
            .O(N__44939),
            .I(N__44889));
    Span4Mux_h I__10854 (
            .O(N__44936),
            .I(N__44884));
    LocalMux I__10853 (
            .O(N__44933),
            .I(N__44884));
    InMux I__10852 (
            .O(N__44932),
            .I(N__44881));
    InMux I__10851 (
            .O(N__44931),
            .I(N__44878));
    LocalMux I__10850 (
            .O(N__44928),
            .I(N__44871));
    LocalMux I__10849 (
            .O(N__44925),
            .I(N__44871));
    LocalMux I__10848 (
            .O(N__44922),
            .I(N__44871));
    LocalMux I__10847 (
            .O(N__44919),
            .I(N__44866));
    LocalMux I__10846 (
            .O(N__44916),
            .I(N__44866));
    InMux I__10845 (
            .O(N__44915),
            .I(N__44863));
    Span4Mux_h I__10844 (
            .O(N__44912),
            .I(N__44859));
    Span4Mux_h I__10843 (
            .O(N__44907),
            .I(N__44854));
    Span4Mux_v I__10842 (
            .O(N__44898),
            .I(N__44854));
    LocalMux I__10841 (
            .O(N__44895),
            .I(N__44851));
    Span4Mux_h I__10840 (
            .O(N__44892),
            .I(N__44840));
    Span4Mux_v I__10839 (
            .O(N__44889),
            .I(N__44840));
    Span4Mux_h I__10838 (
            .O(N__44884),
            .I(N__44840));
    LocalMux I__10837 (
            .O(N__44881),
            .I(N__44840));
    LocalMux I__10836 (
            .O(N__44878),
            .I(N__44840));
    Span4Mux_v I__10835 (
            .O(N__44871),
            .I(N__44833));
    Span4Mux_h I__10834 (
            .O(N__44866),
            .I(N__44833));
    LocalMux I__10833 (
            .O(N__44863),
            .I(N__44833));
    InMux I__10832 (
            .O(N__44862),
            .I(N__44830));
    Odrv4 I__10831 (
            .O(N__44859),
            .I(\c0.n9369 ));
    Odrv4 I__10830 (
            .O(N__44854),
            .I(\c0.n9369 ));
    Odrv4 I__10829 (
            .O(N__44851),
            .I(\c0.n9369 ));
    Odrv4 I__10828 (
            .O(N__44840),
            .I(\c0.n9369 ));
    Odrv4 I__10827 (
            .O(N__44833),
            .I(\c0.n9369 ));
    LocalMux I__10826 (
            .O(N__44830),
            .I(\c0.n9369 ));
    InMux I__10825 (
            .O(N__44817),
            .I(N__44814));
    LocalMux I__10824 (
            .O(N__44814),
            .I(N__44808));
    InMux I__10823 (
            .O(N__44813),
            .I(N__44805));
    InMux I__10822 (
            .O(N__44812),
            .I(N__44802));
    InMux I__10821 (
            .O(N__44811),
            .I(N__44795));
    Span4Mux_v I__10820 (
            .O(N__44808),
            .I(N__44792));
    LocalMux I__10819 (
            .O(N__44805),
            .I(N__44787));
    LocalMux I__10818 (
            .O(N__44802),
            .I(N__44787));
    InMux I__10817 (
            .O(N__44801),
            .I(N__44784));
    InMux I__10816 (
            .O(N__44800),
            .I(N__44781));
    InMux I__10815 (
            .O(N__44799),
            .I(N__44778));
    InMux I__10814 (
            .O(N__44798),
            .I(N__44773));
    LocalMux I__10813 (
            .O(N__44795),
            .I(N__44769));
    Span4Mux_h I__10812 (
            .O(N__44792),
            .I(N__44757));
    Span4Mux_v I__10811 (
            .O(N__44787),
            .I(N__44757));
    LocalMux I__10810 (
            .O(N__44784),
            .I(N__44757));
    LocalMux I__10809 (
            .O(N__44781),
            .I(N__44757));
    LocalMux I__10808 (
            .O(N__44778),
            .I(N__44757));
    InMux I__10807 (
            .O(N__44777),
            .I(N__44754));
    InMux I__10806 (
            .O(N__44776),
            .I(N__44751));
    LocalMux I__10805 (
            .O(N__44773),
            .I(N__44748));
    InMux I__10804 (
            .O(N__44772),
            .I(N__44745));
    Span4Mux_v I__10803 (
            .O(N__44769),
            .I(N__44742));
    InMux I__10802 (
            .O(N__44768),
            .I(N__44739));
    Span4Mux_v I__10801 (
            .O(N__44757),
            .I(N__44730));
    LocalMux I__10800 (
            .O(N__44754),
            .I(N__44730));
    LocalMux I__10799 (
            .O(N__44751),
            .I(N__44730));
    Span4Mux_h I__10798 (
            .O(N__44748),
            .I(N__44725));
    LocalMux I__10797 (
            .O(N__44745),
            .I(N__44725));
    Span4Mux_h I__10796 (
            .O(N__44742),
            .I(N__44719));
    LocalMux I__10795 (
            .O(N__44739),
            .I(N__44719));
    InMux I__10794 (
            .O(N__44738),
            .I(N__44715));
    InMux I__10793 (
            .O(N__44737),
            .I(N__44711));
    Span4Mux_h I__10792 (
            .O(N__44730),
            .I(N__44706));
    Span4Mux_v I__10791 (
            .O(N__44725),
            .I(N__44706));
    InMux I__10790 (
            .O(N__44724),
            .I(N__44703));
    Span4Mux_v I__10789 (
            .O(N__44719),
            .I(N__44699));
    InMux I__10788 (
            .O(N__44718),
            .I(N__44696));
    LocalMux I__10787 (
            .O(N__44715),
            .I(N__44693));
    InMux I__10786 (
            .O(N__44714),
            .I(N__44690));
    LocalMux I__10785 (
            .O(N__44711),
            .I(N__44687));
    Span4Mux_h I__10784 (
            .O(N__44706),
            .I(N__44682));
    LocalMux I__10783 (
            .O(N__44703),
            .I(N__44682));
    InMux I__10782 (
            .O(N__44702),
            .I(N__44679));
    Span4Mux_h I__10781 (
            .O(N__44699),
            .I(N__44668));
    LocalMux I__10780 (
            .O(N__44696),
            .I(N__44668));
    Span4Mux_h I__10779 (
            .O(N__44693),
            .I(N__44663));
    LocalMux I__10778 (
            .O(N__44690),
            .I(N__44663));
    Span4Mux_v I__10777 (
            .O(N__44687),
            .I(N__44656));
    Span4Mux_h I__10776 (
            .O(N__44682),
            .I(N__44656));
    LocalMux I__10775 (
            .O(N__44679),
            .I(N__44656));
    InMux I__10774 (
            .O(N__44678),
            .I(N__44653));
    InMux I__10773 (
            .O(N__44677),
            .I(N__44650));
    InMux I__10772 (
            .O(N__44676),
            .I(N__44647));
    InMux I__10771 (
            .O(N__44675),
            .I(N__44644));
    InMux I__10770 (
            .O(N__44674),
            .I(N__44641));
    InMux I__10769 (
            .O(N__44673),
            .I(N__44638));
    Odrv4 I__10768 (
            .O(N__44668),
            .I(\c0.n276 ));
    Odrv4 I__10767 (
            .O(N__44663),
            .I(\c0.n276 ));
    Odrv4 I__10766 (
            .O(N__44656),
            .I(\c0.n276 ));
    LocalMux I__10765 (
            .O(N__44653),
            .I(\c0.n276 ));
    LocalMux I__10764 (
            .O(N__44650),
            .I(\c0.n276 ));
    LocalMux I__10763 (
            .O(N__44647),
            .I(\c0.n276 ));
    LocalMux I__10762 (
            .O(N__44644),
            .I(\c0.n276 ));
    LocalMux I__10761 (
            .O(N__44641),
            .I(\c0.n276 ));
    LocalMux I__10760 (
            .O(N__44638),
            .I(\c0.n276 ));
    CascadeMux I__10759 (
            .O(N__44619),
            .I(N__44612));
    CascadeMux I__10758 (
            .O(N__44618),
            .I(N__44607));
    InMux I__10757 (
            .O(N__44617),
            .I(N__44596));
    CascadeMux I__10756 (
            .O(N__44616),
            .I(N__44593));
    InMux I__10755 (
            .O(N__44615),
            .I(N__44590));
    InMux I__10754 (
            .O(N__44612),
            .I(N__44587));
    InMux I__10753 (
            .O(N__44611),
            .I(N__44584));
    InMux I__10752 (
            .O(N__44610),
            .I(N__44580));
    InMux I__10751 (
            .O(N__44607),
            .I(N__44577));
    InMux I__10750 (
            .O(N__44606),
            .I(N__44574));
    InMux I__10749 (
            .O(N__44605),
            .I(N__44570));
    CascadeMux I__10748 (
            .O(N__44604),
            .I(N__44567));
    CascadeMux I__10747 (
            .O(N__44603),
            .I(N__44561));
    InMux I__10746 (
            .O(N__44602),
            .I(N__44558));
    InMux I__10745 (
            .O(N__44601),
            .I(N__44555));
    InMux I__10744 (
            .O(N__44600),
            .I(N__44552));
    InMux I__10743 (
            .O(N__44599),
            .I(N__44549));
    LocalMux I__10742 (
            .O(N__44596),
            .I(N__44546));
    InMux I__10741 (
            .O(N__44593),
            .I(N__44543));
    LocalMux I__10740 (
            .O(N__44590),
            .I(N__44539));
    LocalMux I__10739 (
            .O(N__44587),
            .I(N__44536));
    LocalMux I__10738 (
            .O(N__44584),
            .I(N__44533));
    InMux I__10737 (
            .O(N__44583),
            .I(N__44530));
    LocalMux I__10736 (
            .O(N__44580),
            .I(N__44523));
    LocalMux I__10735 (
            .O(N__44577),
            .I(N__44523));
    LocalMux I__10734 (
            .O(N__44574),
            .I(N__44523));
    InMux I__10733 (
            .O(N__44573),
            .I(N__44520));
    LocalMux I__10732 (
            .O(N__44570),
            .I(N__44517));
    InMux I__10731 (
            .O(N__44567),
            .I(N__44514));
    InMux I__10730 (
            .O(N__44566),
            .I(N__44507));
    InMux I__10729 (
            .O(N__44565),
            .I(N__44504));
    InMux I__10728 (
            .O(N__44564),
            .I(N__44501));
    InMux I__10727 (
            .O(N__44561),
            .I(N__44498));
    LocalMux I__10726 (
            .O(N__44558),
            .I(N__44493));
    LocalMux I__10725 (
            .O(N__44555),
            .I(N__44493));
    LocalMux I__10724 (
            .O(N__44552),
            .I(N__44486));
    LocalMux I__10723 (
            .O(N__44549),
            .I(N__44486));
    Span4Mux_h I__10722 (
            .O(N__44546),
            .I(N__44486));
    LocalMux I__10721 (
            .O(N__44543),
            .I(N__44483));
    InMux I__10720 (
            .O(N__44542),
            .I(N__44480));
    Span4Mux_h I__10719 (
            .O(N__44539),
            .I(N__44473));
    Span4Mux_s3_v I__10718 (
            .O(N__44536),
            .I(N__44473));
    Span4Mux_s3_v I__10717 (
            .O(N__44533),
            .I(N__44473));
    LocalMux I__10716 (
            .O(N__44530),
            .I(N__44470));
    Span4Mux_v I__10715 (
            .O(N__44523),
            .I(N__44467));
    LocalMux I__10714 (
            .O(N__44520),
            .I(N__44460));
    Span4Mux_h I__10713 (
            .O(N__44517),
            .I(N__44460));
    LocalMux I__10712 (
            .O(N__44514),
            .I(N__44460));
    InMux I__10711 (
            .O(N__44513),
            .I(N__44457));
    InMux I__10710 (
            .O(N__44512),
            .I(N__44454));
    InMux I__10709 (
            .O(N__44511),
            .I(N__44451));
    InMux I__10708 (
            .O(N__44510),
            .I(N__44448));
    LocalMux I__10707 (
            .O(N__44507),
            .I(N__44445));
    LocalMux I__10706 (
            .O(N__44504),
            .I(N__44442));
    LocalMux I__10705 (
            .O(N__44501),
            .I(N__44437));
    LocalMux I__10704 (
            .O(N__44498),
            .I(N__44437));
    Span4Mux_h I__10703 (
            .O(N__44493),
            .I(N__44430));
    Span4Mux_h I__10702 (
            .O(N__44486),
            .I(N__44430));
    Span4Mux_h I__10701 (
            .O(N__44483),
            .I(N__44430));
    LocalMux I__10700 (
            .O(N__44480),
            .I(N__44425));
    Sp12to4 I__10699 (
            .O(N__44473),
            .I(N__44425));
    Span4Mux_h I__10698 (
            .O(N__44470),
            .I(N__44415));
    Span4Mux_h I__10697 (
            .O(N__44467),
            .I(N__44415));
    Span4Mux_v I__10696 (
            .O(N__44460),
            .I(N__44415));
    LocalMux I__10695 (
            .O(N__44457),
            .I(N__44415));
    LocalMux I__10694 (
            .O(N__44454),
            .I(N__44407));
    LocalMux I__10693 (
            .O(N__44451),
            .I(N__44407));
    LocalMux I__10692 (
            .O(N__44448),
            .I(N__44407));
    Span4Mux_h I__10691 (
            .O(N__44445),
            .I(N__44400));
    Span4Mux_h I__10690 (
            .O(N__44442),
            .I(N__44400));
    Span4Mux_h I__10689 (
            .O(N__44437),
            .I(N__44400));
    Sp12to4 I__10688 (
            .O(N__44430),
            .I(N__44395));
    Span12Mux_s10_h I__10687 (
            .O(N__44425),
            .I(N__44395));
    InMux I__10686 (
            .O(N__44424),
            .I(N__44392));
    Span4Mux_h I__10685 (
            .O(N__44415),
            .I(N__44389));
    InMux I__10684 (
            .O(N__44414),
            .I(N__44386));
    Odrv12 I__10683 (
            .O(N__44407),
            .I(FRAME_MATCHER_i_31__N_1275));
    Odrv4 I__10682 (
            .O(N__44400),
            .I(FRAME_MATCHER_i_31__N_1275));
    Odrv12 I__10681 (
            .O(N__44395),
            .I(FRAME_MATCHER_i_31__N_1275));
    LocalMux I__10680 (
            .O(N__44392),
            .I(FRAME_MATCHER_i_31__N_1275));
    Odrv4 I__10679 (
            .O(N__44389),
            .I(FRAME_MATCHER_i_31__N_1275));
    LocalMux I__10678 (
            .O(N__44386),
            .I(FRAME_MATCHER_i_31__N_1275));
    InMux I__10677 (
            .O(N__44373),
            .I(N__44366));
    InMux I__10676 (
            .O(N__44372),
            .I(N__44366));
    CascadeMux I__10675 (
            .O(N__44371),
            .I(N__44363));
    LocalMux I__10674 (
            .O(N__44366),
            .I(N__44360));
    InMux I__10673 (
            .O(N__44363),
            .I(N__44357));
    Span4Mux_v I__10672 (
            .O(N__44360),
            .I(N__44354));
    LocalMux I__10671 (
            .O(N__44357),
            .I(\c0.FRAME_MATCHER_state_22 ));
    Odrv4 I__10670 (
            .O(N__44354),
            .I(\c0.FRAME_MATCHER_state_22 ));
    SRMux I__10669 (
            .O(N__44349),
            .I(N__44346));
    LocalMux I__10668 (
            .O(N__44346),
            .I(N__44343));
    Span4Mux_v I__10667 (
            .O(N__44343),
            .I(N__44340));
    Span4Mux_h I__10666 (
            .O(N__44340),
            .I(N__44337));
    Odrv4 I__10665 (
            .O(N__44337),
            .I(\c0.n16714 ));
    InMux I__10664 (
            .O(N__44334),
            .I(N__44328));
    InMux I__10663 (
            .O(N__44333),
            .I(N__44328));
    LocalMux I__10662 (
            .O(N__44328),
            .I(data_out_1_7));
    InMux I__10661 (
            .O(N__44325),
            .I(N__44322));
    LocalMux I__10660 (
            .O(N__44322),
            .I(N__44319));
    Span4Mux_v I__10659 (
            .O(N__44319),
            .I(N__44316));
    Odrv4 I__10658 (
            .O(N__44316),
            .I(\c0.n8_adj_2352 ));
    CascadeMux I__10657 (
            .O(N__44313),
            .I(n5142_cascade_));
    InMux I__10656 (
            .O(N__44310),
            .I(N__44307));
    LocalMux I__10655 (
            .O(N__44307),
            .I(N__44304));
    Odrv4 I__10654 (
            .O(N__44304),
            .I(\c0.tx.n6759 ));
    InMux I__10653 (
            .O(N__44301),
            .I(N__44298));
    LocalMux I__10652 (
            .O(N__44298),
            .I(\c0.tx.n13702 ));
    InMux I__10651 (
            .O(N__44295),
            .I(N__44292));
    LocalMux I__10650 (
            .O(N__44292),
            .I(\c0.tx_active_prev ));
    InMux I__10649 (
            .O(N__44289),
            .I(N__44282));
    InMux I__10648 (
            .O(N__44288),
            .I(N__44279));
    InMux I__10647 (
            .O(N__44287),
            .I(N__44274));
    InMux I__10646 (
            .O(N__44286),
            .I(N__44274));
    InMux I__10645 (
            .O(N__44285),
            .I(N__44271));
    LocalMux I__10644 (
            .O(N__44282),
            .I(N__44268));
    LocalMux I__10643 (
            .O(N__44279),
            .I(N__44265));
    LocalMux I__10642 (
            .O(N__44274),
            .I(N__44262));
    LocalMux I__10641 (
            .O(N__44271),
            .I(N__44259));
    Span4Mux_s2_v I__10640 (
            .O(N__44268),
            .I(N__44256));
    Span4Mux_h I__10639 (
            .O(N__44265),
            .I(N__44253));
    Span4Mux_h I__10638 (
            .O(N__44262),
            .I(N__44250));
    Span4Mux_h I__10637 (
            .O(N__44259),
            .I(N__44245));
    Span4Mux_h I__10636 (
            .O(N__44256),
            .I(N__44245));
    Odrv4 I__10635 (
            .O(N__44253),
            .I(\c0.data_out_5_5 ));
    Odrv4 I__10634 (
            .O(N__44250),
            .I(\c0.data_out_5_5 ));
    Odrv4 I__10633 (
            .O(N__44245),
            .I(\c0.data_out_5_5 ));
    InMux I__10632 (
            .O(N__44238),
            .I(N__44235));
    LocalMux I__10631 (
            .O(N__44235),
            .I(N__44232));
    Span12Mux_s2_v I__10630 (
            .O(N__44232),
            .I(N__44229));
    Odrv12 I__10629 (
            .O(N__44229),
            .I(\c0.n5_adj_2163 ));
    CascadeMux I__10628 (
            .O(N__44226),
            .I(\c0.n17581_cascade_ ));
    CascadeMux I__10627 (
            .O(N__44223),
            .I(N__44220));
    InMux I__10626 (
            .O(N__44220),
            .I(N__44217));
    LocalMux I__10625 (
            .O(N__44217),
            .I(n10_adj_2432));
    InMux I__10624 (
            .O(N__44214),
            .I(N__44209));
    CascadeMux I__10623 (
            .O(N__44213),
            .I(N__44205));
    CascadeMux I__10622 (
            .O(N__44212),
            .I(N__44200));
    LocalMux I__10621 (
            .O(N__44209),
            .I(N__44197));
    InMux I__10620 (
            .O(N__44208),
            .I(N__44194));
    InMux I__10619 (
            .O(N__44205),
            .I(N__44188));
    InMux I__10618 (
            .O(N__44204),
            .I(N__44181));
    InMux I__10617 (
            .O(N__44203),
            .I(N__44181));
    InMux I__10616 (
            .O(N__44200),
            .I(N__44181));
    Span4Mux_v I__10615 (
            .O(N__44197),
            .I(N__44173));
    LocalMux I__10614 (
            .O(N__44194),
            .I(N__44173));
    CascadeMux I__10613 (
            .O(N__44193),
            .I(N__44170));
    CascadeMux I__10612 (
            .O(N__44192),
            .I(N__44167));
    CascadeMux I__10611 (
            .O(N__44191),
            .I(N__44164));
    LocalMux I__10610 (
            .O(N__44188),
            .I(N__44161));
    LocalMux I__10609 (
            .O(N__44181),
            .I(N__44158));
    InMux I__10608 (
            .O(N__44180),
            .I(N__44155));
    InMux I__10607 (
            .O(N__44179),
            .I(N__44152));
    InMux I__10606 (
            .O(N__44178),
            .I(N__44149));
    Span4Mux_h I__10605 (
            .O(N__44173),
            .I(N__44146));
    InMux I__10604 (
            .O(N__44170),
            .I(N__44139));
    InMux I__10603 (
            .O(N__44167),
            .I(N__44139));
    InMux I__10602 (
            .O(N__44164),
            .I(N__44139));
    Span4Mux_h I__10601 (
            .O(N__44161),
            .I(N__44134));
    Span4Mux_v I__10600 (
            .O(N__44158),
            .I(N__44134));
    LocalMux I__10599 (
            .O(N__44155),
            .I(\c0.tx.r_SM_Main_1 ));
    LocalMux I__10598 (
            .O(N__44152),
            .I(\c0.tx.r_SM_Main_1 ));
    LocalMux I__10597 (
            .O(N__44149),
            .I(\c0.tx.r_SM_Main_1 ));
    Odrv4 I__10596 (
            .O(N__44146),
            .I(\c0.tx.r_SM_Main_1 ));
    LocalMux I__10595 (
            .O(N__44139),
            .I(\c0.tx.r_SM_Main_1 ));
    Odrv4 I__10594 (
            .O(N__44134),
            .I(\c0.tx.r_SM_Main_1 ));
    InMux I__10593 (
            .O(N__44121),
            .I(N__44118));
    LocalMux I__10592 (
            .O(N__44118),
            .I(\c0.tx.n10613 ));
    InMux I__10591 (
            .O(N__44115),
            .I(N__44112));
    LocalMux I__10590 (
            .O(N__44112),
            .I(\c0.tx.n12_adj_2134 ));
    CascadeMux I__10589 (
            .O(N__44109),
            .I(\c0.n8_cascade_ ));
    CascadeMux I__10588 (
            .O(N__44106),
            .I(N__44100));
    InMux I__10587 (
            .O(N__44105),
            .I(N__44094));
    InMux I__10586 (
            .O(N__44104),
            .I(N__44091));
    InMux I__10585 (
            .O(N__44103),
            .I(N__44088));
    InMux I__10584 (
            .O(N__44100),
            .I(N__44085));
    InMux I__10583 (
            .O(N__44099),
            .I(N__44082));
    CascadeMux I__10582 (
            .O(N__44098),
            .I(N__44079));
    CascadeMux I__10581 (
            .O(N__44097),
            .I(N__44076));
    LocalMux I__10580 (
            .O(N__44094),
            .I(N__44072));
    LocalMux I__10579 (
            .O(N__44091),
            .I(N__44069));
    LocalMux I__10578 (
            .O(N__44088),
            .I(N__44066));
    LocalMux I__10577 (
            .O(N__44085),
            .I(N__44063));
    LocalMux I__10576 (
            .O(N__44082),
            .I(N__44060));
    InMux I__10575 (
            .O(N__44079),
            .I(N__44055));
    InMux I__10574 (
            .O(N__44076),
            .I(N__44055));
    CascadeMux I__10573 (
            .O(N__44075),
            .I(N__44052));
    Span4Mux_h I__10572 (
            .O(N__44072),
            .I(N__44049));
    Span4Mux_h I__10571 (
            .O(N__44069),
            .I(N__44044));
    Span4Mux_h I__10570 (
            .O(N__44066),
            .I(N__44044));
    Span4Mux_h I__10569 (
            .O(N__44063),
            .I(N__44039));
    Span4Mux_h I__10568 (
            .O(N__44060),
            .I(N__44039));
    LocalMux I__10567 (
            .O(N__44055),
            .I(N__44036));
    InMux I__10566 (
            .O(N__44052),
            .I(N__44033));
    Odrv4 I__10565 (
            .O(N__44049),
            .I(n9257));
    Odrv4 I__10564 (
            .O(N__44044),
            .I(n9257));
    Odrv4 I__10563 (
            .O(N__44039),
            .I(n9257));
    Odrv12 I__10562 (
            .O(N__44036),
            .I(n9257));
    LocalMux I__10561 (
            .O(N__44033),
            .I(n9257));
    InMux I__10560 (
            .O(N__44022),
            .I(N__44019));
    LocalMux I__10559 (
            .O(N__44019),
            .I(\c0.n65_adj_2192 ));
    InMux I__10558 (
            .O(N__44016),
            .I(N__44011));
    InMux I__10557 (
            .O(N__44015),
            .I(N__44008));
    InMux I__10556 (
            .O(N__44014),
            .I(N__44005));
    LocalMux I__10555 (
            .O(N__44011),
            .I(N__44000));
    LocalMux I__10554 (
            .O(N__44008),
            .I(N__43993));
    LocalMux I__10553 (
            .O(N__44005),
            .I(N__43993));
    CascadeMux I__10552 (
            .O(N__44004),
            .I(N__43990));
    CascadeMux I__10551 (
            .O(N__44003),
            .I(N__43987));
    Span4Mux_h I__10550 (
            .O(N__44000),
            .I(N__43982));
    InMux I__10549 (
            .O(N__43999),
            .I(N__43977));
    InMux I__10548 (
            .O(N__43998),
            .I(N__43977));
    Span4Mux_h I__10547 (
            .O(N__43993),
            .I(N__43974));
    InMux I__10546 (
            .O(N__43990),
            .I(N__43965));
    InMux I__10545 (
            .O(N__43987),
            .I(N__43965));
    InMux I__10544 (
            .O(N__43986),
            .I(N__43965));
    InMux I__10543 (
            .O(N__43985),
            .I(N__43965));
    Odrv4 I__10542 (
            .O(N__43982),
            .I(\c0.tx.r_SM_Main_0 ));
    LocalMux I__10541 (
            .O(N__43977),
            .I(\c0.tx.r_SM_Main_0 ));
    Odrv4 I__10540 (
            .O(N__43974),
            .I(\c0.tx.r_SM_Main_0 ));
    LocalMux I__10539 (
            .O(N__43965),
            .I(\c0.tx.r_SM_Main_0 ));
    InMux I__10538 (
            .O(N__43956),
            .I(N__43953));
    LocalMux I__10537 (
            .O(N__43953),
            .I(N__43947));
    InMux I__10536 (
            .O(N__43952),
            .I(N__43942));
    InMux I__10535 (
            .O(N__43951),
            .I(N__43942));
    InMux I__10534 (
            .O(N__43950),
            .I(N__43939));
    Span4Mux_v I__10533 (
            .O(N__43947),
            .I(N__43933));
    LocalMux I__10532 (
            .O(N__43942),
            .I(N__43930));
    LocalMux I__10531 (
            .O(N__43939),
            .I(N__43927));
    InMux I__10530 (
            .O(N__43938),
            .I(N__43924));
    InMux I__10529 (
            .O(N__43937),
            .I(N__43919));
    InMux I__10528 (
            .O(N__43936),
            .I(N__43919));
    Odrv4 I__10527 (
            .O(N__43933),
            .I(\c0.tx.n83 ));
    Odrv12 I__10526 (
            .O(N__43930),
            .I(\c0.tx.n83 ));
    Odrv12 I__10525 (
            .O(N__43927),
            .I(\c0.tx.n83 ));
    LocalMux I__10524 (
            .O(N__43924),
            .I(\c0.tx.n83 ));
    LocalMux I__10523 (
            .O(N__43919),
            .I(\c0.tx.n83 ));
    InMux I__10522 (
            .O(N__43908),
            .I(N__43905));
    LocalMux I__10521 (
            .O(N__43905),
            .I(N__43902));
    Odrv4 I__10520 (
            .O(N__43902),
            .I(n10_adj_2422));
    CascadeMux I__10519 (
            .O(N__43899),
            .I(\c0.tx.n77_cascade_ ));
    InMux I__10518 (
            .O(N__43896),
            .I(N__43893));
    LocalMux I__10517 (
            .O(N__43893),
            .I(N__43890));
    Odrv4 I__10516 (
            .O(N__43890),
            .I(\c0.tx.n12 ));
    IoInMux I__10515 (
            .O(N__43887),
            .I(N__43884));
    LocalMux I__10514 (
            .O(N__43884),
            .I(N__43881));
    IoSpan4Mux I__10513 (
            .O(N__43881),
            .I(N__43877));
    InMux I__10512 (
            .O(N__43880),
            .I(N__43874));
    Span4Mux_s3_v I__10511 (
            .O(N__43877),
            .I(N__43871));
    LocalMux I__10510 (
            .O(N__43874),
            .I(N__43868));
    Span4Mux_h I__10509 (
            .O(N__43871),
            .I(N__43863));
    Span4Mux_h I__10508 (
            .O(N__43868),
            .I(N__43863));
    Span4Mux_h I__10507 (
            .O(N__43863),
            .I(N__43859));
    InMux I__10506 (
            .O(N__43862),
            .I(N__43856));
    Odrv4 I__10505 (
            .O(N__43859),
            .I(tx_o));
    LocalMux I__10504 (
            .O(N__43856),
            .I(tx_o));
    InMux I__10503 (
            .O(N__43851),
            .I(N__43848));
    LocalMux I__10502 (
            .O(N__43848),
            .I(\c0.tx.n10 ));
    InMux I__10501 (
            .O(N__43845),
            .I(N__43837));
    InMux I__10500 (
            .O(N__43844),
            .I(N__43831));
    InMux I__10499 (
            .O(N__43843),
            .I(N__43831));
    CascadeMux I__10498 (
            .O(N__43842),
            .I(N__43828));
    InMux I__10497 (
            .O(N__43841),
            .I(N__43825));
    InMux I__10496 (
            .O(N__43840),
            .I(N__43822));
    LocalMux I__10495 (
            .O(N__43837),
            .I(N__43819));
    InMux I__10494 (
            .O(N__43836),
            .I(N__43816));
    LocalMux I__10493 (
            .O(N__43831),
            .I(N__43810));
    InMux I__10492 (
            .O(N__43828),
            .I(N__43807));
    LocalMux I__10491 (
            .O(N__43825),
            .I(N__43804));
    LocalMux I__10490 (
            .O(N__43822),
            .I(N__43801));
    Span4Mux_s2_v I__10489 (
            .O(N__43819),
            .I(N__43796));
    LocalMux I__10488 (
            .O(N__43816),
            .I(N__43796));
    InMux I__10487 (
            .O(N__43815),
            .I(N__43793));
    InMux I__10486 (
            .O(N__43814),
            .I(N__43788));
    InMux I__10485 (
            .O(N__43813),
            .I(N__43788));
    Span4Mux_h I__10484 (
            .O(N__43810),
            .I(N__43785));
    LocalMux I__10483 (
            .O(N__43807),
            .I(N__43778));
    Span4Mux_v I__10482 (
            .O(N__43804),
            .I(N__43778));
    Span4Mux_h I__10481 (
            .O(N__43801),
            .I(N__43778));
    Span4Mux_v I__10480 (
            .O(N__43796),
            .I(N__43775));
    LocalMux I__10479 (
            .O(N__43793),
            .I(byte_transmit_counter_4));
    LocalMux I__10478 (
            .O(N__43788),
            .I(byte_transmit_counter_4));
    Odrv4 I__10477 (
            .O(N__43785),
            .I(byte_transmit_counter_4));
    Odrv4 I__10476 (
            .O(N__43778),
            .I(byte_transmit_counter_4));
    Odrv4 I__10475 (
            .O(N__43775),
            .I(byte_transmit_counter_4));
    InMux I__10474 (
            .O(N__43764),
            .I(N__43761));
    LocalMux I__10473 (
            .O(N__43761),
            .I(n10_adj_2443));
    InMux I__10472 (
            .O(N__43758),
            .I(N__43754));
    InMux I__10471 (
            .O(N__43757),
            .I(N__43751));
    LocalMux I__10470 (
            .O(N__43754),
            .I(N__43748));
    LocalMux I__10469 (
            .O(N__43751),
            .I(r_Tx_Data_6));
    Odrv4 I__10468 (
            .O(N__43748),
            .I(r_Tx_Data_6));
    InMux I__10467 (
            .O(N__43743),
            .I(N__43740));
    LocalMux I__10466 (
            .O(N__43740),
            .I(N__43737));
    Span4Mux_v I__10465 (
            .O(N__43737),
            .I(N__43733));
    CascadeMux I__10464 (
            .O(N__43736),
            .I(N__43730));
    Span4Mux_h I__10463 (
            .O(N__43733),
            .I(N__43727));
    InMux I__10462 (
            .O(N__43730),
            .I(N__43724));
    Odrv4 I__10461 (
            .O(N__43727),
            .I(rand_setpoint_5));
    LocalMux I__10460 (
            .O(N__43724),
            .I(rand_setpoint_5));
    CascadeMux I__10459 (
            .O(N__43719),
            .I(N__43712));
    CascadeMux I__10458 (
            .O(N__43718),
            .I(N__43709));
    InMux I__10457 (
            .O(N__43717),
            .I(N__43706));
    CascadeMux I__10456 (
            .O(N__43716),
            .I(N__43703));
    CascadeMux I__10455 (
            .O(N__43715),
            .I(N__43700));
    InMux I__10454 (
            .O(N__43712),
            .I(N__43697));
    InMux I__10453 (
            .O(N__43709),
            .I(N__43694));
    LocalMux I__10452 (
            .O(N__43706),
            .I(N__43690));
    InMux I__10451 (
            .O(N__43703),
            .I(N__43687));
    InMux I__10450 (
            .O(N__43700),
            .I(N__43684));
    LocalMux I__10449 (
            .O(N__43697),
            .I(N__43681));
    LocalMux I__10448 (
            .O(N__43694),
            .I(N__43678));
    InMux I__10447 (
            .O(N__43693),
            .I(N__43675));
    Span4Mux_h I__10446 (
            .O(N__43690),
            .I(N__43668));
    LocalMux I__10445 (
            .O(N__43687),
            .I(N__43668));
    LocalMux I__10444 (
            .O(N__43684),
            .I(N__43668));
    Span4Mux_v I__10443 (
            .O(N__43681),
            .I(N__43665));
    Span4Mux_h I__10442 (
            .O(N__43678),
            .I(N__43662));
    LocalMux I__10441 (
            .O(N__43675),
            .I(N__43657));
    Span4Mux_v I__10440 (
            .O(N__43668),
            .I(N__43657));
    Odrv4 I__10439 (
            .O(N__43665),
            .I(n2594));
    Odrv4 I__10438 (
            .O(N__43662),
            .I(n2594));
    Odrv4 I__10437 (
            .O(N__43657),
            .I(n2594));
    CascadeMux I__10436 (
            .O(N__43650),
            .I(N__43647));
    InMux I__10435 (
            .O(N__43647),
            .I(N__43643));
    CascadeMux I__10434 (
            .O(N__43646),
            .I(N__43640));
    LocalMux I__10433 (
            .O(N__43643),
            .I(N__43637));
    InMux I__10432 (
            .O(N__43640),
            .I(N__43634));
    Odrv12 I__10431 (
            .O(N__43637),
            .I(rand_setpoint_13));
    LocalMux I__10430 (
            .O(N__43634),
            .I(rand_setpoint_13));
    InMux I__10429 (
            .O(N__43629),
            .I(N__43626));
    LocalMux I__10428 (
            .O(N__43626),
            .I(N__43621));
    InMux I__10427 (
            .O(N__43625),
            .I(N__43616));
    InMux I__10426 (
            .O(N__43624),
            .I(N__43616));
    Span12Mux_s6_v I__10425 (
            .O(N__43621),
            .I(N__43613));
    LocalMux I__10424 (
            .O(N__43616),
            .I(\c0.data_out_7_5 ));
    Odrv12 I__10423 (
            .O(N__43613),
            .I(\c0.data_out_7_5 ));
    CascadeMux I__10422 (
            .O(N__43608),
            .I(N__43605));
    InMux I__10421 (
            .O(N__43605),
            .I(N__43602));
    LocalMux I__10420 (
            .O(N__43602),
            .I(N__43598));
    InMux I__10419 (
            .O(N__43601),
            .I(N__43595));
    Span4Mux_h I__10418 (
            .O(N__43598),
            .I(N__43592));
    LocalMux I__10417 (
            .O(N__43595),
            .I(r_Tx_Data_7));
    Odrv4 I__10416 (
            .O(N__43592),
            .I(r_Tx_Data_7));
    InMux I__10415 (
            .O(N__43587),
            .I(N__43584));
    LocalMux I__10414 (
            .O(N__43584),
            .I(N__43581));
    Span4Mux_h I__10413 (
            .O(N__43581),
            .I(N__43578));
    Odrv4 I__10412 (
            .O(N__43578),
            .I(\c0.data_out_1_1 ));
    InMux I__10411 (
            .O(N__43575),
            .I(N__43571));
    InMux I__10410 (
            .O(N__43574),
            .I(N__43568));
    LocalMux I__10409 (
            .O(N__43571),
            .I(data_out_0_1));
    LocalMux I__10408 (
            .O(N__43568),
            .I(data_out_0_1));
    InMux I__10407 (
            .O(N__43563),
            .I(N__43560));
    LocalMux I__10406 (
            .O(N__43560),
            .I(n1_adj_2449));
    InMux I__10405 (
            .O(N__43557),
            .I(N__43554));
    LocalMux I__10404 (
            .O(N__43554),
            .I(\c0.n12630 ));
    InMux I__10403 (
            .O(N__43551),
            .I(N__43546));
    InMux I__10402 (
            .O(N__43550),
            .I(N__43543));
    InMux I__10401 (
            .O(N__43549),
            .I(N__43540));
    LocalMux I__10400 (
            .O(N__43546),
            .I(\c0.data_out_7_0 ));
    LocalMux I__10399 (
            .O(N__43543),
            .I(\c0.data_out_7_0 ));
    LocalMux I__10398 (
            .O(N__43540),
            .I(\c0.data_out_7_0 ));
    InMux I__10397 (
            .O(N__43533),
            .I(N__43530));
    LocalMux I__10396 (
            .O(N__43530),
            .I(N__43526));
    InMux I__10395 (
            .O(N__43529),
            .I(N__43523));
    Odrv4 I__10394 (
            .O(N__43526),
            .I(\c0.n10395 ));
    LocalMux I__10393 (
            .O(N__43523),
            .I(\c0.n10395 ));
    CascadeMux I__10392 (
            .O(N__43518),
            .I(\c0.n10_adj_2189_cascade_ ));
    InMux I__10391 (
            .O(N__43515),
            .I(N__43512));
    LocalMux I__10390 (
            .O(N__43512),
            .I(N__43508));
    InMux I__10389 (
            .O(N__43511),
            .I(N__43505));
    Span4Mux_h I__10388 (
            .O(N__43508),
            .I(N__43502));
    LocalMux I__10387 (
            .O(N__43505),
            .I(r_Tx_Data_0));
    Odrv4 I__10386 (
            .O(N__43502),
            .I(r_Tx_Data_0));
    InMux I__10385 (
            .O(N__43497),
            .I(N__43494));
    LocalMux I__10384 (
            .O(N__43494),
            .I(\c0.n8_adj_2157 ));
    InMux I__10383 (
            .O(N__43491),
            .I(N__43488));
    LocalMux I__10382 (
            .O(N__43488),
            .I(\c0.n15_adj_2177 ));
    CascadeMux I__10381 (
            .O(N__43485),
            .I(N__43482));
    InMux I__10380 (
            .O(N__43482),
            .I(N__43479));
    LocalMux I__10379 (
            .O(N__43479),
            .I(N__43476));
    Span4Mux_v I__10378 (
            .O(N__43476),
            .I(N__43473));
    Odrv4 I__10377 (
            .O(N__43473),
            .I(\c0.n17270 ));
    InMux I__10376 (
            .O(N__43470),
            .I(N__43466));
    InMux I__10375 (
            .O(N__43469),
            .I(N__43462));
    LocalMux I__10374 (
            .O(N__43466),
            .I(N__43459));
    InMux I__10373 (
            .O(N__43465),
            .I(N__43456));
    LocalMux I__10372 (
            .O(N__43462),
            .I(N__43453));
    Span4Mux_v I__10371 (
            .O(N__43459),
            .I(N__43450));
    LocalMux I__10370 (
            .O(N__43456),
            .I(N__43447));
    Span12Mux_v I__10369 (
            .O(N__43453),
            .I(N__43444));
    Span4Mux_h I__10368 (
            .O(N__43450),
            .I(N__43441));
    Span4Mux_h I__10367 (
            .O(N__43447),
            .I(N__43438));
    Odrv12 I__10366 (
            .O(N__43444),
            .I(\c0.data_out_7_2 ));
    Odrv4 I__10365 (
            .O(N__43441),
            .I(\c0.data_out_7_2 ));
    Odrv4 I__10364 (
            .O(N__43438),
            .I(\c0.data_out_7_2 ));
    InMux I__10363 (
            .O(N__43431),
            .I(N__43428));
    LocalMux I__10362 (
            .O(N__43428),
            .I(\c0.n10316 ));
    InMux I__10361 (
            .O(N__43425),
            .I(N__43422));
    LocalMux I__10360 (
            .O(N__43422),
            .I(\c0.n17201 ));
    CascadeMux I__10359 (
            .O(N__43419),
            .I(\c0.n10316_cascade_ ));
    InMux I__10358 (
            .O(N__43416),
            .I(N__43410));
    InMux I__10357 (
            .O(N__43415),
            .I(N__43410));
    LocalMux I__10356 (
            .O(N__43410),
            .I(\c0.n17177 ));
    InMux I__10355 (
            .O(N__43407),
            .I(N__43403));
    InMux I__10354 (
            .O(N__43406),
            .I(N__43400));
    LocalMux I__10353 (
            .O(N__43403),
            .I(N__43395));
    LocalMux I__10352 (
            .O(N__43400),
            .I(N__43392));
    InMux I__10351 (
            .O(N__43399),
            .I(N__43387));
    InMux I__10350 (
            .O(N__43398),
            .I(N__43387));
    Span4Mux_h I__10349 (
            .O(N__43395),
            .I(N__43383));
    Span4Mux_v I__10348 (
            .O(N__43392),
            .I(N__43378));
    LocalMux I__10347 (
            .O(N__43387),
            .I(N__43378));
    InMux I__10346 (
            .O(N__43386),
            .I(N__43375));
    Span4Mux_v I__10345 (
            .O(N__43383),
            .I(N__43372));
    Span4Mux_h I__10344 (
            .O(N__43378),
            .I(N__43369));
    LocalMux I__10343 (
            .O(N__43375),
            .I(data_out_8_6));
    Odrv4 I__10342 (
            .O(N__43372),
            .I(data_out_8_6));
    Odrv4 I__10341 (
            .O(N__43369),
            .I(data_out_8_6));
    InMux I__10340 (
            .O(N__43362),
            .I(N__43353));
    InMux I__10339 (
            .O(N__43361),
            .I(N__43353));
    InMux I__10338 (
            .O(N__43360),
            .I(N__43350));
    InMux I__10337 (
            .O(N__43359),
            .I(N__43345));
    InMux I__10336 (
            .O(N__43358),
            .I(N__43345));
    LocalMux I__10335 (
            .O(N__43353),
            .I(N__43342));
    LocalMux I__10334 (
            .O(N__43350),
            .I(N__43337));
    LocalMux I__10333 (
            .O(N__43345),
            .I(N__43337));
    Span4Mux_v I__10332 (
            .O(N__43342),
            .I(N__43334));
    Span4Mux_v I__10331 (
            .O(N__43337),
            .I(N__43331));
    Sp12to4 I__10330 (
            .O(N__43334),
            .I(N__43326));
    Sp12to4 I__10329 (
            .O(N__43331),
            .I(N__43326));
    Span12Mux_h I__10328 (
            .O(N__43326),
            .I(N__43323));
    Odrv12 I__10327 (
            .O(N__43323),
            .I(\c0.data_out_6__1__N_537 ));
    InMux I__10326 (
            .O(N__43320),
            .I(N__43317));
    LocalMux I__10325 (
            .O(N__43317),
            .I(N__43314));
    Span4Mux_v I__10324 (
            .O(N__43314),
            .I(N__43310));
    InMux I__10323 (
            .O(N__43313),
            .I(N__43305));
    Sp12to4 I__10322 (
            .O(N__43310),
            .I(N__43302));
    InMux I__10321 (
            .O(N__43309),
            .I(N__43297));
    InMux I__10320 (
            .O(N__43308),
            .I(N__43297));
    LocalMux I__10319 (
            .O(N__43305),
            .I(\c0.data_out_7_7 ));
    Odrv12 I__10318 (
            .O(N__43302),
            .I(\c0.data_out_7_7 ));
    LocalMux I__10317 (
            .O(N__43297),
            .I(\c0.data_out_7_7 ));
    InMux I__10316 (
            .O(N__43290),
            .I(N__43287));
    LocalMux I__10315 (
            .O(N__43287),
            .I(n10_adj_2483));
    InMux I__10314 (
            .O(N__43284),
            .I(N__43281));
    LocalMux I__10313 (
            .O(N__43281),
            .I(N__43277));
    InMux I__10312 (
            .O(N__43280),
            .I(N__43274));
    Span4Mux_v I__10311 (
            .O(N__43277),
            .I(N__43271));
    LocalMux I__10310 (
            .O(N__43274),
            .I(\c0.data_out_3_6 ));
    Odrv4 I__10309 (
            .O(N__43271),
            .I(\c0.data_out_3_6 ));
    CascadeMux I__10308 (
            .O(N__43266),
            .I(N__43261));
    InMux I__10307 (
            .O(N__43265),
            .I(N__43256));
    InMux I__10306 (
            .O(N__43264),
            .I(N__43256));
    InMux I__10305 (
            .O(N__43261),
            .I(N__43253));
    LocalMux I__10304 (
            .O(N__43256),
            .I(N__43250));
    LocalMux I__10303 (
            .O(N__43253),
            .I(N__43245));
    Span4Mux_v I__10302 (
            .O(N__43250),
            .I(N__43245));
    Odrv4 I__10301 (
            .O(N__43245),
            .I(\c0.FRAME_MATCHER_state_25 ));
    SRMux I__10300 (
            .O(N__43242),
            .I(N__43239));
    LocalMux I__10299 (
            .O(N__43239),
            .I(N__43236));
    Span4Mux_v I__10298 (
            .O(N__43236),
            .I(N__43233));
    Odrv4 I__10297 (
            .O(N__43233),
            .I(\c0.n16690 ));
    CascadeMux I__10296 (
            .O(N__43230),
            .I(N__43226));
    InMux I__10295 (
            .O(N__43229),
            .I(N__43222));
    InMux I__10294 (
            .O(N__43226),
            .I(N__43219));
    InMux I__10293 (
            .O(N__43225),
            .I(N__43216));
    LocalMux I__10292 (
            .O(N__43222),
            .I(N__43211));
    LocalMux I__10291 (
            .O(N__43219),
            .I(N__43211));
    LocalMux I__10290 (
            .O(N__43216),
            .I(N__43206));
    Span4Mux_v I__10289 (
            .O(N__43211),
            .I(N__43206));
    Odrv4 I__10288 (
            .O(N__43206),
            .I(\c0.FRAME_MATCHER_state_26 ));
    SRMux I__10287 (
            .O(N__43203),
            .I(N__43200));
    LocalMux I__10286 (
            .O(N__43200),
            .I(N__43197));
    Span4Mux_h I__10285 (
            .O(N__43197),
            .I(N__43194));
    Odrv4 I__10284 (
            .O(N__43194),
            .I(\c0.n16702 ));
    InMux I__10283 (
            .O(N__43191),
            .I(N__43187));
    CascadeMux I__10282 (
            .O(N__43190),
            .I(N__43184));
    LocalMux I__10281 (
            .O(N__43187),
            .I(N__43180));
    InMux I__10280 (
            .O(N__43184),
            .I(N__43177));
    InMux I__10279 (
            .O(N__43183),
            .I(N__43174));
    Span4Mux_h I__10278 (
            .O(N__43180),
            .I(N__43171));
    LocalMux I__10277 (
            .O(N__43177),
            .I(\c0.FRAME_MATCHER_state_15 ));
    LocalMux I__10276 (
            .O(N__43174),
            .I(\c0.FRAME_MATCHER_state_15 ));
    Odrv4 I__10275 (
            .O(N__43171),
            .I(\c0.FRAME_MATCHER_state_15 ));
    SRMux I__10274 (
            .O(N__43164),
            .I(N__43161));
    LocalMux I__10273 (
            .O(N__43161),
            .I(\c0.n8_adj_2330 ));
    InMux I__10272 (
            .O(N__43158),
            .I(N__43154));
    CascadeMux I__10271 (
            .O(N__43157),
            .I(N__43151));
    LocalMux I__10270 (
            .O(N__43154),
            .I(N__43147));
    InMux I__10269 (
            .O(N__43151),
            .I(N__43144));
    InMux I__10268 (
            .O(N__43150),
            .I(N__43141));
    Span4Mux_h I__10267 (
            .O(N__43147),
            .I(N__43138));
    LocalMux I__10266 (
            .O(N__43144),
            .I(\c0.FRAME_MATCHER_state_21 ));
    LocalMux I__10265 (
            .O(N__43141),
            .I(\c0.FRAME_MATCHER_state_21 ));
    Odrv4 I__10264 (
            .O(N__43138),
            .I(\c0.FRAME_MATCHER_state_21 ));
    SRMux I__10263 (
            .O(N__43131),
            .I(N__43128));
    LocalMux I__10262 (
            .O(N__43128),
            .I(N__43125));
    Span4Mux_v I__10261 (
            .O(N__43125),
            .I(N__43122));
    Odrv4 I__10260 (
            .O(N__43122),
            .I(\c0.n16686 ));
    CascadeMux I__10259 (
            .O(N__43119),
            .I(N__43115));
    InMux I__10258 (
            .O(N__43118),
            .I(N__43111));
    InMux I__10257 (
            .O(N__43115),
            .I(N__43108));
    CascadeMux I__10256 (
            .O(N__43114),
            .I(N__43105));
    LocalMux I__10255 (
            .O(N__43111),
            .I(N__43100));
    LocalMux I__10254 (
            .O(N__43108),
            .I(N__43100));
    InMux I__10253 (
            .O(N__43105),
            .I(N__43097));
    Span4Mux_h I__10252 (
            .O(N__43100),
            .I(N__43094));
    LocalMux I__10251 (
            .O(N__43097),
            .I(\c0.FRAME_MATCHER_state_24 ));
    Odrv4 I__10250 (
            .O(N__43094),
            .I(\c0.FRAME_MATCHER_state_24 ));
    SRMux I__10249 (
            .O(N__43089),
            .I(N__43086));
    LocalMux I__10248 (
            .O(N__43086),
            .I(N__43083));
    Odrv4 I__10247 (
            .O(N__43083),
            .I(\c0.n16688 ));
    CascadeMux I__10246 (
            .O(N__43080),
            .I(\c0.n68_cascade_ ));
    InMux I__10245 (
            .O(N__43077),
            .I(N__43072));
    InMux I__10244 (
            .O(N__43076),
            .I(N__43069));
    InMux I__10243 (
            .O(N__43075),
            .I(N__43066));
    LocalMux I__10242 (
            .O(N__43072),
            .I(tx_transmit_N_1947_7));
    LocalMux I__10241 (
            .O(N__43069),
            .I(tx_transmit_N_1947_7));
    LocalMux I__10240 (
            .O(N__43066),
            .I(tx_transmit_N_1947_7));
    SRMux I__10239 (
            .O(N__43059),
            .I(N__43056));
    LocalMux I__10238 (
            .O(N__43056),
            .I(N__43053));
    Odrv4 I__10237 (
            .O(N__43053),
            .I(\c0.n4650 ));
    InMux I__10236 (
            .O(N__43050),
            .I(N__43047));
    LocalMux I__10235 (
            .O(N__43047),
            .I(N__43044));
    Span4Mux_h I__10234 (
            .O(N__43044),
            .I(N__43035));
    InMux I__10233 (
            .O(N__43043),
            .I(N__43030));
    InMux I__10232 (
            .O(N__43042),
            .I(N__43030));
    InMux I__10231 (
            .O(N__43041),
            .I(N__43027));
    InMux I__10230 (
            .O(N__43040),
            .I(N__43022));
    InMux I__10229 (
            .O(N__43039),
            .I(N__43022));
    InMux I__10228 (
            .O(N__43038),
            .I(N__43019));
    Odrv4 I__10227 (
            .O(N__43035),
            .I(tx_transmit_N_1947_3));
    LocalMux I__10226 (
            .O(N__43030),
            .I(tx_transmit_N_1947_3));
    LocalMux I__10225 (
            .O(N__43027),
            .I(tx_transmit_N_1947_3));
    LocalMux I__10224 (
            .O(N__43022),
            .I(tx_transmit_N_1947_3));
    LocalMux I__10223 (
            .O(N__43019),
            .I(tx_transmit_N_1947_3));
    InMux I__10222 (
            .O(N__43008),
            .I(N__43005));
    LocalMux I__10221 (
            .O(N__43005),
            .I(\c0.n59 ));
    CascadeMux I__10220 (
            .O(N__43002),
            .I(N__42999));
    InMux I__10219 (
            .O(N__42999),
            .I(N__42996));
    LocalMux I__10218 (
            .O(N__42996),
            .I(\c0.n65 ));
    InMux I__10217 (
            .O(N__42993),
            .I(N__42990));
    LocalMux I__10216 (
            .O(N__42990),
            .I(N__42986));
    CascadeMux I__10215 (
            .O(N__42989),
            .I(N__42982));
    Span4Mux_h I__10214 (
            .O(N__42986),
            .I(N__42979));
    InMux I__10213 (
            .O(N__42985),
            .I(N__42976));
    InMux I__10212 (
            .O(N__42982),
            .I(N__42973));
    Odrv4 I__10211 (
            .O(N__42979),
            .I(tx_transmit_N_1947_4));
    LocalMux I__10210 (
            .O(N__42976),
            .I(tx_transmit_N_1947_4));
    LocalMux I__10209 (
            .O(N__42973),
            .I(tx_transmit_N_1947_4));
    CascadeMux I__10208 (
            .O(N__42966),
            .I(N__42963));
    InMux I__10207 (
            .O(N__42963),
            .I(N__42958));
    InMux I__10206 (
            .O(N__42962),
            .I(N__42955));
    InMux I__10205 (
            .O(N__42961),
            .I(N__42952));
    LocalMux I__10204 (
            .O(N__42958),
            .I(tx_transmit_N_1947_5));
    LocalMux I__10203 (
            .O(N__42955),
            .I(tx_transmit_N_1947_5));
    LocalMux I__10202 (
            .O(N__42952),
            .I(tx_transmit_N_1947_5));
    InMux I__10201 (
            .O(N__42945),
            .I(N__42942));
    LocalMux I__10200 (
            .O(N__42942),
            .I(N__42939));
    Span4Mux_h I__10199 (
            .O(N__42939),
            .I(N__42936));
    Span4Mux_v I__10198 (
            .O(N__42936),
            .I(N__42931));
    InMux I__10197 (
            .O(N__42935),
            .I(N__42928));
    InMux I__10196 (
            .O(N__42934),
            .I(N__42925));
    Odrv4 I__10195 (
            .O(N__42931),
            .I(tx_transmit_N_1947_6));
    LocalMux I__10194 (
            .O(N__42928),
            .I(tx_transmit_N_1947_6));
    LocalMux I__10193 (
            .O(N__42925),
            .I(tx_transmit_N_1947_6));
    InMux I__10192 (
            .O(N__42918),
            .I(N__42915));
    LocalMux I__10191 (
            .O(N__42915),
            .I(\c0.n17404 ));
    InMux I__10190 (
            .O(N__42912),
            .I(N__42909));
    LocalMux I__10189 (
            .O(N__42909),
            .I(N__42906));
    Span4Mux_h I__10188 (
            .O(N__42906),
            .I(N__42902));
    InMux I__10187 (
            .O(N__42905),
            .I(N__42899));
    Odrv4 I__10186 (
            .O(N__42902),
            .I(tx_transmit_N_1947_1));
    LocalMux I__10185 (
            .O(N__42899),
            .I(tx_transmit_N_1947_1));
    InMux I__10184 (
            .O(N__42894),
            .I(N__42891));
    LocalMux I__10183 (
            .O(N__42891),
            .I(N__42888));
    Span4Mux_v I__10182 (
            .O(N__42888),
            .I(N__42884));
    InMux I__10181 (
            .O(N__42887),
            .I(N__42881));
    Odrv4 I__10180 (
            .O(N__42884),
            .I(tx_transmit_N_1947_0));
    LocalMux I__10179 (
            .O(N__42881),
            .I(tx_transmit_N_1947_0));
    InMux I__10178 (
            .O(N__42876),
            .I(N__42871));
    InMux I__10177 (
            .O(N__42875),
            .I(N__42868));
    InMux I__10176 (
            .O(N__42874),
            .I(N__42865));
    LocalMux I__10175 (
            .O(N__42871),
            .I(N__42862));
    LocalMux I__10174 (
            .O(N__42868),
            .I(\c0.n13662 ));
    LocalMux I__10173 (
            .O(N__42865),
            .I(\c0.n13662 ));
    Odrv4 I__10172 (
            .O(N__42862),
            .I(\c0.n13662 ));
    CascadeMux I__10171 (
            .O(N__42855),
            .I(\c0.n13662_cascade_ ));
    InMux I__10170 (
            .O(N__42852),
            .I(N__42849));
    LocalMux I__10169 (
            .O(N__42849),
            .I(N__42846));
    Span4Mux_h I__10168 (
            .O(N__42846),
            .I(N__42838));
    InMux I__10167 (
            .O(N__42845),
            .I(N__42835));
    InMux I__10166 (
            .O(N__42844),
            .I(N__42832));
    InMux I__10165 (
            .O(N__42843),
            .I(N__42825));
    InMux I__10164 (
            .O(N__42842),
            .I(N__42825));
    InMux I__10163 (
            .O(N__42841),
            .I(N__42825));
    Odrv4 I__10162 (
            .O(N__42838),
            .I(tx_transmit_N_1947_2));
    LocalMux I__10161 (
            .O(N__42835),
            .I(tx_transmit_N_1947_2));
    LocalMux I__10160 (
            .O(N__42832),
            .I(tx_transmit_N_1947_2));
    LocalMux I__10159 (
            .O(N__42825),
            .I(tx_transmit_N_1947_2));
    InMux I__10158 (
            .O(N__42816),
            .I(N__42813));
    LocalMux I__10157 (
            .O(N__42813),
            .I(N__42810));
    Odrv4 I__10156 (
            .O(N__42810),
            .I(\c0.n13726 ));
    SRMux I__10155 (
            .O(N__42807),
            .I(N__42803));
    SRMux I__10154 (
            .O(N__42806),
            .I(N__42800));
    LocalMux I__10153 (
            .O(N__42803),
            .I(N__42797));
    LocalMux I__10152 (
            .O(N__42800),
            .I(N__42794));
    Sp12to4 I__10151 (
            .O(N__42797),
            .I(N__42790));
    Span4Mux_h I__10150 (
            .O(N__42794),
            .I(N__42787));
    SRMux I__10149 (
            .O(N__42793),
            .I(N__42784));
    Span12Mux_s8_h I__10148 (
            .O(N__42790),
            .I(N__42781));
    Span4Mux_h I__10147 (
            .O(N__42787),
            .I(N__42778));
    LocalMux I__10146 (
            .O(N__42784),
            .I(N__42775));
    Odrv12 I__10145 (
            .O(N__42781),
            .I(\c0.n10815 ));
    Odrv4 I__10144 (
            .O(N__42778),
            .I(\c0.n10815 ));
    Odrv12 I__10143 (
            .O(N__42775),
            .I(\c0.n10815 ));
    InMux I__10142 (
            .O(N__42768),
            .I(N__42765));
    LocalMux I__10141 (
            .O(N__42765),
            .I(N__42762));
    Span4Mux_h I__10140 (
            .O(N__42762),
            .I(N__42758));
    InMux I__10139 (
            .O(N__42761),
            .I(N__42755));
    Span4Mux_v I__10138 (
            .O(N__42758),
            .I(N__42752));
    LocalMux I__10137 (
            .O(N__42755),
            .I(data_out_0_3));
    Odrv4 I__10136 (
            .O(N__42752),
            .I(data_out_0_3));
    InMux I__10135 (
            .O(N__42747),
            .I(\c0.n16110 ));
    InMux I__10134 (
            .O(N__42744),
            .I(\c0.n16111 ));
    InMux I__10133 (
            .O(N__42741),
            .I(\c0.n16112 ));
    InMux I__10132 (
            .O(N__42738),
            .I(\c0.n16113 ));
    InMux I__10131 (
            .O(N__42735),
            .I(N__42731));
    InMux I__10130 (
            .O(N__42734),
            .I(N__42728));
    LocalMux I__10129 (
            .O(N__42731),
            .I(byte_transmit_counter_5));
    LocalMux I__10128 (
            .O(N__42728),
            .I(byte_transmit_counter_5));
    InMux I__10127 (
            .O(N__42723),
            .I(\c0.n16114 ));
    InMux I__10126 (
            .O(N__42720),
            .I(N__42717));
    LocalMux I__10125 (
            .O(N__42717),
            .I(N__42713));
    InMux I__10124 (
            .O(N__42716),
            .I(N__42710));
    Span4Mux_v I__10123 (
            .O(N__42713),
            .I(N__42707));
    LocalMux I__10122 (
            .O(N__42710),
            .I(byte_transmit_counter_6));
    Odrv4 I__10121 (
            .O(N__42707),
            .I(byte_transmit_counter_6));
    InMux I__10120 (
            .O(N__42702),
            .I(\c0.n16115 ));
    InMux I__10119 (
            .O(N__42699),
            .I(N__42695));
    InMux I__10118 (
            .O(N__42698),
            .I(N__42692));
    LocalMux I__10117 (
            .O(N__42695),
            .I(byte_transmit_counter_7));
    LocalMux I__10116 (
            .O(N__42692),
            .I(byte_transmit_counter_7));
    InMux I__10115 (
            .O(N__42687),
            .I(\c0.n16116 ));
    CascadeMux I__10114 (
            .O(N__42684),
            .I(n5_adj_2448_cascade_));
    CascadeMux I__10113 (
            .O(N__42681),
            .I(n31_cascade_));
    InMux I__10112 (
            .O(N__42678),
            .I(N__42675));
    LocalMux I__10111 (
            .O(N__42675),
            .I(n22));
    InMux I__10110 (
            .O(N__42672),
            .I(N__42667));
    InMux I__10109 (
            .O(N__42671),
            .I(N__42662));
    InMux I__10108 (
            .O(N__42670),
            .I(N__42662));
    LocalMux I__10107 (
            .O(N__42667),
            .I(n9524));
    LocalMux I__10106 (
            .O(N__42662),
            .I(n9524));
    InMux I__10105 (
            .O(N__42657),
            .I(N__42650));
    InMux I__10104 (
            .O(N__42656),
            .I(N__42650));
    InMux I__10103 (
            .O(N__42655),
            .I(N__42647));
    LocalMux I__10102 (
            .O(N__42650),
            .I(n450));
    LocalMux I__10101 (
            .O(N__42647),
            .I(n450));
    InMux I__10100 (
            .O(N__42642),
            .I(N__42637));
    CascadeMux I__10099 (
            .O(N__42641),
            .I(N__42633));
    InMux I__10098 (
            .O(N__42640),
            .I(N__42630));
    LocalMux I__10097 (
            .O(N__42637),
            .I(N__42627));
    CascadeMux I__10096 (
            .O(N__42636),
            .I(N__42621));
    InMux I__10095 (
            .O(N__42633),
            .I(N__42618));
    LocalMux I__10094 (
            .O(N__42630),
            .I(N__42615));
    Span4Mux_h I__10093 (
            .O(N__42627),
            .I(N__42612));
    InMux I__10092 (
            .O(N__42626),
            .I(N__42607));
    InMux I__10091 (
            .O(N__42625),
            .I(N__42607));
    InMux I__10090 (
            .O(N__42624),
            .I(N__42602));
    InMux I__10089 (
            .O(N__42621),
            .I(N__42602));
    LocalMux I__10088 (
            .O(N__42618),
            .I(r_Bit_Index_1));
    Odrv4 I__10087 (
            .O(N__42615),
            .I(r_Bit_Index_1));
    Odrv4 I__10086 (
            .O(N__42612),
            .I(r_Bit_Index_1));
    LocalMux I__10085 (
            .O(N__42607),
            .I(r_Bit_Index_1));
    LocalMux I__10084 (
            .O(N__42602),
            .I(r_Bit_Index_1));
    CascadeMux I__10083 (
            .O(N__42591),
            .I(N__42588));
    InMux I__10082 (
            .O(N__42588),
            .I(N__42585));
    LocalMux I__10081 (
            .O(N__42585),
            .I(N__42580));
    InMux I__10080 (
            .O(N__42584),
            .I(N__42575));
    InMux I__10079 (
            .O(N__42583),
            .I(N__42572));
    Span4Mux_h I__10078 (
            .O(N__42580),
            .I(N__42569));
    InMux I__10077 (
            .O(N__42579),
            .I(N__42564));
    InMux I__10076 (
            .O(N__42578),
            .I(N__42564));
    LocalMux I__10075 (
            .O(N__42575),
            .I(\c0.tx.r_Bit_Index_0 ));
    LocalMux I__10074 (
            .O(N__42572),
            .I(\c0.tx.r_Bit_Index_0 ));
    Odrv4 I__10073 (
            .O(N__42569),
            .I(\c0.tx.r_Bit_Index_0 ));
    LocalMux I__10072 (
            .O(N__42564),
            .I(\c0.tx.r_Bit_Index_0 ));
    InMux I__10071 (
            .O(N__42555),
            .I(N__42551));
    InMux I__10070 (
            .O(N__42554),
            .I(N__42547));
    LocalMux I__10069 (
            .O(N__42551),
            .I(N__42543));
    InMux I__10068 (
            .O(N__42550),
            .I(N__42540));
    LocalMux I__10067 (
            .O(N__42547),
            .I(N__42537));
    InMux I__10066 (
            .O(N__42546),
            .I(N__42534));
    Span4Mux_h I__10065 (
            .O(N__42543),
            .I(N__42531));
    LocalMux I__10064 (
            .O(N__42540),
            .I(r_Bit_Index_2));
    Odrv4 I__10063 (
            .O(N__42537),
            .I(r_Bit_Index_2));
    LocalMux I__10062 (
            .O(N__42534),
            .I(r_Bit_Index_2));
    Odrv4 I__10061 (
            .O(N__42531),
            .I(r_Bit_Index_2));
    CascadeMux I__10060 (
            .O(N__42522),
            .I(\c0.tx.n17673_cascade_ ));
    CascadeMux I__10059 (
            .O(N__42519),
            .I(N__42515));
    InMux I__10058 (
            .O(N__42518),
            .I(N__42512));
    InMux I__10057 (
            .O(N__42515),
            .I(N__42509));
    LocalMux I__10056 (
            .O(N__42512),
            .I(N__42506));
    LocalMux I__10055 (
            .O(N__42509),
            .I(N__42503));
    Span4Mux_h I__10054 (
            .O(N__42506),
            .I(N__42500));
    Span4Mux_h I__10053 (
            .O(N__42503),
            .I(N__42497));
    Odrv4 I__10052 (
            .O(N__42500),
            .I(\c0.n10326 ));
    Odrv4 I__10051 (
            .O(N__42497),
            .I(\c0.n10326 ));
    InMux I__10050 (
            .O(N__42492),
            .I(N__42489));
    LocalMux I__10049 (
            .O(N__42489),
            .I(N__42486));
    Span4Mux_h I__10048 (
            .O(N__42486),
            .I(N__42483));
    Span4Mux_h I__10047 (
            .O(N__42483),
            .I(N__42480));
    Odrv4 I__10046 (
            .O(N__42480),
            .I(\c0.n17126 ));
    CascadeMux I__10045 (
            .O(N__42477),
            .I(\c0.n17126_cascade_ ));
    InMux I__10044 (
            .O(N__42474),
            .I(N__42471));
    LocalMux I__10043 (
            .O(N__42471),
            .I(N__42468));
    Span4Mux_h I__10042 (
            .O(N__42468),
            .I(N__42465));
    Odrv4 I__10041 (
            .O(N__42465),
            .I(\c0.n17651 ));
    CascadeMux I__10040 (
            .O(N__42462),
            .I(N__42457));
    CascadeMux I__10039 (
            .O(N__42461),
            .I(N__42453));
    InMux I__10038 (
            .O(N__42460),
            .I(N__42449));
    InMux I__10037 (
            .O(N__42457),
            .I(N__42443));
    InMux I__10036 (
            .O(N__42456),
            .I(N__42438));
    InMux I__10035 (
            .O(N__42453),
            .I(N__42438));
    CascadeMux I__10034 (
            .O(N__42452),
            .I(N__42435));
    LocalMux I__10033 (
            .O(N__42449),
            .I(N__42432));
    CascadeMux I__10032 (
            .O(N__42448),
            .I(N__42429));
    CascadeMux I__10031 (
            .O(N__42447),
            .I(N__42426));
    CascadeMux I__10030 (
            .O(N__42446),
            .I(N__42423));
    LocalMux I__10029 (
            .O(N__42443),
            .I(N__42418));
    LocalMux I__10028 (
            .O(N__42438),
            .I(N__42418));
    InMux I__10027 (
            .O(N__42435),
            .I(N__42415));
    Span4Mux_v I__10026 (
            .O(N__42432),
            .I(N__42412));
    InMux I__10025 (
            .O(N__42429),
            .I(N__42405));
    InMux I__10024 (
            .O(N__42426),
            .I(N__42405));
    InMux I__10023 (
            .O(N__42423),
            .I(N__42405));
    Span4Mux_v I__10022 (
            .O(N__42418),
            .I(N__42402));
    LocalMux I__10021 (
            .O(N__42415),
            .I(N__42399));
    Span4Mux_v I__10020 (
            .O(N__42412),
            .I(N__42396));
    LocalMux I__10019 (
            .O(N__42405),
            .I(N__42393));
    Span4Mux_v I__10018 (
            .O(N__42402),
            .I(N__42390));
    Span4Mux_h I__10017 (
            .O(N__42399),
            .I(N__42387));
    Span4Mux_h I__10016 (
            .O(N__42396),
            .I(N__42382));
    Span4Mux_v I__10015 (
            .O(N__42393),
            .I(N__42382));
    Span4Mux_h I__10014 (
            .O(N__42390),
            .I(N__42377));
    Span4Mux_v I__10013 (
            .O(N__42387),
            .I(N__42377));
    Span4Mux_v I__10012 (
            .O(N__42382),
            .I(N__42374));
    Odrv4 I__10011 (
            .O(N__42377),
            .I(n10705));
    Odrv4 I__10010 (
            .O(N__42374),
            .I(n10705));
    InMux I__10009 (
            .O(N__42369),
            .I(N__42358));
    InMux I__10008 (
            .O(N__42368),
            .I(N__42358));
    InMux I__10007 (
            .O(N__42367),
            .I(N__42358));
    InMux I__10006 (
            .O(N__42366),
            .I(N__42355));
    InMux I__10005 (
            .O(N__42365),
            .I(N__42352));
    LocalMux I__10004 (
            .O(N__42358),
            .I(N__42345));
    LocalMux I__10003 (
            .O(N__42355),
            .I(N__42345));
    LocalMux I__10002 (
            .O(N__42352),
            .I(N__42342));
    InMux I__10001 (
            .O(N__42351),
            .I(N__42339));
    InMux I__10000 (
            .O(N__42350),
            .I(N__42336));
    Odrv4 I__9999 (
            .O(N__42345),
            .I(n10_adj_2444));
    Odrv4 I__9998 (
            .O(N__42342),
            .I(n10_adj_2444));
    LocalMux I__9997 (
            .O(N__42339),
            .I(n10_adj_2444));
    LocalMux I__9996 (
            .O(N__42336),
            .I(n10_adj_2444));
    CascadeMux I__9995 (
            .O(N__42327),
            .I(n18187_cascade_));
    InMux I__9994 (
            .O(N__42324),
            .I(N__42320));
    InMux I__9993 (
            .O(N__42323),
            .I(N__42317));
    LocalMux I__9992 (
            .O(N__42320),
            .I(N__42312));
    LocalMux I__9991 (
            .O(N__42317),
            .I(N__42312));
    Odrv4 I__9990 (
            .O(N__42312),
            .I(\c0.data_out_6_6 ));
    CascadeMux I__9989 (
            .O(N__42309),
            .I(N__42306));
    InMux I__9988 (
            .O(N__42306),
            .I(N__42303));
    LocalMux I__9987 (
            .O(N__42303),
            .I(\c0.n5_adj_2159 ));
    InMux I__9986 (
            .O(N__42300),
            .I(N__42297));
    LocalMux I__9985 (
            .O(N__42297),
            .I(N__42294));
    Span4Mux_h I__9984 (
            .O(N__42294),
            .I(N__42290));
    CascadeMux I__9983 (
            .O(N__42293),
            .I(N__42287));
    Span4Mux_h I__9982 (
            .O(N__42290),
            .I(N__42284));
    InMux I__9981 (
            .O(N__42287),
            .I(N__42281));
    Odrv4 I__9980 (
            .O(N__42284),
            .I(rand_setpoint_30));
    LocalMux I__9979 (
            .O(N__42281),
            .I(rand_setpoint_30));
    InMux I__9978 (
            .O(N__42276),
            .I(N__42273));
    LocalMux I__9977 (
            .O(N__42273),
            .I(\c0.n17698 ));
    InMux I__9976 (
            .O(N__42270),
            .I(N__42267));
    LocalMux I__9975 (
            .O(N__42267),
            .I(\c0.n17612 ));
    CascadeMux I__9974 (
            .O(N__42264),
            .I(N__42261));
    InMux I__9973 (
            .O(N__42261),
            .I(N__42258));
    LocalMux I__9972 (
            .O(N__42258),
            .I(N__42255));
    Span4Mux_v I__9971 (
            .O(N__42255),
            .I(N__42252));
    Span4Mux_h I__9970 (
            .O(N__42252),
            .I(N__42249));
    Odrv4 I__9969 (
            .O(N__42249),
            .I(\c0.n17626 ));
    CascadeMux I__9968 (
            .O(N__42246),
            .I(N__42243));
    InMux I__9967 (
            .O(N__42243),
            .I(N__42240));
    LocalMux I__9966 (
            .O(N__42240),
            .I(N__42237));
    Span4Mux_h I__9965 (
            .O(N__42237),
            .I(N__42234));
    Odrv4 I__9964 (
            .O(N__42234),
            .I(n25));
    InMux I__9963 (
            .O(N__42231),
            .I(N__42228));
    LocalMux I__9962 (
            .O(N__42228),
            .I(N__42225));
    Odrv4 I__9961 (
            .O(N__42225),
            .I(n28));
    SRMux I__9960 (
            .O(N__42222),
            .I(N__42219));
    LocalMux I__9959 (
            .O(N__42219),
            .I(\c0.n16704 ));
    InMux I__9958 (
            .O(N__42216),
            .I(N__42213));
    LocalMux I__9957 (
            .O(N__42213),
            .I(N__42210));
    Odrv4 I__9956 (
            .O(N__42210),
            .I(\c0.n3_adj_2193 ));
    CascadeMux I__9955 (
            .O(N__42207),
            .I(N__42204));
    InMux I__9954 (
            .O(N__42204),
            .I(N__42201));
    LocalMux I__9953 (
            .O(N__42201),
            .I(N__42198));
    Span4Mux_h I__9952 (
            .O(N__42198),
            .I(N__42195));
    Odrv4 I__9951 (
            .O(N__42195),
            .I(n10_adj_2431));
    InMux I__9950 (
            .O(N__42192),
            .I(N__42189));
    LocalMux I__9949 (
            .O(N__42189),
            .I(N__42186));
    Span4Mux_v I__9948 (
            .O(N__42186),
            .I(N__42183));
    Span4Mux_h I__9947 (
            .O(N__42183),
            .I(N__42180));
    Odrv4 I__9946 (
            .O(N__42180),
            .I(\c0.n6_adj_2221 ));
    InMux I__9945 (
            .O(N__42177),
            .I(N__42171));
    InMux I__9944 (
            .O(N__42176),
            .I(N__42171));
    LocalMux I__9943 (
            .O(N__42171),
            .I(\c0.n17147 ));
    InMux I__9942 (
            .O(N__42168),
            .I(N__42164));
    CascadeMux I__9941 (
            .O(N__42167),
            .I(N__42161));
    LocalMux I__9940 (
            .O(N__42164),
            .I(N__42158));
    InMux I__9939 (
            .O(N__42161),
            .I(N__42155));
    Odrv12 I__9938 (
            .O(N__42158),
            .I(rand_setpoint_8));
    LocalMux I__9937 (
            .O(N__42155),
            .I(rand_setpoint_8));
    InMux I__9936 (
            .O(N__42150),
            .I(N__42147));
    LocalMux I__9935 (
            .O(N__42147),
            .I(\c0.n17653 ));
    InMux I__9934 (
            .O(N__42144),
            .I(N__42140));
    InMux I__9933 (
            .O(N__42143),
            .I(N__42137));
    LocalMux I__9932 (
            .O(N__42140),
            .I(N__42133));
    LocalMux I__9931 (
            .O(N__42137),
            .I(N__42130));
    InMux I__9930 (
            .O(N__42136),
            .I(N__42126));
    Span4Mux_h I__9929 (
            .O(N__42133),
            .I(N__42123));
    Span4Mux_v I__9928 (
            .O(N__42130),
            .I(N__42120));
    InMux I__9927 (
            .O(N__42129),
            .I(N__42117));
    LocalMux I__9926 (
            .O(N__42126),
            .I(data_out_8_1));
    Odrv4 I__9925 (
            .O(N__42123),
            .I(data_out_8_1));
    Odrv4 I__9924 (
            .O(N__42120),
            .I(data_out_8_1));
    LocalMux I__9923 (
            .O(N__42117),
            .I(data_out_8_1));
    InMux I__9922 (
            .O(N__42108),
            .I(N__42105));
    LocalMux I__9921 (
            .O(N__42105),
            .I(N__42102));
    Odrv12 I__9920 (
            .O(N__42102),
            .I(\c0.n1_adj_2160 ));
    CascadeMux I__9919 (
            .O(N__42099),
            .I(\c0.n18184_cascade_ ));
    InMux I__9918 (
            .O(N__42096),
            .I(N__42090));
    InMux I__9917 (
            .O(N__42095),
            .I(N__42087));
    InMux I__9916 (
            .O(N__42094),
            .I(N__42081));
    InMux I__9915 (
            .O(N__42093),
            .I(N__42078));
    LocalMux I__9914 (
            .O(N__42090),
            .I(N__42075));
    LocalMux I__9913 (
            .O(N__42087),
            .I(N__42072));
    InMux I__9912 (
            .O(N__42086),
            .I(N__42069));
    InMux I__9911 (
            .O(N__42085),
            .I(N__42066));
    InMux I__9910 (
            .O(N__42084),
            .I(N__42063));
    LocalMux I__9909 (
            .O(N__42081),
            .I(N__42060));
    LocalMux I__9908 (
            .O(N__42078),
            .I(N__42057));
    Span4Mux_v I__9907 (
            .O(N__42075),
            .I(N__42054));
    Span4Mux_v I__9906 (
            .O(N__42072),
            .I(N__42050));
    LocalMux I__9905 (
            .O(N__42069),
            .I(N__42047));
    LocalMux I__9904 (
            .O(N__42066),
            .I(N__42044));
    LocalMux I__9903 (
            .O(N__42063),
            .I(N__42041));
    Span4Mux_h I__9902 (
            .O(N__42060),
            .I(N__42035));
    Span4Mux_h I__9901 (
            .O(N__42057),
            .I(N__42035));
    Sp12to4 I__9900 (
            .O(N__42054),
            .I(N__42032));
    InMux I__9899 (
            .O(N__42053),
            .I(N__42029));
    Span4Mux_h I__9898 (
            .O(N__42050),
            .I(N__42024));
    Span4Mux_v I__9897 (
            .O(N__42047),
            .I(N__42024));
    Span4Mux_v I__9896 (
            .O(N__42044),
            .I(N__42019));
    Span4Mux_h I__9895 (
            .O(N__42041),
            .I(N__42019));
    InMux I__9894 (
            .O(N__42040),
            .I(N__42016));
    Span4Mux_v I__9893 (
            .O(N__42035),
            .I(N__42011));
    Span12Mux_h I__9892 (
            .O(N__42032),
            .I(N__42006));
    LocalMux I__9891 (
            .O(N__42029),
            .I(N__42006));
    Span4Mux_h I__9890 (
            .O(N__42024),
            .I(N__42003));
    Span4Mux_v I__9889 (
            .O(N__42019),
            .I(N__42000));
    LocalMux I__9888 (
            .O(N__42016),
            .I(N__41997));
    InMux I__9887 (
            .O(N__42015),
            .I(N__41994));
    InMux I__9886 (
            .O(N__42014),
            .I(N__41991));
    Odrv4 I__9885 (
            .O(N__42011),
            .I(FRAME_MATCHER_i_31__N_1272));
    Odrv12 I__9884 (
            .O(N__42006),
            .I(FRAME_MATCHER_i_31__N_1272));
    Odrv4 I__9883 (
            .O(N__42003),
            .I(FRAME_MATCHER_i_31__N_1272));
    Odrv4 I__9882 (
            .O(N__42000),
            .I(FRAME_MATCHER_i_31__N_1272));
    Odrv4 I__9881 (
            .O(N__41997),
            .I(FRAME_MATCHER_i_31__N_1272));
    LocalMux I__9880 (
            .O(N__41994),
            .I(FRAME_MATCHER_i_31__N_1272));
    LocalMux I__9879 (
            .O(N__41991),
            .I(FRAME_MATCHER_i_31__N_1272));
    CascadeMux I__9878 (
            .O(N__41976),
            .I(N__41973));
    InMux I__9877 (
            .O(N__41973),
            .I(N__41969));
    InMux I__9876 (
            .O(N__41972),
            .I(N__41964));
    LocalMux I__9875 (
            .O(N__41969),
            .I(N__41961));
    InMux I__9874 (
            .O(N__41968),
            .I(N__41958));
    InMux I__9873 (
            .O(N__41967),
            .I(N__41953));
    LocalMux I__9872 (
            .O(N__41964),
            .I(N__41950));
    Span4Mux_h I__9871 (
            .O(N__41961),
            .I(N__41947));
    LocalMux I__9870 (
            .O(N__41958),
            .I(N__41943));
    InMux I__9869 (
            .O(N__41957),
            .I(N__41938));
    InMux I__9868 (
            .O(N__41956),
            .I(N__41938));
    LocalMux I__9867 (
            .O(N__41953),
            .I(N__41935));
    Span4Mux_v I__9866 (
            .O(N__41950),
            .I(N__41932));
    Span4Mux_v I__9865 (
            .O(N__41947),
            .I(N__41929));
    InMux I__9864 (
            .O(N__41946),
            .I(N__41926));
    Span4Mux_h I__9863 (
            .O(N__41943),
            .I(N__41919));
    LocalMux I__9862 (
            .O(N__41938),
            .I(N__41919));
    Span4Mux_v I__9861 (
            .O(N__41935),
            .I(N__41919));
    Span4Mux_v I__9860 (
            .O(N__41932),
            .I(N__41916));
    Odrv4 I__9859 (
            .O(N__41929),
            .I(n488));
    LocalMux I__9858 (
            .O(N__41926),
            .I(n488));
    Odrv4 I__9857 (
            .O(N__41919),
            .I(n488));
    Odrv4 I__9856 (
            .O(N__41916),
            .I(n488));
    InMux I__9855 (
            .O(N__41907),
            .I(N__41892));
    InMux I__9854 (
            .O(N__41906),
            .I(N__41892));
    InMux I__9853 (
            .O(N__41905),
            .I(N__41892));
    InMux I__9852 (
            .O(N__41904),
            .I(N__41892));
    InMux I__9851 (
            .O(N__41903),
            .I(N__41892));
    LocalMux I__9850 (
            .O(N__41892),
            .I(N__41855));
    InMux I__9849 (
            .O(N__41891),
            .I(N__41825));
    InMux I__9848 (
            .O(N__41890),
            .I(N__41825));
    InMux I__9847 (
            .O(N__41889),
            .I(N__41825));
    InMux I__9846 (
            .O(N__41888),
            .I(N__41825));
    InMux I__9845 (
            .O(N__41887),
            .I(N__41825));
    InMux I__9844 (
            .O(N__41886),
            .I(N__41814));
    InMux I__9843 (
            .O(N__41885),
            .I(N__41814));
    InMux I__9842 (
            .O(N__41884),
            .I(N__41814));
    InMux I__9841 (
            .O(N__41883),
            .I(N__41814));
    InMux I__9840 (
            .O(N__41882),
            .I(N__41814));
    InMux I__9839 (
            .O(N__41881),
            .I(N__41801));
    InMux I__9838 (
            .O(N__41880),
            .I(N__41801));
    InMux I__9837 (
            .O(N__41879),
            .I(N__41801));
    InMux I__9836 (
            .O(N__41878),
            .I(N__41801));
    InMux I__9835 (
            .O(N__41877),
            .I(N__41801));
    InMux I__9834 (
            .O(N__41876),
            .I(N__41801));
    InMux I__9833 (
            .O(N__41875),
            .I(N__41794));
    InMux I__9832 (
            .O(N__41874),
            .I(N__41794));
    InMux I__9831 (
            .O(N__41873),
            .I(N__41794));
    InMux I__9830 (
            .O(N__41872),
            .I(N__41779));
    InMux I__9829 (
            .O(N__41871),
            .I(N__41779));
    InMux I__9828 (
            .O(N__41870),
            .I(N__41779));
    InMux I__9827 (
            .O(N__41869),
            .I(N__41779));
    InMux I__9826 (
            .O(N__41868),
            .I(N__41779));
    InMux I__9825 (
            .O(N__41867),
            .I(N__41779));
    InMux I__9824 (
            .O(N__41866),
            .I(N__41779));
    InMux I__9823 (
            .O(N__41865),
            .I(N__41766));
    InMux I__9822 (
            .O(N__41864),
            .I(N__41766));
    InMux I__9821 (
            .O(N__41863),
            .I(N__41766));
    InMux I__9820 (
            .O(N__41862),
            .I(N__41766));
    InMux I__9819 (
            .O(N__41861),
            .I(N__41766));
    InMux I__9818 (
            .O(N__41860),
            .I(N__41766));
    InMux I__9817 (
            .O(N__41859),
            .I(N__41760));
    InMux I__9816 (
            .O(N__41858),
            .I(N__41760));
    Span4Mux_v I__9815 (
            .O(N__41855),
            .I(N__41757));
    InMux I__9814 (
            .O(N__41854),
            .I(N__41742));
    InMux I__9813 (
            .O(N__41853),
            .I(N__41742));
    InMux I__9812 (
            .O(N__41852),
            .I(N__41742));
    InMux I__9811 (
            .O(N__41851),
            .I(N__41742));
    InMux I__9810 (
            .O(N__41850),
            .I(N__41742));
    InMux I__9809 (
            .O(N__41849),
            .I(N__41742));
    InMux I__9808 (
            .O(N__41848),
            .I(N__41742));
    InMux I__9807 (
            .O(N__41847),
            .I(N__41730));
    InMux I__9806 (
            .O(N__41846),
            .I(N__41730));
    InMux I__9805 (
            .O(N__41845),
            .I(N__41730));
    InMux I__9804 (
            .O(N__41844),
            .I(N__41730));
    InMux I__9803 (
            .O(N__41843),
            .I(N__41730));
    InMux I__9802 (
            .O(N__41842),
            .I(N__41715));
    InMux I__9801 (
            .O(N__41841),
            .I(N__41715));
    InMux I__9800 (
            .O(N__41840),
            .I(N__41715));
    InMux I__9799 (
            .O(N__41839),
            .I(N__41715));
    InMux I__9798 (
            .O(N__41838),
            .I(N__41715));
    InMux I__9797 (
            .O(N__41837),
            .I(N__41715));
    InMux I__9796 (
            .O(N__41836),
            .I(N__41715));
    LocalMux I__9795 (
            .O(N__41825),
            .I(N__41704));
    LocalMux I__9794 (
            .O(N__41814),
            .I(N__41704));
    LocalMux I__9793 (
            .O(N__41801),
            .I(N__41704));
    LocalMux I__9792 (
            .O(N__41794),
            .I(N__41704));
    LocalMux I__9791 (
            .O(N__41779),
            .I(N__41704));
    LocalMux I__9790 (
            .O(N__41766),
            .I(N__41701));
    InMux I__9789 (
            .O(N__41765),
            .I(N__41697));
    LocalMux I__9788 (
            .O(N__41760),
            .I(N__41694));
    Span4Mux_h I__9787 (
            .O(N__41757),
            .I(N__41689));
    LocalMux I__9786 (
            .O(N__41742),
            .I(N__41689));
    InMux I__9785 (
            .O(N__41741),
            .I(N__41686));
    LocalMux I__9784 (
            .O(N__41730),
            .I(N__41683));
    LocalMux I__9783 (
            .O(N__41715),
            .I(N__41676));
    Span4Mux_v I__9782 (
            .O(N__41704),
            .I(N__41676));
    Span4Mux_h I__9781 (
            .O(N__41701),
            .I(N__41676));
    InMux I__9780 (
            .O(N__41700),
            .I(N__41665));
    LocalMux I__9779 (
            .O(N__41697),
            .I(N__41662));
    Span4Mux_h I__9778 (
            .O(N__41694),
            .I(N__41657));
    Span4Mux_v I__9777 (
            .O(N__41689),
            .I(N__41657));
    LocalMux I__9776 (
            .O(N__41686),
            .I(N__41654));
    Span4Mux_v I__9775 (
            .O(N__41683),
            .I(N__41649));
    Span4Mux_h I__9774 (
            .O(N__41676),
            .I(N__41649));
    InMux I__9773 (
            .O(N__41675),
            .I(N__41636));
    InMux I__9772 (
            .O(N__41674),
            .I(N__41636));
    InMux I__9771 (
            .O(N__41673),
            .I(N__41636));
    InMux I__9770 (
            .O(N__41672),
            .I(N__41636));
    InMux I__9769 (
            .O(N__41671),
            .I(N__41636));
    InMux I__9768 (
            .O(N__41670),
            .I(N__41636));
    InMux I__9767 (
            .O(N__41669),
            .I(N__41633));
    InMux I__9766 (
            .O(N__41668),
            .I(N__41630));
    LocalMux I__9765 (
            .O(N__41665),
            .I(\c0.n13146 ));
    Odrv4 I__9764 (
            .O(N__41662),
            .I(\c0.n13146 ));
    Odrv4 I__9763 (
            .O(N__41657),
            .I(\c0.n13146 ));
    Odrv4 I__9762 (
            .O(N__41654),
            .I(\c0.n13146 ));
    Odrv4 I__9761 (
            .O(N__41649),
            .I(\c0.n13146 ));
    LocalMux I__9760 (
            .O(N__41636),
            .I(\c0.n13146 ));
    LocalMux I__9759 (
            .O(N__41633),
            .I(\c0.n13146 ));
    LocalMux I__9758 (
            .O(N__41630),
            .I(\c0.n13146 ));
    CascadeMux I__9757 (
            .O(N__41613),
            .I(N__41610));
    InMux I__9756 (
            .O(N__41610),
            .I(N__41607));
    LocalMux I__9755 (
            .O(N__41607),
            .I(N__41602));
    InMux I__9754 (
            .O(N__41606),
            .I(N__41599));
    InMux I__9753 (
            .O(N__41605),
            .I(N__41596));
    Span4Mux_v I__9752 (
            .O(N__41602),
            .I(N__41593));
    LocalMux I__9751 (
            .O(N__41599),
            .I(N__41589));
    LocalMux I__9750 (
            .O(N__41596),
            .I(N__41586));
    Span4Mux_h I__9749 (
            .O(N__41593),
            .I(N__41583));
    InMux I__9748 (
            .O(N__41592),
            .I(N__41580));
    Span4Mux_v I__9747 (
            .O(N__41589),
            .I(N__41577));
    Sp12to4 I__9746 (
            .O(N__41586),
            .I(N__41570));
    Sp12to4 I__9745 (
            .O(N__41583),
            .I(N__41570));
    LocalMux I__9744 (
            .O(N__41580),
            .I(N__41570));
    Span4Mux_h I__9743 (
            .O(N__41577),
            .I(N__41567));
    Span12Mux_h I__9742 (
            .O(N__41570),
            .I(N__41564));
    Odrv4 I__9741 (
            .O(N__41567),
            .I(n4408));
    Odrv12 I__9740 (
            .O(N__41564),
            .I(n4408));
    CascadeMux I__9739 (
            .O(N__41559),
            .I(\c0.n276_cascade_ ));
    InMux I__9738 (
            .O(N__41556),
            .I(N__41553));
    LocalMux I__9737 (
            .O(N__41553),
            .I(N__41549));
    InMux I__9736 (
            .O(N__41552),
            .I(N__41546));
    Span12Mux_h I__9735 (
            .O(N__41549),
            .I(N__41542));
    LocalMux I__9734 (
            .O(N__41546),
            .I(N__41539));
    InMux I__9733 (
            .O(N__41545),
            .I(N__41536));
    Odrv12 I__9732 (
            .O(N__41542),
            .I(\c0.n4_adj_2135 ));
    Odrv4 I__9731 (
            .O(N__41539),
            .I(\c0.n4_adj_2135 ));
    LocalMux I__9730 (
            .O(N__41536),
            .I(\c0.n4_adj_2135 ));
    CascadeMux I__9729 (
            .O(N__41529),
            .I(\c0.n4_adj_2135_cascade_ ));
    InMux I__9728 (
            .O(N__41526),
            .I(N__41519));
    InMux I__9727 (
            .O(N__41525),
            .I(N__41519));
    InMux I__9726 (
            .O(N__41524),
            .I(N__41516));
    LocalMux I__9725 (
            .O(N__41519),
            .I(\c0.FRAME_MATCHER_state_31 ));
    LocalMux I__9724 (
            .O(N__41516),
            .I(\c0.FRAME_MATCHER_state_31 ));
    SRMux I__9723 (
            .O(N__41511),
            .I(N__41508));
    LocalMux I__9722 (
            .O(N__41508),
            .I(N__41505));
    Span4Mux_h I__9721 (
            .O(N__41505),
            .I(N__41502));
    Odrv4 I__9720 (
            .O(N__41502),
            .I(\c0.n16700 ));
    CascadeMux I__9719 (
            .O(N__41499),
            .I(N__41495));
    InMux I__9718 (
            .O(N__41498),
            .I(N__41482));
    InMux I__9717 (
            .O(N__41495),
            .I(N__41482));
    InMux I__9716 (
            .O(N__41494),
            .I(N__41482));
    InMux I__9715 (
            .O(N__41493),
            .I(N__41482));
    CascadeMux I__9714 (
            .O(N__41492),
            .I(N__41479));
    CascadeMux I__9713 (
            .O(N__41491),
            .I(N__41475));
    LocalMux I__9712 (
            .O(N__41482),
            .I(N__41469));
    InMux I__9711 (
            .O(N__41479),
            .I(N__41458));
    InMux I__9710 (
            .O(N__41478),
            .I(N__41458));
    InMux I__9709 (
            .O(N__41475),
            .I(N__41458));
    InMux I__9708 (
            .O(N__41474),
            .I(N__41458));
    InMux I__9707 (
            .O(N__41473),
            .I(N__41458));
    InMux I__9706 (
            .O(N__41472),
            .I(N__41454));
    Span4Mux_h I__9705 (
            .O(N__41469),
            .I(N__41449));
    LocalMux I__9704 (
            .O(N__41458),
            .I(N__41449));
    InMux I__9703 (
            .O(N__41457),
            .I(N__41446));
    LocalMux I__9702 (
            .O(N__41454),
            .I(N__41442));
    Span4Mux_h I__9701 (
            .O(N__41449),
            .I(N__41437));
    LocalMux I__9700 (
            .O(N__41446),
            .I(N__41437));
    InMux I__9699 (
            .O(N__41445),
            .I(N__41434));
    Odrv4 I__9698 (
            .O(N__41442),
            .I(\c0.n9334 ));
    Odrv4 I__9697 (
            .O(N__41437),
            .I(\c0.n9334 ));
    LocalMux I__9696 (
            .O(N__41434),
            .I(\c0.n9334 ));
    CascadeMux I__9695 (
            .O(N__41427),
            .I(N__41424));
    InMux I__9694 (
            .O(N__41424),
            .I(N__41414));
    CascadeMux I__9693 (
            .O(N__41423),
            .I(N__41411));
    CascadeMux I__9692 (
            .O(N__41422),
            .I(N__41408));
    CascadeMux I__9691 (
            .O(N__41421),
            .I(N__41404));
    CascadeMux I__9690 (
            .O(N__41420),
            .I(N__41401));
    CascadeMux I__9689 (
            .O(N__41419),
            .I(N__41397));
    CascadeMux I__9688 (
            .O(N__41418),
            .I(N__41393));
    CascadeMux I__9687 (
            .O(N__41417),
            .I(N__41390));
    LocalMux I__9686 (
            .O(N__41414),
            .I(N__41386));
    InMux I__9685 (
            .O(N__41411),
            .I(N__41383));
    InMux I__9684 (
            .O(N__41408),
            .I(N__41374));
    InMux I__9683 (
            .O(N__41407),
            .I(N__41374));
    InMux I__9682 (
            .O(N__41404),
            .I(N__41374));
    InMux I__9681 (
            .O(N__41401),
            .I(N__41374));
    InMux I__9680 (
            .O(N__41400),
            .I(N__41363));
    InMux I__9679 (
            .O(N__41397),
            .I(N__41363));
    InMux I__9678 (
            .O(N__41396),
            .I(N__41363));
    InMux I__9677 (
            .O(N__41393),
            .I(N__41363));
    InMux I__9676 (
            .O(N__41390),
            .I(N__41363));
    InMux I__9675 (
            .O(N__41389),
            .I(N__41359));
    Span4Mux_h I__9674 (
            .O(N__41386),
            .I(N__41354));
    LocalMux I__9673 (
            .O(N__41383),
            .I(N__41354));
    LocalMux I__9672 (
            .O(N__41374),
            .I(N__41349));
    LocalMux I__9671 (
            .O(N__41363),
            .I(N__41349));
    InMux I__9670 (
            .O(N__41362),
            .I(N__41346));
    LocalMux I__9669 (
            .O(N__41359),
            .I(n44));
    Odrv4 I__9668 (
            .O(N__41354),
            .I(n44));
    Odrv4 I__9667 (
            .O(N__41349),
            .I(n44));
    LocalMux I__9666 (
            .O(N__41346),
            .I(n44));
    InMux I__9665 (
            .O(N__41337),
            .I(N__41323));
    InMux I__9664 (
            .O(N__41336),
            .I(N__41323));
    InMux I__9663 (
            .O(N__41335),
            .I(N__41323));
    InMux I__9662 (
            .O(N__41334),
            .I(N__41323));
    InMux I__9661 (
            .O(N__41333),
            .I(N__41315));
    InMux I__9660 (
            .O(N__41332),
            .I(N__41312));
    LocalMux I__9659 (
            .O(N__41323),
            .I(N__41309));
    InMux I__9658 (
            .O(N__41322),
            .I(N__41298));
    InMux I__9657 (
            .O(N__41321),
            .I(N__41298));
    InMux I__9656 (
            .O(N__41320),
            .I(N__41298));
    InMux I__9655 (
            .O(N__41319),
            .I(N__41298));
    InMux I__9654 (
            .O(N__41318),
            .I(N__41298));
    LocalMux I__9653 (
            .O(N__41315),
            .I(N__41293));
    LocalMux I__9652 (
            .O(N__41312),
            .I(N__41290));
    Span4Mux_h I__9651 (
            .O(N__41309),
            .I(N__41285));
    LocalMux I__9650 (
            .O(N__41298),
            .I(N__41285));
    InMux I__9649 (
            .O(N__41297),
            .I(N__41282));
    InMux I__9648 (
            .O(N__41296),
            .I(N__41279));
    Odrv4 I__9647 (
            .O(N__41293),
            .I(\c0.n17069 ));
    Odrv4 I__9646 (
            .O(N__41290),
            .I(\c0.n17069 ));
    Odrv4 I__9645 (
            .O(N__41285),
            .I(\c0.n17069 ));
    LocalMux I__9644 (
            .O(N__41282),
            .I(\c0.n17069 ));
    LocalMux I__9643 (
            .O(N__41279),
            .I(\c0.n17069 ));
    InMux I__9642 (
            .O(N__41268),
            .I(N__41265));
    LocalMux I__9641 (
            .O(N__41265),
            .I(N__41260));
    CascadeMux I__9640 (
            .O(N__41264),
            .I(N__41257));
    InMux I__9639 (
            .O(N__41263),
            .I(N__41254));
    Span4Mux_v I__9638 (
            .O(N__41260),
            .I(N__41251));
    InMux I__9637 (
            .O(N__41257),
            .I(N__41248));
    LocalMux I__9636 (
            .O(N__41254),
            .I(N__41245));
    Span4Mux_h I__9635 (
            .O(N__41251),
            .I(N__41242));
    LocalMux I__9634 (
            .O(N__41248),
            .I(\c0.FRAME_MATCHER_state_17 ));
    Odrv4 I__9633 (
            .O(N__41245),
            .I(\c0.FRAME_MATCHER_state_17 ));
    Odrv4 I__9632 (
            .O(N__41242),
            .I(\c0.FRAME_MATCHER_state_17 ));
    CascadeMux I__9631 (
            .O(N__41235),
            .I(N__41232));
    InMux I__9630 (
            .O(N__41232),
            .I(N__41229));
    LocalMux I__9629 (
            .O(N__41229),
            .I(N__41224));
    InMux I__9628 (
            .O(N__41228),
            .I(N__41221));
    InMux I__9627 (
            .O(N__41227),
            .I(N__41218));
    Span4Mux_h I__9626 (
            .O(N__41224),
            .I(N__41215));
    LocalMux I__9625 (
            .O(N__41221),
            .I(\c0.FRAME_MATCHER_state_29 ));
    LocalMux I__9624 (
            .O(N__41218),
            .I(\c0.FRAME_MATCHER_state_29 ));
    Odrv4 I__9623 (
            .O(N__41215),
            .I(\c0.FRAME_MATCHER_state_29 ));
    SRMux I__9622 (
            .O(N__41208),
            .I(N__41205));
    LocalMux I__9621 (
            .O(N__41205),
            .I(N__41202));
    Span4Mux_v I__9620 (
            .O(N__41202),
            .I(N__41199));
    Span4Mux_h I__9619 (
            .O(N__41199),
            .I(N__41196));
    Odrv4 I__9618 (
            .O(N__41196),
            .I(\c0.n16658 ));
    CascadeMux I__9617 (
            .O(N__41193),
            .I(N__41189));
    CascadeMux I__9616 (
            .O(N__41192),
            .I(N__41185));
    InMux I__9615 (
            .O(N__41189),
            .I(N__41182));
    InMux I__9614 (
            .O(N__41188),
            .I(N__41179));
    InMux I__9613 (
            .O(N__41185),
            .I(N__41176));
    LocalMux I__9612 (
            .O(N__41182),
            .I(\c0.FRAME_MATCHER_state_10 ));
    LocalMux I__9611 (
            .O(N__41179),
            .I(\c0.FRAME_MATCHER_state_10 ));
    LocalMux I__9610 (
            .O(N__41176),
            .I(\c0.FRAME_MATCHER_state_10 ));
    SRMux I__9609 (
            .O(N__41169),
            .I(N__41166));
    LocalMux I__9608 (
            .O(N__41166),
            .I(N__41163));
    Span4Mux_h I__9607 (
            .O(N__41163),
            .I(N__41160));
    Odrv4 I__9606 (
            .O(N__41160),
            .I(\c0.n16710 ));
    CascadeMux I__9605 (
            .O(N__41157),
            .I(N__41153));
    InMux I__9604 (
            .O(N__41156),
            .I(N__41150));
    InMux I__9603 (
            .O(N__41153),
            .I(N__41146));
    LocalMux I__9602 (
            .O(N__41150),
            .I(N__41141));
    InMux I__9601 (
            .O(N__41149),
            .I(N__41138));
    LocalMux I__9600 (
            .O(N__41146),
            .I(N__41135));
    InMux I__9599 (
            .O(N__41145),
            .I(N__41132));
    InMux I__9598 (
            .O(N__41144),
            .I(N__41129));
    Span4Mux_h I__9597 (
            .O(N__41141),
            .I(N__41126));
    LocalMux I__9596 (
            .O(N__41138),
            .I(N__41123));
    Span12Mux_v I__9595 (
            .O(N__41135),
            .I(N__41118));
    LocalMux I__9594 (
            .O(N__41132),
            .I(N__41118));
    LocalMux I__9593 (
            .O(N__41129),
            .I(data_out_frame2_13_4));
    Odrv4 I__9592 (
            .O(N__41126),
            .I(data_out_frame2_13_4));
    Odrv12 I__9591 (
            .O(N__41123),
            .I(data_out_frame2_13_4));
    Odrv12 I__9590 (
            .O(N__41118),
            .I(data_out_frame2_13_4));
    InMux I__9589 (
            .O(N__41109),
            .I(N__41102));
    InMux I__9588 (
            .O(N__41108),
            .I(N__41099));
    InMux I__9587 (
            .O(N__41107),
            .I(N__41093));
    InMux I__9586 (
            .O(N__41106),
            .I(N__41093));
    CascadeMux I__9585 (
            .O(N__41105),
            .I(N__41090));
    LocalMux I__9584 (
            .O(N__41102),
            .I(N__41087));
    LocalMux I__9583 (
            .O(N__41099),
            .I(N__41084));
    InMux I__9582 (
            .O(N__41098),
            .I(N__41081));
    LocalMux I__9581 (
            .O(N__41093),
            .I(N__41078));
    InMux I__9580 (
            .O(N__41090),
            .I(N__41075));
    Span4Mux_h I__9579 (
            .O(N__41087),
            .I(N__41072));
    Span4Mux_v I__9578 (
            .O(N__41084),
            .I(N__41065));
    LocalMux I__9577 (
            .O(N__41081),
            .I(N__41065));
    Span4Mux_v I__9576 (
            .O(N__41078),
            .I(N__41065));
    LocalMux I__9575 (
            .O(N__41075),
            .I(N__41060));
    Span4Mux_h I__9574 (
            .O(N__41072),
            .I(N__41060));
    Odrv4 I__9573 (
            .O(N__41065),
            .I(data_out_frame2_9_0));
    Odrv4 I__9572 (
            .O(N__41060),
            .I(data_out_frame2_9_0));
    CascadeMux I__9571 (
            .O(N__41055),
            .I(N__41052));
    InMux I__9570 (
            .O(N__41052),
            .I(N__41049));
    LocalMux I__9569 (
            .O(N__41049),
            .I(N__41046));
    Span4Mux_v I__9568 (
            .O(N__41046),
            .I(N__41043));
    Span4Mux_h I__9567 (
            .O(N__41043),
            .I(N__41040));
    Span4Mux_h I__9566 (
            .O(N__41040),
            .I(N__41037));
    Odrv4 I__9565 (
            .O(N__41037),
            .I(\c0.n17315 ));
    CascadeMux I__9564 (
            .O(N__41034),
            .I(N__41027));
    InMux I__9563 (
            .O(N__41033),
            .I(N__41024));
    InMux I__9562 (
            .O(N__41032),
            .I(N__41021));
    InMux I__9561 (
            .O(N__41031),
            .I(N__41018));
    InMux I__9560 (
            .O(N__41030),
            .I(N__41015));
    InMux I__9559 (
            .O(N__41027),
            .I(N__41012));
    LocalMux I__9558 (
            .O(N__41024),
            .I(N__41009));
    LocalMux I__9557 (
            .O(N__41021),
            .I(N__41006));
    LocalMux I__9556 (
            .O(N__41018),
            .I(N__41003));
    LocalMux I__9555 (
            .O(N__41015),
            .I(N__41000));
    LocalMux I__9554 (
            .O(N__41012),
            .I(\c0.data_in_frame_0_0 ));
    Odrv12 I__9553 (
            .O(N__41009),
            .I(\c0.data_in_frame_0_0 ));
    Odrv4 I__9552 (
            .O(N__41006),
            .I(\c0.data_in_frame_0_0 ));
    Odrv4 I__9551 (
            .O(N__41003),
            .I(\c0.data_in_frame_0_0 ));
    Odrv4 I__9550 (
            .O(N__41000),
            .I(\c0.data_in_frame_0_0 ));
    CascadeMux I__9549 (
            .O(N__40989),
            .I(N__40985));
    InMux I__9548 (
            .O(N__40988),
            .I(N__40979));
    InMux I__9547 (
            .O(N__40985),
            .I(N__40979));
    CascadeMux I__9546 (
            .O(N__40984),
            .I(N__40975));
    LocalMux I__9545 (
            .O(N__40979),
            .I(N__40972));
    InMux I__9544 (
            .O(N__40978),
            .I(N__40969));
    InMux I__9543 (
            .O(N__40975),
            .I(N__40966));
    Span4Mux_h I__9542 (
            .O(N__40972),
            .I(N__40963));
    LocalMux I__9541 (
            .O(N__40969),
            .I(N__40960));
    LocalMux I__9540 (
            .O(N__40966),
            .I(\c0.data_in_frame_1_7 ));
    Odrv4 I__9539 (
            .O(N__40963),
            .I(\c0.data_in_frame_1_7 ));
    Odrv4 I__9538 (
            .O(N__40960),
            .I(\c0.data_in_frame_1_7 ));
    InMux I__9537 (
            .O(N__40953),
            .I(N__40947));
    InMux I__9536 (
            .O(N__40952),
            .I(N__40947));
    LocalMux I__9535 (
            .O(N__40947),
            .I(N__40944));
    Span4Mux_h I__9534 (
            .O(N__40944),
            .I(N__40941));
    Odrv4 I__9533 (
            .O(N__40941),
            .I(\c0.n17213 ));
    CascadeMux I__9532 (
            .O(N__40938),
            .I(N__40935));
    InMux I__9531 (
            .O(N__40935),
            .I(N__40930));
    CascadeMux I__9530 (
            .O(N__40934),
            .I(N__40926));
    InMux I__9529 (
            .O(N__40933),
            .I(N__40922));
    LocalMux I__9528 (
            .O(N__40930),
            .I(N__40919));
    InMux I__9527 (
            .O(N__40929),
            .I(N__40914));
    InMux I__9526 (
            .O(N__40926),
            .I(N__40914));
    InMux I__9525 (
            .O(N__40925),
            .I(N__40911));
    LocalMux I__9524 (
            .O(N__40922),
            .I(N__40908));
    Span4Mux_v I__9523 (
            .O(N__40919),
            .I(N__40903));
    LocalMux I__9522 (
            .O(N__40914),
            .I(N__40903));
    LocalMux I__9521 (
            .O(N__40911),
            .I(data_out_frame2_8_5));
    Odrv12 I__9520 (
            .O(N__40908),
            .I(data_out_frame2_8_5));
    Odrv4 I__9519 (
            .O(N__40903),
            .I(data_out_frame2_8_5));
    InMux I__9518 (
            .O(N__40896),
            .I(N__40893));
    LocalMux I__9517 (
            .O(N__40893),
            .I(N__40888));
    InMux I__9516 (
            .O(N__40892),
            .I(N__40885));
    InMux I__9515 (
            .O(N__40891),
            .I(N__40882));
    Span4Mux_v I__9514 (
            .O(N__40888),
            .I(N__40879));
    LocalMux I__9513 (
            .O(N__40885),
            .I(N__40876));
    LocalMux I__9512 (
            .O(N__40882),
            .I(N__40873));
    Span4Mux_h I__9511 (
            .O(N__40879),
            .I(N__40868));
    Span4Mux_v I__9510 (
            .O(N__40876),
            .I(N__40868));
    Span4Mux_v I__9509 (
            .O(N__40873),
            .I(N__40865));
    Span4Mux_h I__9508 (
            .O(N__40868),
            .I(N__40858));
    Span4Mux_h I__9507 (
            .O(N__40865),
            .I(N__40858));
    InMux I__9506 (
            .O(N__40864),
            .I(N__40855));
    InMux I__9505 (
            .O(N__40863),
            .I(N__40852));
    Sp12to4 I__9504 (
            .O(N__40858),
            .I(N__40849));
    LocalMux I__9503 (
            .O(N__40855),
            .I(data_out_frame2_6_6));
    LocalMux I__9502 (
            .O(N__40852),
            .I(data_out_frame2_6_6));
    Odrv12 I__9501 (
            .O(N__40849),
            .I(data_out_frame2_6_6));
    CascadeMux I__9500 (
            .O(N__40842),
            .I(N__40839));
    InMux I__9499 (
            .O(N__40839),
            .I(N__40836));
    LocalMux I__9498 (
            .O(N__40836),
            .I(N__40833));
    Span4Mux_v I__9497 (
            .O(N__40833),
            .I(N__40830));
    Sp12to4 I__9496 (
            .O(N__40830),
            .I(N__40827));
    Span12Mux_s5_h I__9495 (
            .O(N__40827),
            .I(N__40824));
    Odrv12 I__9494 (
            .O(N__40824),
            .I(\c0.n10472 ));
    InMux I__9493 (
            .O(N__40821),
            .I(N__40815));
    InMux I__9492 (
            .O(N__40820),
            .I(N__40815));
    LocalMux I__9491 (
            .O(N__40815),
            .I(N__40811));
    InMux I__9490 (
            .O(N__40814),
            .I(N__40808));
    Span4Mux_v I__9489 (
            .O(N__40811),
            .I(N__40802));
    LocalMux I__9488 (
            .O(N__40808),
            .I(N__40802));
    InMux I__9487 (
            .O(N__40807),
            .I(N__40799));
    Span4Mux_h I__9486 (
            .O(N__40802),
            .I(N__40789));
    LocalMux I__9485 (
            .O(N__40799),
            .I(N__40786));
    InMux I__9484 (
            .O(N__40798),
            .I(N__40773));
    InMux I__9483 (
            .O(N__40797),
            .I(N__40773));
    InMux I__9482 (
            .O(N__40796),
            .I(N__40773));
    InMux I__9481 (
            .O(N__40795),
            .I(N__40773));
    InMux I__9480 (
            .O(N__40794),
            .I(N__40773));
    InMux I__9479 (
            .O(N__40793),
            .I(N__40773));
    InMux I__9478 (
            .O(N__40792),
            .I(N__40770));
    Odrv4 I__9477 (
            .O(N__40789),
            .I(\c0.n15821 ));
    Odrv4 I__9476 (
            .O(N__40786),
            .I(\c0.n15821 ));
    LocalMux I__9475 (
            .O(N__40773),
            .I(\c0.n15821 ));
    LocalMux I__9474 (
            .O(N__40770),
            .I(\c0.n15821 ));
    CascadeMux I__9473 (
            .O(N__40761),
            .I(N__40756));
    CascadeMux I__9472 (
            .O(N__40760),
            .I(N__40753));
    InMux I__9471 (
            .O(N__40759),
            .I(N__40750));
    InMux I__9470 (
            .O(N__40756),
            .I(N__40747));
    InMux I__9469 (
            .O(N__40753),
            .I(N__40744));
    LocalMux I__9468 (
            .O(N__40750),
            .I(N__40741));
    LocalMux I__9467 (
            .O(N__40747),
            .I(N__40738));
    LocalMux I__9466 (
            .O(N__40744),
            .I(\c0.FRAME_MATCHER_state_18 ));
    Odrv4 I__9465 (
            .O(N__40741),
            .I(\c0.FRAME_MATCHER_state_18 ));
    Odrv4 I__9464 (
            .O(N__40738),
            .I(\c0.FRAME_MATCHER_state_18 ));
    SRMux I__9463 (
            .O(N__40731),
            .I(N__40728));
    LocalMux I__9462 (
            .O(N__40728),
            .I(N__40725));
    Span4Mux_h I__9461 (
            .O(N__40725),
            .I(N__40722));
    Odrv4 I__9460 (
            .O(N__40722),
            .I(\c0.n8_adj_2329 ));
    InMux I__9459 (
            .O(N__40719),
            .I(N__40715));
    InMux I__9458 (
            .O(N__40718),
            .I(N__40712));
    LocalMux I__9457 (
            .O(N__40715),
            .I(N__40706));
    LocalMux I__9456 (
            .O(N__40712),
            .I(N__40706));
    CascadeMux I__9455 (
            .O(N__40711),
            .I(N__40703));
    Span4Mux_h I__9454 (
            .O(N__40706),
            .I(N__40699));
    InMux I__9453 (
            .O(N__40703),
            .I(N__40694));
    InMux I__9452 (
            .O(N__40702),
            .I(N__40694));
    Odrv4 I__9451 (
            .O(N__40699),
            .I(\c0.n8_adj_2385 ));
    LocalMux I__9450 (
            .O(N__40694),
            .I(\c0.n8_adj_2385 ));
    InMux I__9449 (
            .O(N__40689),
            .I(N__40686));
    LocalMux I__9448 (
            .O(N__40686),
            .I(N__40683));
    Odrv12 I__9447 (
            .O(N__40683),
            .I(\c0.n46 ));
    CascadeMux I__9446 (
            .O(N__40680),
            .I(N__40677));
    InMux I__9445 (
            .O(N__40677),
            .I(N__40674));
    LocalMux I__9444 (
            .O(N__40674),
            .I(N__40669));
    InMux I__9443 (
            .O(N__40673),
            .I(N__40664));
    InMux I__9442 (
            .O(N__40672),
            .I(N__40664));
    Span4Mux_h I__9441 (
            .O(N__40669),
            .I(N__40660));
    LocalMux I__9440 (
            .O(N__40664),
            .I(N__40657));
    CascadeMux I__9439 (
            .O(N__40663),
            .I(N__40654));
    Sp12to4 I__9438 (
            .O(N__40660),
            .I(N__40651));
    Span4Mux_h I__9437 (
            .O(N__40657),
            .I(N__40648));
    InMux I__9436 (
            .O(N__40654),
            .I(N__40645));
    Span12Mux_v I__9435 (
            .O(N__40651),
            .I(N__40642));
    Span4Mux_h I__9434 (
            .O(N__40648),
            .I(N__40639));
    LocalMux I__9433 (
            .O(N__40645),
            .I(\c0.data_out_frame2_0_0 ));
    Odrv12 I__9432 (
            .O(N__40642),
            .I(\c0.data_out_frame2_0_0 ));
    Odrv4 I__9431 (
            .O(N__40639),
            .I(\c0.data_out_frame2_0_0 ));
    InMux I__9430 (
            .O(N__40632),
            .I(N__40629));
    LocalMux I__9429 (
            .O(N__40629),
            .I(\c0.n17490 ));
    CascadeMux I__9428 (
            .O(N__40626),
            .I(N__40620));
    CascadeMux I__9427 (
            .O(N__40625),
            .I(N__40615));
    CascadeMux I__9426 (
            .O(N__40624),
            .I(N__40611));
    CascadeMux I__9425 (
            .O(N__40623),
            .I(N__40607));
    InMux I__9424 (
            .O(N__40620),
            .I(N__40601));
    InMux I__9423 (
            .O(N__40619),
            .I(N__40601));
    InMux I__9422 (
            .O(N__40618),
            .I(N__40595));
    InMux I__9421 (
            .O(N__40615),
            .I(N__40592));
    InMux I__9420 (
            .O(N__40614),
            .I(N__40587));
    InMux I__9419 (
            .O(N__40611),
            .I(N__40587));
    InMux I__9418 (
            .O(N__40610),
            .I(N__40584));
    InMux I__9417 (
            .O(N__40607),
            .I(N__40579));
    InMux I__9416 (
            .O(N__40606),
            .I(N__40579));
    LocalMux I__9415 (
            .O(N__40601),
            .I(N__40574));
    InMux I__9414 (
            .O(N__40600),
            .I(N__40571));
    InMux I__9413 (
            .O(N__40599),
            .I(N__40568));
    InMux I__9412 (
            .O(N__40598),
            .I(N__40564));
    LocalMux I__9411 (
            .O(N__40595),
            .I(N__40561));
    LocalMux I__9410 (
            .O(N__40592),
            .I(N__40558));
    LocalMux I__9409 (
            .O(N__40587),
            .I(N__40553));
    LocalMux I__9408 (
            .O(N__40584),
            .I(N__40553));
    LocalMux I__9407 (
            .O(N__40579),
            .I(N__40550));
    InMux I__9406 (
            .O(N__40578),
            .I(N__40545));
    InMux I__9405 (
            .O(N__40577),
            .I(N__40545));
    Span4Mux_v I__9404 (
            .O(N__40574),
            .I(N__40538));
    LocalMux I__9403 (
            .O(N__40571),
            .I(N__40538));
    LocalMux I__9402 (
            .O(N__40568),
            .I(N__40538));
    InMux I__9401 (
            .O(N__40567),
            .I(N__40535));
    LocalMux I__9400 (
            .O(N__40564),
            .I(N__40528));
    Span4Mux_v I__9399 (
            .O(N__40561),
            .I(N__40528));
    Span4Mux_v I__9398 (
            .O(N__40558),
            .I(N__40528));
    Span4Mux_h I__9397 (
            .O(N__40553),
            .I(N__40525));
    Span4Mux_v I__9396 (
            .O(N__40550),
            .I(N__40518));
    LocalMux I__9395 (
            .O(N__40545),
            .I(N__40518));
    Span4Mux_v I__9394 (
            .O(N__40538),
            .I(N__40518));
    LocalMux I__9393 (
            .O(N__40535),
            .I(\c0.n15171 ));
    Odrv4 I__9392 (
            .O(N__40528),
            .I(\c0.n15171 ));
    Odrv4 I__9391 (
            .O(N__40525),
            .I(\c0.n15171 ));
    Odrv4 I__9390 (
            .O(N__40518),
            .I(\c0.n15171 ));
    CascadeMux I__9389 (
            .O(N__40509),
            .I(N__40506));
    InMux I__9388 (
            .O(N__40506),
            .I(N__40496));
    InMux I__9387 (
            .O(N__40505),
            .I(N__40493));
    InMux I__9386 (
            .O(N__40504),
            .I(N__40490));
    InMux I__9385 (
            .O(N__40503),
            .I(N__40487));
    CascadeMux I__9384 (
            .O(N__40502),
            .I(N__40484));
    CascadeMux I__9383 (
            .O(N__40501),
            .I(N__40481));
    InMux I__9382 (
            .O(N__40500),
            .I(N__40478));
    InMux I__9381 (
            .O(N__40499),
            .I(N__40475));
    LocalMux I__9380 (
            .O(N__40496),
            .I(N__40472));
    LocalMux I__9379 (
            .O(N__40493),
            .I(N__40467));
    LocalMux I__9378 (
            .O(N__40490),
            .I(N__40467));
    LocalMux I__9377 (
            .O(N__40487),
            .I(N__40464));
    InMux I__9376 (
            .O(N__40484),
            .I(N__40461));
    InMux I__9375 (
            .O(N__40481),
            .I(N__40458));
    LocalMux I__9374 (
            .O(N__40478),
            .I(N__40455));
    LocalMux I__9373 (
            .O(N__40475),
            .I(N__40450));
    Span4Mux_h I__9372 (
            .O(N__40472),
            .I(N__40450));
    Span4Mux_v I__9371 (
            .O(N__40467),
            .I(N__40445));
    Span4Mux_v I__9370 (
            .O(N__40464),
            .I(N__40445));
    LocalMux I__9369 (
            .O(N__40461),
            .I(rx_data_7));
    LocalMux I__9368 (
            .O(N__40458),
            .I(rx_data_7));
    Odrv12 I__9367 (
            .O(N__40455),
            .I(rx_data_7));
    Odrv4 I__9366 (
            .O(N__40450),
            .I(rx_data_7));
    Odrv4 I__9365 (
            .O(N__40445),
            .I(rx_data_7));
    CascadeMux I__9364 (
            .O(N__40434),
            .I(N__40415));
    CascadeMux I__9363 (
            .O(N__40433),
            .I(N__40412));
    InMux I__9362 (
            .O(N__40432),
            .I(N__40403));
    InMux I__9361 (
            .O(N__40431),
            .I(N__40400));
    InMux I__9360 (
            .O(N__40430),
            .I(N__40397));
    InMux I__9359 (
            .O(N__40429),
            .I(N__40390));
    InMux I__9358 (
            .O(N__40428),
            .I(N__40390));
    InMux I__9357 (
            .O(N__40427),
            .I(N__40390));
    InMux I__9356 (
            .O(N__40426),
            .I(N__40387));
    InMux I__9355 (
            .O(N__40425),
            .I(N__40382));
    InMux I__9354 (
            .O(N__40424),
            .I(N__40382));
    InMux I__9353 (
            .O(N__40423),
            .I(N__40379));
    InMux I__9352 (
            .O(N__40422),
            .I(N__40374));
    InMux I__9351 (
            .O(N__40421),
            .I(N__40374));
    InMux I__9350 (
            .O(N__40420),
            .I(N__40367));
    InMux I__9349 (
            .O(N__40419),
            .I(N__40367));
    InMux I__9348 (
            .O(N__40418),
            .I(N__40367));
    InMux I__9347 (
            .O(N__40415),
            .I(N__40358));
    InMux I__9346 (
            .O(N__40412),
            .I(N__40358));
    InMux I__9345 (
            .O(N__40411),
            .I(N__40358));
    InMux I__9344 (
            .O(N__40410),
            .I(N__40358));
    InMux I__9343 (
            .O(N__40409),
            .I(N__40349));
    InMux I__9342 (
            .O(N__40408),
            .I(N__40349));
    InMux I__9341 (
            .O(N__40407),
            .I(N__40349));
    InMux I__9340 (
            .O(N__40406),
            .I(N__40349));
    LocalMux I__9339 (
            .O(N__40403),
            .I(N__40346));
    LocalMux I__9338 (
            .O(N__40400),
            .I(N__40341));
    LocalMux I__9337 (
            .O(N__40397),
            .I(N__40341));
    LocalMux I__9336 (
            .O(N__40390),
            .I(N__40338));
    LocalMux I__9335 (
            .O(N__40387),
            .I(\c0.n17076 ));
    LocalMux I__9334 (
            .O(N__40382),
            .I(\c0.n17076 ));
    LocalMux I__9333 (
            .O(N__40379),
            .I(\c0.n17076 ));
    LocalMux I__9332 (
            .O(N__40374),
            .I(\c0.n17076 ));
    LocalMux I__9331 (
            .O(N__40367),
            .I(\c0.n17076 ));
    LocalMux I__9330 (
            .O(N__40358),
            .I(\c0.n17076 ));
    LocalMux I__9329 (
            .O(N__40349),
            .I(\c0.n17076 ));
    Odrv4 I__9328 (
            .O(N__40346),
            .I(\c0.n17076 ));
    Odrv4 I__9327 (
            .O(N__40341),
            .I(\c0.n17076 ));
    Odrv4 I__9326 (
            .O(N__40338),
            .I(\c0.n17076 ));
    InMux I__9325 (
            .O(N__40317),
            .I(N__40310));
    InMux I__9324 (
            .O(N__40316),
            .I(N__40305));
    InMux I__9323 (
            .O(N__40315),
            .I(N__40305));
    InMux I__9322 (
            .O(N__40314),
            .I(N__40300));
    InMux I__9321 (
            .O(N__40313),
            .I(N__40300));
    LocalMux I__9320 (
            .O(N__40310),
            .I(\c0.n26_adj_2174 ));
    LocalMux I__9319 (
            .O(N__40305),
            .I(\c0.n26_adj_2174 ));
    LocalMux I__9318 (
            .O(N__40300),
            .I(\c0.n26_adj_2174 ));
    CascadeMux I__9317 (
            .O(N__40293),
            .I(\c0.n17487_cascade_ ));
    InMux I__9316 (
            .O(N__40290),
            .I(N__40287));
    LocalMux I__9315 (
            .O(N__40287),
            .I(N__40283));
    InMux I__9314 (
            .O(N__40286),
            .I(N__40280));
    Span4Mux_v I__9313 (
            .O(N__40283),
            .I(N__40277));
    LocalMux I__9312 (
            .O(N__40280),
            .I(N__40274));
    Span4Mux_h I__9311 (
            .O(N__40277),
            .I(N__40267));
    Span4Mux_h I__9310 (
            .O(N__40274),
            .I(N__40267));
    InMux I__9309 (
            .O(N__40273),
            .I(N__40264));
    InMux I__9308 (
            .O(N__40272),
            .I(N__40261));
    Span4Mux_h I__9307 (
            .O(N__40267),
            .I(N__40258));
    LocalMux I__9306 (
            .O(N__40264),
            .I(N__40255));
    LocalMux I__9305 (
            .O(N__40261),
            .I(\c0.data_out_frame2_0_1 ));
    Odrv4 I__9304 (
            .O(N__40258),
            .I(\c0.data_out_frame2_0_1 ));
    Odrv12 I__9303 (
            .O(N__40255),
            .I(\c0.data_out_frame2_0_1 ));
    InMux I__9302 (
            .O(N__40248),
            .I(N__40240));
    InMux I__9301 (
            .O(N__40247),
            .I(N__40236));
    InMux I__9300 (
            .O(N__40246),
            .I(N__40227));
    InMux I__9299 (
            .O(N__40245),
            .I(N__40227));
    InMux I__9298 (
            .O(N__40244),
            .I(N__40227));
    InMux I__9297 (
            .O(N__40243),
            .I(N__40224));
    LocalMux I__9296 (
            .O(N__40240),
            .I(N__40221));
    InMux I__9295 (
            .O(N__40239),
            .I(N__40216));
    LocalMux I__9294 (
            .O(N__40236),
            .I(N__40213));
    InMux I__9293 (
            .O(N__40235),
            .I(N__40208));
    InMux I__9292 (
            .O(N__40234),
            .I(N__40208));
    LocalMux I__9291 (
            .O(N__40227),
            .I(N__40203));
    LocalMux I__9290 (
            .O(N__40224),
            .I(N__40203));
    Span4Mux_h I__9289 (
            .O(N__40221),
            .I(N__40200));
    CascadeMux I__9288 (
            .O(N__40220),
            .I(N__40194));
    InMux I__9287 (
            .O(N__40219),
            .I(N__40189));
    LocalMux I__9286 (
            .O(N__40216),
            .I(N__40186));
    Span4Mux_h I__9285 (
            .O(N__40213),
            .I(N__40181));
    LocalMux I__9284 (
            .O(N__40208),
            .I(N__40181));
    Span4Mux_v I__9283 (
            .O(N__40203),
            .I(N__40176));
    Span4Mux_h I__9282 (
            .O(N__40200),
            .I(N__40176));
    InMux I__9281 (
            .O(N__40199),
            .I(N__40171));
    InMux I__9280 (
            .O(N__40198),
            .I(N__40171));
    InMux I__9279 (
            .O(N__40197),
            .I(N__40168));
    InMux I__9278 (
            .O(N__40194),
            .I(N__40161));
    InMux I__9277 (
            .O(N__40193),
            .I(N__40161));
    InMux I__9276 (
            .O(N__40192),
            .I(N__40161));
    LocalMux I__9275 (
            .O(N__40189),
            .I(FRAME_MATCHER_state_0));
    Odrv4 I__9274 (
            .O(N__40186),
            .I(FRAME_MATCHER_state_0));
    Odrv4 I__9273 (
            .O(N__40181),
            .I(FRAME_MATCHER_state_0));
    Odrv4 I__9272 (
            .O(N__40176),
            .I(FRAME_MATCHER_state_0));
    LocalMux I__9271 (
            .O(N__40171),
            .I(FRAME_MATCHER_state_0));
    LocalMux I__9270 (
            .O(N__40168),
            .I(FRAME_MATCHER_state_0));
    LocalMux I__9269 (
            .O(N__40161),
            .I(FRAME_MATCHER_state_0));
    CascadeMux I__9268 (
            .O(N__40146),
            .I(N__40137));
    InMux I__9267 (
            .O(N__40145),
            .I(N__40134));
    InMux I__9266 (
            .O(N__40144),
            .I(N__40129));
    InMux I__9265 (
            .O(N__40143),
            .I(N__40129));
    InMux I__9264 (
            .O(N__40142),
            .I(N__40126));
    InMux I__9263 (
            .O(N__40141),
            .I(N__40121));
    InMux I__9262 (
            .O(N__40140),
            .I(N__40121));
    InMux I__9261 (
            .O(N__40137),
            .I(N__40118));
    LocalMux I__9260 (
            .O(N__40134),
            .I(\c0.n12491 ));
    LocalMux I__9259 (
            .O(N__40129),
            .I(\c0.n12491 ));
    LocalMux I__9258 (
            .O(N__40126),
            .I(\c0.n12491 ));
    LocalMux I__9257 (
            .O(N__40121),
            .I(\c0.n12491 ));
    LocalMux I__9256 (
            .O(N__40118),
            .I(\c0.n12491 ));
    CascadeMux I__9255 (
            .O(N__40107),
            .I(\c0.n17690_cascade_ ));
    InMux I__9254 (
            .O(N__40104),
            .I(N__40100));
    InMux I__9253 (
            .O(N__40103),
            .I(N__40097));
    LocalMux I__9252 (
            .O(N__40100),
            .I(N__40094));
    LocalMux I__9251 (
            .O(N__40097),
            .I(N__40090));
    Span4Mux_v I__9250 (
            .O(N__40094),
            .I(N__40086));
    InMux I__9249 (
            .O(N__40093),
            .I(N__40083));
    Span4Mux_h I__9248 (
            .O(N__40090),
            .I(N__40080));
    CascadeMux I__9247 (
            .O(N__40089),
            .I(N__40076));
    Sp12to4 I__9246 (
            .O(N__40086),
            .I(N__40071));
    LocalMux I__9245 (
            .O(N__40083),
            .I(N__40071));
    Span4Mux_h I__9244 (
            .O(N__40080),
            .I(N__40068));
    InMux I__9243 (
            .O(N__40079),
            .I(N__40063));
    InMux I__9242 (
            .O(N__40076),
            .I(N__40063));
    Span12Mux_s5_h I__9241 (
            .O(N__40071),
            .I(N__40060));
    Span4Mux_h I__9240 (
            .O(N__40068),
            .I(N__40057));
    LocalMux I__9239 (
            .O(N__40063),
            .I(\c0.data_out_frame2_0_2 ));
    Odrv12 I__9238 (
            .O(N__40060),
            .I(\c0.data_out_frame2_0_2 ));
    Odrv4 I__9237 (
            .O(N__40057),
            .I(\c0.data_out_frame2_0_2 ));
    InMux I__9236 (
            .O(N__40050),
            .I(N__40046));
    InMux I__9235 (
            .O(N__40049),
            .I(N__40043));
    LocalMux I__9234 (
            .O(N__40046),
            .I(N__40040));
    LocalMux I__9233 (
            .O(N__40043),
            .I(N__40037));
    Span4Mux_h I__9232 (
            .O(N__40040),
            .I(N__40034));
    Span4Mux_h I__9231 (
            .O(N__40037),
            .I(N__40031));
    Odrv4 I__9230 (
            .O(N__40034),
            .I(\c0.data_in_frame_5_2 ));
    Odrv4 I__9229 (
            .O(N__40031),
            .I(\c0.data_in_frame_5_2 ));
    InMux I__9228 (
            .O(N__40026),
            .I(N__40023));
    LocalMux I__9227 (
            .O(N__40023),
            .I(N__40016));
    InMux I__9226 (
            .O(N__40022),
            .I(N__40011));
    InMux I__9225 (
            .O(N__40021),
            .I(N__40011));
    InMux I__9224 (
            .O(N__40020),
            .I(N__40006));
    InMux I__9223 (
            .O(N__40019),
            .I(N__40006));
    Odrv12 I__9222 (
            .O(N__40016),
            .I(\c0.data_in_frame_1_0 ));
    LocalMux I__9221 (
            .O(N__40011),
            .I(\c0.data_in_frame_1_0 ));
    LocalMux I__9220 (
            .O(N__40006),
            .I(\c0.data_in_frame_1_0 ));
    InMux I__9219 (
            .O(N__39999),
            .I(N__39995));
    CascadeMux I__9218 (
            .O(N__39998),
            .I(N__39990));
    LocalMux I__9217 (
            .O(N__39995),
            .I(N__39987));
    InMux I__9216 (
            .O(N__39994),
            .I(N__39984));
    InMux I__9215 (
            .O(N__39993),
            .I(N__39980));
    InMux I__9214 (
            .O(N__39990),
            .I(N__39977));
    Span4Mux_h I__9213 (
            .O(N__39987),
            .I(N__39972));
    LocalMux I__9212 (
            .O(N__39984),
            .I(N__39972));
    InMux I__9211 (
            .O(N__39983),
            .I(N__39969));
    LocalMux I__9210 (
            .O(N__39980),
            .I(N__39966));
    LocalMux I__9209 (
            .O(N__39977),
            .I(\c0.data_in_frame_1_1 ));
    Odrv4 I__9208 (
            .O(N__39972),
            .I(\c0.data_in_frame_1_1 ));
    LocalMux I__9207 (
            .O(N__39969),
            .I(\c0.data_in_frame_1_1 ));
    Odrv4 I__9206 (
            .O(N__39966),
            .I(\c0.data_in_frame_1_1 ));
    InMux I__9205 (
            .O(N__39957),
            .I(N__39954));
    LocalMux I__9204 (
            .O(N__39954),
            .I(\c0.n17102 ));
    InMux I__9203 (
            .O(N__39951),
            .I(N__39948));
    LocalMux I__9202 (
            .O(N__39948),
            .I(N__39940));
    InMux I__9201 (
            .O(N__39947),
            .I(N__39937));
    InMux I__9200 (
            .O(N__39946),
            .I(N__39929));
    InMux I__9199 (
            .O(N__39945),
            .I(N__39929));
    InMux I__9198 (
            .O(N__39944),
            .I(N__39924));
    InMux I__9197 (
            .O(N__39943),
            .I(N__39924));
    Span4Mux_v I__9196 (
            .O(N__39940),
            .I(N__39921));
    LocalMux I__9195 (
            .O(N__39937),
            .I(N__39918));
    InMux I__9194 (
            .O(N__39936),
            .I(N__39915));
    InMux I__9193 (
            .O(N__39935),
            .I(N__39910));
    InMux I__9192 (
            .O(N__39934),
            .I(N__39910));
    LocalMux I__9191 (
            .O(N__39929),
            .I(N__39905));
    LocalMux I__9190 (
            .O(N__39924),
            .I(N__39905));
    Sp12to4 I__9189 (
            .O(N__39921),
            .I(N__39902));
    Span4Mux_h I__9188 (
            .O(N__39918),
            .I(N__39899));
    LocalMux I__9187 (
            .O(N__39915),
            .I(N__39896));
    LocalMux I__9186 (
            .O(N__39910),
            .I(N__39893));
    Span4Mux_h I__9185 (
            .O(N__39905),
            .I(N__39890));
    Odrv12 I__9184 (
            .O(N__39902),
            .I(\c0.n5815 ));
    Odrv4 I__9183 (
            .O(N__39899),
            .I(\c0.n5815 ));
    Odrv4 I__9182 (
            .O(N__39896),
            .I(\c0.n5815 ));
    Odrv4 I__9181 (
            .O(N__39893),
            .I(\c0.n5815 ));
    Odrv4 I__9180 (
            .O(N__39890),
            .I(\c0.n5815 ));
    InMux I__9179 (
            .O(N__39879),
            .I(N__39871));
    InMux I__9178 (
            .O(N__39878),
            .I(N__39866));
    InMux I__9177 (
            .O(N__39877),
            .I(N__39866));
    InMux I__9176 (
            .O(N__39876),
            .I(N__39863));
    InMux I__9175 (
            .O(N__39875),
            .I(N__39860));
    InMux I__9174 (
            .O(N__39874),
            .I(N__39857));
    LocalMux I__9173 (
            .O(N__39871),
            .I(\c0.n4494 ));
    LocalMux I__9172 (
            .O(N__39866),
            .I(\c0.n4494 ));
    LocalMux I__9171 (
            .O(N__39863),
            .I(\c0.n4494 ));
    LocalMux I__9170 (
            .O(N__39860),
            .I(\c0.n4494 ));
    LocalMux I__9169 (
            .O(N__39857),
            .I(\c0.n4494 ));
    CascadeMux I__9168 (
            .O(N__39846),
            .I(N__39841));
    CascadeMux I__9167 (
            .O(N__39845),
            .I(N__39838));
    CascadeMux I__9166 (
            .O(N__39844),
            .I(N__39832));
    InMux I__9165 (
            .O(N__39841),
            .I(N__39828));
    InMux I__9164 (
            .O(N__39838),
            .I(N__39821));
    InMux I__9163 (
            .O(N__39837),
            .I(N__39818));
    InMux I__9162 (
            .O(N__39836),
            .I(N__39815));
    InMux I__9161 (
            .O(N__39835),
            .I(N__39812));
    InMux I__9160 (
            .O(N__39832),
            .I(N__39807));
    InMux I__9159 (
            .O(N__39831),
            .I(N__39807));
    LocalMux I__9158 (
            .O(N__39828),
            .I(N__39804));
    InMux I__9157 (
            .O(N__39827),
            .I(N__39795));
    InMux I__9156 (
            .O(N__39826),
            .I(N__39795));
    InMux I__9155 (
            .O(N__39825),
            .I(N__39795));
    InMux I__9154 (
            .O(N__39824),
            .I(N__39795));
    LocalMux I__9153 (
            .O(N__39821),
            .I(N__39792));
    LocalMux I__9152 (
            .O(N__39818),
            .I(N__39789));
    LocalMux I__9151 (
            .O(N__39815),
            .I(N__39782));
    LocalMux I__9150 (
            .O(N__39812),
            .I(N__39782));
    LocalMux I__9149 (
            .O(N__39807),
            .I(N__39782));
    Span4Mux_h I__9148 (
            .O(N__39804),
            .I(N__39779));
    LocalMux I__9147 (
            .O(N__39795),
            .I(N__39776));
    Span4Mux_h I__9146 (
            .O(N__39792),
            .I(N__39773));
    Span4Mux_v I__9145 (
            .O(N__39789),
            .I(N__39768));
    Span4Mux_v I__9144 (
            .O(N__39782),
            .I(N__39768));
    Odrv4 I__9143 (
            .O(N__39779),
            .I(\c0.n5817 ));
    Odrv4 I__9142 (
            .O(N__39776),
            .I(\c0.n5817 ));
    Odrv4 I__9141 (
            .O(N__39773),
            .I(\c0.n5817 ));
    Odrv4 I__9140 (
            .O(N__39768),
            .I(\c0.n5817 ));
    InMux I__9139 (
            .O(N__39759),
            .I(N__39755));
    InMux I__9138 (
            .O(N__39758),
            .I(N__39750));
    LocalMux I__9137 (
            .O(N__39755),
            .I(N__39747));
    InMux I__9136 (
            .O(N__39754),
            .I(N__39742));
    InMux I__9135 (
            .O(N__39753),
            .I(N__39742));
    LocalMux I__9134 (
            .O(N__39750),
            .I(N__39739));
    Span12Mux_h I__9133 (
            .O(N__39747),
            .I(N__39734));
    LocalMux I__9132 (
            .O(N__39742),
            .I(N__39734));
    Odrv12 I__9131 (
            .O(N__39739),
            .I(n31_adj_2415));
    Odrv12 I__9130 (
            .O(N__39734),
            .I(n31_adj_2415));
    CascadeMux I__9129 (
            .O(N__39729),
            .I(N__39726));
    InMux I__9128 (
            .O(N__39726),
            .I(N__39719));
    InMux I__9127 (
            .O(N__39725),
            .I(N__39719));
    InMux I__9126 (
            .O(N__39724),
            .I(N__39716));
    LocalMux I__9125 (
            .O(N__39719),
            .I(\c0.n18202 ));
    LocalMux I__9124 (
            .O(N__39716),
            .I(\c0.n18202 ));
    InMux I__9123 (
            .O(N__39711),
            .I(N__39708));
    LocalMux I__9122 (
            .O(N__39708),
            .I(N__39705));
    Odrv12 I__9121 (
            .O(N__39705),
            .I(\c0.n17712 ));
    InMux I__9120 (
            .O(N__39702),
            .I(N__39698));
    CascadeMux I__9119 (
            .O(N__39701),
            .I(N__39694));
    LocalMux I__9118 (
            .O(N__39698),
            .I(N__39690));
    CascadeMux I__9117 (
            .O(N__39697),
            .I(N__39687));
    InMux I__9116 (
            .O(N__39694),
            .I(N__39684));
    CascadeMux I__9115 (
            .O(N__39693),
            .I(N__39680));
    Sp12to4 I__9114 (
            .O(N__39690),
            .I(N__39675));
    InMux I__9113 (
            .O(N__39687),
            .I(N__39672));
    LocalMux I__9112 (
            .O(N__39684),
            .I(N__39669));
    CascadeMux I__9111 (
            .O(N__39683),
            .I(N__39666));
    InMux I__9110 (
            .O(N__39680),
            .I(N__39663));
    CascadeMux I__9109 (
            .O(N__39679),
            .I(N__39660));
    CascadeMux I__9108 (
            .O(N__39678),
            .I(N__39657));
    Span12Mux_v I__9107 (
            .O(N__39675),
            .I(N__39652));
    LocalMux I__9106 (
            .O(N__39672),
            .I(N__39652));
    Span4Mux_v I__9105 (
            .O(N__39669),
            .I(N__39649));
    InMux I__9104 (
            .O(N__39666),
            .I(N__39646));
    LocalMux I__9103 (
            .O(N__39663),
            .I(N__39643));
    InMux I__9102 (
            .O(N__39660),
            .I(N__39640));
    InMux I__9101 (
            .O(N__39657),
            .I(N__39637));
    Odrv12 I__9100 (
            .O(N__39652),
            .I(\c0.n11867 ));
    Odrv4 I__9099 (
            .O(N__39649),
            .I(\c0.n11867 ));
    LocalMux I__9098 (
            .O(N__39646),
            .I(\c0.n11867 ));
    Odrv4 I__9097 (
            .O(N__39643),
            .I(\c0.n11867 ));
    LocalMux I__9096 (
            .O(N__39640),
            .I(\c0.n11867 ));
    LocalMux I__9095 (
            .O(N__39637),
            .I(\c0.n11867 ));
    InMux I__9094 (
            .O(N__39624),
            .I(N__39619));
    InMux I__9093 (
            .O(N__39623),
            .I(N__39616));
    CascadeMux I__9092 (
            .O(N__39622),
            .I(N__39613));
    LocalMux I__9091 (
            .O(N__39619),
            .I(N__39609));
    LocalMux I__9090 (
            .O(N__39616),
            .I(N__39606));
    InMux I__9089 (
            .O(N__39613),
            .I(N__39603));
    InMux I__9088 (
            .O(N__39612),
            .I(N__39600));
    Span4Mux_v I__9087 (
            .O(N__39609),
            .I(N__39593));
    Span4Mux_h I__9086 (
            .O(N__39606),
            .I(N__39593));
    LocalMux I__9085 (
            .O(N__39603),
            .I(N__39593));
    LocalMux I__9084 (
            .O(N__39600),
            .I(\c0.byte_transmit_counter2_5 ));
    Odrv4 I__9083 (
            .O(N__39593),
            .I(\c0.byte_transmit_counter2_5 ));
    SRMux I__9082 (
            .O(N__39588),
            .I(N__39585));
    LocalMux I__9081 (
            .O(N__39585),
            .I(N__39582));
    Span4Mux_h I__9080 (
            .O(N__39582),
            .I(N__39579));
    Odrv4 I__9079 (
            .O(N__39579),
            .I(\c0.n4_adj_2147 ));
    InMux I__9078 (
            .O(N__39576),
            .I(N__39573));
    LocalMux I__9077 (
            .O(N__39573),
            .I(N__39569));
    InMux I__9076 (
            .O(N__39572),
            .I(N__39566));
    Span4Mux_v I__9075 (
            .O(N__39569),
            .I(N__39563));
    LocalMux I__9074 (
            .O(N__39566),
            .I(N__39560));
    Odrv4 I__9073 (
            .O(N__39563),
            .I(n13116));
    Odrv12 I__9072 (
            .O(N__39560),
            .I(n13116));
    CascadeMux I__9071 (
            .O(N__39555),
            .I(N__39549));
    CascadeMux I__9070 (
            .O(N__39554),
            .I(N__39546));
    InMux I__9069 (
            .O(N__39553),
            .I(N__39542));
    InMux I__9068 (
            .O(N__39552),
            .I(N__39538));
    InMux I__9067 (
            .O(N__39549),
            .I(N__39535));
    InMux I__9066 (
            .O(N__39546),
            .I(N__39530));
    InMux I__9065 (
            .O(N__39545),
            .I(N__39530));
    LocalMux I__9064 (
            .O(N__39542),
            .I(N__39527));
    InMux I__9063 (
            .O(N__39541),
            .I(N__39524));
    LocalMux I__9062 (
            .O(N__39538),
            .I(N__39520));
    LocalMux I__9061 (
            .O(N__39535),
            .I(N__39516));
    LocalMux I__9060 (
            .O(N__39530),
            .I(N__39511));
    Span4Mux_v I__9059 (
            .O(N__39527),
            .I(N__39511));
    LocalMux I__9058 (
            .O(N__39524),
            .I(N__39508));
    CascadeMux I__9057 (
            .O(N__39523),
            .I(N__39505));
    Span4Mux_h I__9056 (
            .O(N__39520),
            .I(N__39502));
    InMux I__9055 (
            .O(N__39519),
            .I(N__39499));
    Span4Mux_v I__9054 (
            .O(N__39516),
            .I(N__39492));
    Span4Mux_h I__9053 (
            .O(N__39511),
            .I(N__39492));
    Span4Mux_v I__9052 (
            .O(N__39508),
            .I(N__39492));
    InMux I__9051 (
            .O(N__39505),
            .I(N__39489));
    Odrv4 I__9050 (
            .O(N__39502),
            .I(rx_data_6));
    LocalMux I__9049 (
            .O(N__39499),
            .I(rx_data_6));
    Odrv4 I__9048 (
            .O(N__39492),
            .I(rx_data_6));
    LocalMux I__9047 (
            .O(N__39489),
            .I(rx_data_6));
    CascadeMux I__9046 (
            .O(N__39480),
            .I(N__39473));
    InMux I__9045 (
            .O(N__39479),
            .I(N__39470));
    CascadeMux I__9044 (
            .O(N__39478),
            .I(N__39466));
    InMux I__9043 (
            .O(N__39477),
            .I(N__39463));
    InMux I__9042 (
            .O(N__39476),
            .I(N__39459));
    InMux I__9041 (
            .O(N__39473),
            .I(N__39456));
    LocalMux I__9040 (
            .O(N__39470),
            .I(N__39453));
    CascadeMux I__9039 (
            .O(N__39469),
            .I(N__39450));
    InMux I__9038 (
            .O(N__39466),
            .I(N__39447));
    LocalMux I__9037 (
            .O(N__39463),
            .I(N__39443));
    CascadeMux I__9036 (
            .O(N__39462),
            .I(N__39440));
    LocalMux I__9035 (
            .O(N__39459),
            .I(N__39433));
    LocalMux I__9034 (
            .O(N__39456),
            .I(N__39433));
    Span4Mux_h I__9033 (
            .O(N__39453),
            .I(N__39433));
    InMux I__9032 (
            .O(N__39450),
            .I(N__39430));
    LocalMux I__9031 (
            .O(N__39447),
            .I(N__39427));
    CascadeMux I__9030 (
            .O(N__39446),
            .I(N__39424));
    Span4Mux_h I__9029 (
            .O(N__39443),
            .I(N__39421));
    InMux I__9028 (
            .O(N__39440),
            .I(N__39418));
    Span4Mux_h I__9027 (
            .O(N__39433),
            .I(N__39415));
    LocalMux I__9026 (
            .O(N__39430),
            .I(N__39410));
    Span4Mux_v I__9025 (
            .O(N__39427),
            .I(N__39410));
    InMux I__9024 (
            .O(N__39424),
            .I(N__39407));
    Odrv4 I__9023 (
            .O(N__39421),
            .I(rx_data_1));
    LocalMux I__9022 (
            .O(N__39418),
            .I(rx_data_1));
    Odrv4 I__9021 (
            .O(N__39415),
            .I(rx_data_1));
    Odrv4 I__9020 (
            .O(N__39410),
            .I(rx_data_1));
    LocalMux I__9019 (
            .O(N__39407),
            .I(rx_data_1));
    CascadeMux I__9018 (
            .O(N__39396),
            .I(N__39391));
    InMux I__9017 (
            .O(N__39395),
            .I(N__39382));
    InMux I__9016 (
            .O(N__39394),
            .I(N__39379));
    InMux I__9015 (
            .O(N__39391),
            .I(N__39376));
    InMux I__9014 (
            .O(N__39390),
            .I(N__39373));
    InMux I__9013 (
            .O(N__39389),
            .I(N__39363));
    InMux I__9012 (
            .O(N__39388),
            .I(N__39363));
    InMux I__9011 (
            .O(N__39387),
            .I(N__39363));
    InMux I__9010 (
            .O(N__39386),
            .I(N__39354));
    InMux I__9009 (
            .O(N__39385),
            .I(N__39354));
    LocalMux I__9008 (
            .O(N__39382),
            .I(N__39351));
    LocalMux I__9007 (
            .O(N__39379),
            .I(N__39348));
    LocalMux I__9006 (
            .O(N__39376),
            .I(N__39343));
    LocalMux I__9005 (
            .O(N__39373),
            .I(N__39343));
    InMux I__9004 (
            .O(N__39372),
            .I(N__39336));
    InMux I__9003 (
            .O(N__39371),
            .I(N__39336));
    InMux I__9002 (
            .O(N__39370),
            .I(N__39336));
    LocalMux I__9001 (
            .O(N__39363),
            .I(N__39333));
    InMux I__9000 (
            .O(N__39362),
            .I(N__39330));
    InMux I__8999 (
            .O(N__39361),
            .I(N__39327));
    InMux I__8998 (
            .O(N__39360),
            .I(N__39324));
    InMux I__8997 (
            .O(N__39359),
            .I(N__39321));
    LocalMux I__8996 (
            .O(N__39354),
            .I(N__39318));
    Span4Mux_h I__8995 (
            .O(N__39351),
            .I(N__39311));
    Span4Mux_h I__8994 (
            .O(N__39348),
            .I(N__39311));
    Span4Mux_v I__8993 (
            .O(N__39343),
            .I(N__39311));
    LocalMux I__8992 (
            .O(N__39336),
            .I(N__39306));
    Span4Mux_v I__8991 (
            .O(N__39333),
            .I(N__39306));
    LocalMux I__8990 (
            .O(N__39330),
            .I(N__39303));
    LocalMux I__8989 (
            .O(N__39327),
            .I(\c0.n17072 ));
    LocalMux I__8988 (
            .O(N__39324),
            .I(\c0.n17072 ));
    LocalMux I__8987 (
            .O(N__39321),
            .I(\c0.n17072 ));
    Odrv4 I__8986 (
            .O(N__39318),
            .I(\c0.n17072 ));
    Odrv4 I__8985 (
            .O(N__39311),
            .I(\c0.n17072 ));
    Odrv4 I__8984 (
            .O(N__39306),
            .I(\c0.n17072 ));
    Odrv4 I__8983 (
            .O(N__39303),
            .I(\c0.n17072 ));
    CascadeMux I__8982 (
            .O(N__39288),
            .I(N__39285));
    InMux I__8981 (
            .O(N__39285),
            .I(N__39282));
    LocalMux I__8980 (
            .O(N__39282),
            .I(N__39278));
    InMux I__8979 (
            .O(N__39281),
            .I(N__39275));
    Span4Mux_h I__8978 (
            .O(N__39278),
            .I(N__39272));
    LocalMux I__8977 (
            .O(N__39275),
            .I(\c0.data_in_frame_3_1 ));
    Odrv4 I__8976 (
            .O(N__39272),
            .I(\c0.data_in_frame_3_1 ));
    CascadeMux I__8975 (
            .O(N__39267),
            .I(\c0.n17472_cascade_ ));
    InMux I__8974 (
            .O(N__39264),
            .I(N__39260));
    InMux I__8973 (
            .O(N__39263),
            .I(N__39255));
    LocalMux I__8972 (
            .O(N__39260),
            .I(N__39252));
    InMux I__8971 (
            .O(N__39259),
            .I(N__39249));
    CascadeMux I__8970 (
            .O(N__39258),
            .I(N__39246));
    LocalMux I__8969 (
            .O(N__39255),
            .I(N__39243));
    Span4Mux_v I__8968 (
            .O(N__39252),
            .I(N__39238));
    LocalMux I__8967 (
            .O(N__39249),
            .I(N__39238));
    InMux I__8966 (
            .O(N__39246),
            .I(N__39235));
    Span4Mux_v I__8965 (
            .O(N__39243),
            .I(N__39232));
    Span4Mux_h I__8964 (
            .O(N__39238),
            .I(N__39229));
    LocalMux I__8963 (
            .O(N__39235),
            .I(\c0.data_out_frame2_0_6 ));
    Odrv4 I__8962 (
            .O(N__39232),
            .I(\c0.data_out_frame2_0_6 ));
    Odrv4 I__8961 (
            .O(N__39229),
            .I(\c0.data_out_frame2_0_6 ));
    InMux I__8960 (
            .O(N__39222),
            .I(N__39201));
    InMux I__8959 (
            .O(N__39221),
            .I(N__39195));
    InMux I__8958 (
            .O(N__39220),
            .I(N__39195));
    CascadeMux I__8957 (
            .O(N__39219),
            .I(N__39191));
    CascadeMux I__8956 (
            .O(N__39218),
            .I(N__39187));
    InMux I__8955 (
            .O(N__39217),
            .I(N__39179));
    InMux I__8954 (
            .O(N__39216),
            .I(N__39179));
    InMux I__8953 (
            .O(N__39215),
            .I(N__39174));
    InMux I__8952 (
            .O(N__39214),
            .I(N__39174));
    InMux I__8951 (
            .O(N__39213),
            .I(N__39163));
    InMux I__8950 (
            .O(N__39212),
            .I(N__39163));
    InMux I__8949 (
            .O(N__39211),
            .I(N__39163));
    InMux I__8948 (
            .O(N__39210),
            .I(N__39163));
    InMux I__8947 (
            .O(N__39209),
            .I(N__39163));
    InMux I__8946 (
            .O(N__39208),
            .I(N__39160));
    InMux I__8945 (
            .O(N__39207),
            .I(N__39157));
    InMux I__8944 (
            .O(N__39206),
            .I(N__39154));
    InMux I__8943 (
            .O(N__39205),
            .I(N__39149));
    InMux I__8942 (
            .O(N__39204),
            .I(N__39149));
    LocalMux I__8941 (
            .O(N__39201),
            .I(N__39146));
    InMux I__8940 (
            .O(N__39200),
            .I(N__39143));
    LocalMux I__8939 (
            .O(N__39195),
            .I(N__39139));
    InMux I__8938 (
            .O(N__39194),
            .I(N__39136));
    InMux I__8937 (
            .O(N__39191),
            .I(N__39133));
    InMux I__8936 (
            .O(N__39190),
            .I(N__39126));
    InMux I__8935 (
            .O(N__39187),
            .I(N__39119));
    InMux I__8934 (
            .O(N__39186),
            .I(N__39119));
    InMux I__8933 (
            .O(N__39185),
            .I(N__39119));
    InMux I__8932 (
            .O(N__39184),
            .I(N__39116));
    LocalMux I__8931 (
            .O(N__39179),
            .I(N__39103));
    LocalMux I__8930 (
            .O(N__39174),
            .I(N__39103));
    LocalMux I__8929 (
            .O(N__39163),
            .I(N__39103));
    LocalMux I__8928 (
            .O(N__39160),
            .I(N__39103));
    LocalMux I__8927 (
            .O(N__39157),
            .I(N__39103));
    LocalMux I__8926 (
            .O(N__39154),
            .I(N__39103));
    LocalMux I__8925 (
            .O(N__39149),
            .I(N__39096));
    Span4Mux_v I__8924 (
            .O(N__39146),
            .I(N__39096));
    LocalMux I__8923 (
            .O(N__39143),
            .I(N__39096));
    InMux I__8922 (
            .O(N__39142),
            .I(N__39090));
    Span4Mux_v I__8921 (
            .O(N__39139),
            .I(N__39087));
    LocalMux I__8920 (
            .O(N__39136),
            .I(N__39082));
    LocalMux I__8919 (
            .O(N__39133),
            .I(N__39082));
    InMux I__8918 (
            .O(N__39132),
            .I(N__39079));
    InMux I__8917 (
            .O(N__39131),
            .I(N__39072));
    InMux I__8916 (
            .O(N__39130),
            .I(N__39072));
    InMux I__8915 (
            .O(N__39129),
            .I(N__39072));
    LocalMux I__8914 (
            .O(N__39126),
            .I(N__39067));
    LocalMux I__8913 (
            .O(N__39119),
            .I(N__39067));
    LocalMux I__8912 (
            .O(N__39116),
            .I(N__39060));
    Span4Mux_v I__8911 (
            .O(N__39103),
            .I(N__39060));
    Span4Mux_h I__8910 (
            .O(N__39096),
            .I(N__39060));
    InMux I__8909 (
            .O(N__39095),
            .I(N__39056));
    InMux I__8908 (
            .O(N__39094),
            .I(N__39051));
    InMux I__8907 (
            .O(N__39093),
            .I(N__39051));
    LocalMux I__8906 (
            .O(N__39090),
            .I(N__39044));
    Span4Mux_h I__8905 (
            .O(N__39087),
            .I(N__39044));
    Span4Mux_v I__8904 (
            .O(N__39082),
            .I(N__39044));
    LocalMux I__8903 (
            .O(N__39079),
            .I(N__39037));
    LocalMux I__8902 (
            .O(N__39072),
            .I(N__39037));
    Span4Mux_v I__8901 (
            .O(N__39067),
            .I(N__39037));
    Span4Mux_h I__8900 (
            .O(N__39060),
            .I(N__39034));
    CascadeMux I__8899 (
            .O(N__39059),
            .I(N__39031));
    LocalMux I__8898 (
            .O(N__39056),
            .I(N__39025));
    LocalMux I__8897 (
            .O(N__39051),
            .I(N__39025));
    Sp12to4 I__8896 (
            .O(N__39044),
            .I(N__39022));
    Span4Mux_h I__8895 (
            .O(N__39037),
            .I(N__39017));
    Span4Mux_v I__8894 (
            .O(N__39034),
            .I(N__39017));
    InMux I__8893 (
            .O(N__39031),
            .I(N__39013));
    InMux I__8892 (
            .O(N__39030),
            .I(N__39010));
    Span12Mux_h I__8891 (
            .O(N__39025),
            .I(N__39007));
    Span12Mux_v I__8890 (
            .O(N__39022),
            .I(N__39004));
    Span4Mux_v I__8889 (
            .O(N__39017),
            .I(N__39001));
    InMux I__8888 (
            .O(N__39016),
            .I(N__38998));
    LocalMux I__8887 (
            .O(N__39013),
            .I(rx_data_ready));
    LocalMux I__8886 (
            .O(N__39010),
            .I(rx_data_ready));
    Odrv12 I__8885 (
            .O(N__39007),
            .I(rx_data_ready));
    Odrv12 I__8884 (
            .O(N__39004),
            .I(rx_data_ready));
    Odrv4 I__8883 (
            .O(N__39001),
            .I(rx_data_ready));
    LocalMux I__8882 (
            .O(N__38998),
            .I(rx_data_ready));
    InMux I__8881 (
            .O(N__38985),
            .I(N__38982));
    LocalMux I__8880 (
            .O(N__38982),
            .I(N__38979));
    Span4Mux_v I__8879 (
            .O(N__38979),
            .I(N__38974));
    InMux I__8878 (
            .O(N__38978),
            .I(N__38971));
    InMux I__8877 (
            .O(N__38977),
            .I(N__38968));
    Span4Mux_h I__8876 (
            .O(N__38974),
            .I(N__38964));
    LocalMux I__8875 (
            .O(N__38971),
            .I(N__38961));
    LocalMux I__8874 (
            .O(N__38968),
            .I(N__38958));
    InMux I__8873 (
            .O(N__38967),
            .I(N__38955));
    Span4Mux_h I__8872 (
            .O(N__38964),
            .I(N__38950));
    Span4Mux_h I__8871 (
            .O(N__38961),
            .I(N__38950));
    Sp12to4 I__8870 (
            .O(N__38958),
            .I(N__38947));
    LocalMux I__8869 (
            .O(N__38955),
            .I(data_in_3_2));
    Odrv4 I__8868 (
            .O(N__38950),
            .I(data_in_3_2));
    Odrv12 I__8867 (
            .O(N__38947),
            .I(data_in_3_2));
    InMux I__8866 (
            .O(N__38940),
            .I(N__38936));
    InMux I__8865 (
            .O(N__38939),
            .I(N__38933));
    LocalMux I__8864 (
            .O(N__38936),
            .I(N__38929));
    LocalMux I__8863 (
            .O(N__38933),
            .I(N__38926));
    InMux I__8862 (
            .O(N__38932),
            .I(N__38923));
    Span4Mux_v I__8861 (
            .O(N__38929),
            .I(N__38919));
    Span4Mux_v I__8860 (
            .O(N__38926),
            .I(N__38914));
    LocalMux I__8859 (
            .O(N__38923),
            .I(N__38914));
    InMux I__8858 (
            .O(N__38922),
            .I(N__38911));
    Span4Mux_h I__8857 (
            .O(N__38919),
            .I(N__38906));
    Span4Mux_h I__8856 (
            .O(N__38914),
            .I(N__38906));
    LocalMux I__8855 (
            .O(N__38911),
            .I(data_in_2_2));
    Odrv4 I__8854 (
            .O(N__38906),
            .I(data_in_2_2));
    InMux I__8853 (
            .O(N__38901),
            .I(N__38896));
    InMux I__8852 (
            .O(N__38900),
            .I(N__38893));
    CascadeMux I__8851 (
            .O(N__38899),
            .I(N__38889));
    LocalMux I__8850 (
            .O(N__38896),
            .I(N__38886));
    LocalMux I__8849 (
            .O(N__38893),
            .I(N__38882));
    InMux I__8848 (
            .O(N__38892),
            .I(N__38879));
    InMux I__8847 (
            .O(N__38889),
            .I(N__38876));
    Span4Mux_v I__8846 (
            .O(N__38886),
            .I(N__38873));
    InMux I__8845 (
            .O(N__38885),
            .I(N__38870));
    Span4Mux_v I__8844 (
            .O(N__38882),
            .I(N__38867));
    LocalMux I__8843 (
            .O(N__38879),
            .I(N__38864));
    LocalMux I__8842 (
            .O(N__38876),
            .I(\c0.data_in_frame_1_3 ));
    Odrv4 I__8841 (
            .O(N__38873),
            .I(\c0.data_in_frame_1_3 ));
    LocalMux I__8840 (
            .O(N__38870),
            .I(\c0.data_in_frame_1_3 ));
    Odrv4 I__8839 (
            .O(N__38867),
            .I(\c0.data_in_frame_1_3 ));
    Odrv4 I__8838 (
            .O(N__38864),
            .I(\c0.data_in_frame_1_3 ));
    CascadeMux I__8837 (
            .O(N__38853),
            .I(N__38850));
    InMux I__8836 (
            .O(N__38850),
            .I(N__38846));
    InMux I__8835 (
            .O(N__38849),
            .I(N__38843));
    LocalMux I__8834 (
            .O(N__38846),
            .I(N__38840));
    LocalMux I__8833 (
            .O(N__38843),
            .I(N__38835));
    Span4Mux_v I__8832 (
            .O(N__38840),
            .I(N__38835));
    Odrv4 I__8831 (
            .O(N__38835),
            .I(\c0.data_in_frame_5_4 ));
    InMux I__8830 (
            .O(N__38832),
            .I(N__38829));
    LocalMux I__8829 (
            .O(N__38829),
            .I(N__38824));
    InMux I__8828 (
            .O(N__38828),
            .I(N__38819));
    InMux I__8827 (
            .O(N__38827),
            .I(N__38816));
    Span4Mux_h I__8826 (
            .O(N__38824),
            .I(N__38813));
    InMux I__8825 (
            .O(N__38823),
            .I(N__38808));
    InMux I__8824 (
            .O(N__38822),
            .I(N__38808));
    LocalMux I__8823 (
            .O(N__38819),
            .I(N__38803));
    LocalMux I__8822 (
            .O(N__38816),
            .I(N__38803));
    Odrv4 I__8821 (
            .O(N__38813),
            .I(\c0.data_in_frame_1_2 ));
    LocalMux I__8820 (
            .O(N__38808),
            .I(\c0.data_in_frame_1_2 ));
    Odrv4 I__8819 (
            .O(N__38803),
            .I(\c0.data_in_frame_1_2 ));
    InMux I__8818 (
            .O(N__38796),
            .I(N__38793));
    LocalMux I__8817 (
            .O(N__38793),
            .I(\c0.n21_adj_2357 ));
    InMux I__8816 (
            .O(N__38790),
            .I(N__38786));
    InMux I__8815 (
            .O(N__38789),
            .I(N__38783));
    LocalMux I__8814 (
            .O(N__38786),
            .I(\c0.delay_counter_12 ));
    LocalMux I__8813 (
            .O(N__38783),
            .I(\c0.delay_counter_12 ));
    InMux I__8812 (
            .O(N__38778),
            .I(N__38775));
    LocalMux I__8811 (
            .O(N__38775),
            .I(\c0.n16_adj_2212 ));
    InMux I__8810 (
            .O(N__38772),
            .I(N__38766));
    InMux I__8809 (
            .O(N__38771),
            .I(N__38766));
    LocalMux I__8808 (
            .O(N__38766),
            .I(\c0.delay_counter_2 ));
    InMux I__8807 (
            .O(N__38763),
            .I(N__38760));
    LocalMux I__8806 (
            .O(N__38760),
            .I(\c0.n26 ));
    InMux I__8805 (
            .O(N__38757),
            .I(N__38753));
    InMux I__8804 (
            .O(N__38756),
            .I(N__38750));
    LocalMux I__8803 (
            .O(N__38753),
            .I(\c0.delay_counter_0 ));
    LocalMux I__8802 (
            .O(N__38750),
            .I(\c0.delay_counter_0 ));
    InMux I__8801 (
            .O(N__38745),
            .I(N__38741));
    InMux I__8800 (
            .O(N__38744),
            .I(N__38738));
    LocalMux I__8799 (
            .O(N__38741),
            .I(\c0.delay_counter_6 ));
    LocalMux I__8798 (
            .O(N__38738),
            .I(\c0.delay_counter_6 ));
    InMux I__8797 (
            .O(N__38733),
            .I(N__38730));
    LocalMux I__8796 (
            .O(N__38730),
            .I(\c0.n22_adj_2390 ));
    InMux I__8795 (
            .O(N__38727),
            .I(N__38721));
    InMux I__8794 (
            .O(N__38726),
            .I(N__38721));
    LocalMux I__8793 (
            .O(N__38721),
            .I(\c0.delay_counter_10 ));
    InMux I__8792 (
            .O(N__38718),
            .I(N__38715));
    LocalMux I__8791 (
            .O(N__38715),
            .I(\c0.n18_adj_2220 ));
    CascadeMux I__8790 (
            .O(N__38712),
            .I(N__38708));
    InMux I__8789 (
            .O(N__38711),
            .I(N__38703));
    InMux I__8788 (
            .O(N__38708),
            .I(N__38703));
    LocalMux I__8787 (
            .O(N__38703),
            .I(\c0.delay_counter_13 ));
    InMux I__8786 (
            .O(N__38700),
            .I(N__38697));
    LocalMux I__8785 (
            .O(N__38697),
            .I(\c0.n15_adj_2211 ));
    InMux I__8784 (
            .O(N__38694),
            .I(N__38691));
    LocalMux I__8783 (
            .O(N__38691),
            .I(N__38687));
    InMux I__8782 (
            .O(N__38690),
            .I(N__38684));
    Span4Mux_h I__8781 (
            .O(N__38687),
            .I(N__38681));
    LocalMux I__8780 (
            .O(N__38684),
            .I(r_Tx_Data_5));
    Odrv4 I__8779 (
            .O(N__38681),
            .I(r_Tx_Data_5));
    InMux I__8778 (
            .O(N__38676),
            .I(N__38672));
    InMux I__8777 (
            .O(N__38675),
            .I(N__38669));
    LocalMux I__8776 (
            .O(N__38672),
            .I(\c0.delay_counter_11 ));
    LocalMux I__8775 (
            .O(N__38669),
            .I(\c0.delay_counter_11 ));
    InMux I__8774 (
            .O(N__38664),
            .I(N__38657));
    CascadeMux I__8773 (
            .O(N__38663),
            .I(N__38654));
    InMux I__8772 (
            .O(N__38662),
            .I(N__38649));
    CascadeMux I__8771 (
            .O(N__38661),
            .I(N__38643));
    CascadeMux I__8770 (
            .O(N__38660),
            .I(N__38640));
    LocalMux I__8769 (
            .O(N__38657),
            .I(N__38632));
    InMux I__8768 (
            .O(N__38654),
            .I(N__38625));
    InMux I__8767 (
            .O(N__38653),
            .I(N__38625));
    InMux I__8766 (
            .O(N__38652),
            .I(N__38625));
    LocalMux I__8765 (
            .O(N__38649),
            .I(N__38622));
    InMux I__8764 (
            .O(N__38648),
            .I(N__38615));
    InMux I__8763 (
            .O(N__38647),
            .I(N__38615));
    InMux I__8762 (
            .O(N__38646),
            .I(N__38615));
    InMux I__8761 (
            .O(N__38643),
            .I(N__38608));
    InMux I__8760 (
            .O(N__38640),
            .I(N__38608));
    InMux I__8759 (
            .O(N__38639),
            .I(N__38608));
    InMux I__8758 (
            .O(N__38638),
            .I(N__38605));
    InMux I__8757 (
            .O(N__38637),
            .I(N__38598));
    InMux I__8756 (
            .O(N__38636),
            .I(N__38598));
    InMux I__8755 (
            .O(N__38635),
            .I(N__38598));
    Span4Mux_h I__8754 (
            .O(N__38632),
            .I(N__38595));
    LocalMux I__8753 (
            .O(N__38625),
            .I(\c0.n9453 ));
    Odrv4 I__8752 (
            .O(N__38622),
            .I(\c0.n9453 ));
    LocalMux I__8751 (
            .O(N__38615),
            .I(\c0.n9453 ));
    LocalMux I__8750 (
            .O(N__38608),
            .I(\c0.n9453 ));
    LocalMux I__8749 (
            .O(N__38605),
            .I(\c0.n9453 ));
    LocalMux I__8748 (
            .O(N__38598),
            .I(\c0.n9453 ));
    Odrv4 I__8747 (
            .O(N__38595),
            .I(\c0.n9453 ));
    InMux I__8746 (
            .O(N__38580),
            .I(N__38571));
    InMux I__8745 (
            .O(N__38579),
            .I(N__38571));
    InMux I__8744 (
            .O(N__38578),
            .I(N__38571));
    LocalMux I__8743 (
            .O(N__38571),
            .I(N__38555));
    InMux I__8742 (
            .O(N__38570),
            .I(N__38552));
    InMux I__8741 (
            .O(N__38569),
            .I(N__38543));
    InMux I__8740 (
            .O(N__38568),
            .I(N__38543));
    InMux I__8739 (
            .O(N__38567),
            .I(N__38543));
    InMux I__8738 (
            .O(N__38566),
            .I(N__38543));
    InMux I__8737 (
            .O(N__38565),
            .I(N__38534));
    InMux I__8736 (
            .O(N__38564),
            .I(N__38534));
    InMux I__8735 (
            .O(N__38563),
            .I(N__38534));
    InMux I__8734 (
            .O(N__38562),
            .I(N__38534));
    InMux I__8733 (
            .O(N__38561),
            .I(N__38527));
    InMux I__8732 (
            .O(N__38560),
            .I(N__38527));
    InMux I__8731 (
            .O(N__38559),
            .I(N__38527));
    InMux I__8730 (
            .O(N__38558),
            .I(N__38524));
    Odrv4 I__8729 (
            .O(N__38555),
            .I(\c0.n16267 ));
    LocalMux I__8728 (
            .O(N__38552),
            .I(\c0.n16267 ));
    LocalMux I__8727 (
            .O(N__38543),
            .I(\c0.n16267 ));
    LocalMux I__8726 (
            .O(N__38534),
            .I(\c0.n16267 ));
    LocalMux I__8725 (
            .O(N__38527),
            .I(\c0.n16267 ));
    LocalMux I__8724 (
            .O(N__38524),
            .I(\c0.n16267 ));
    InMux I__8723 (
            .O(N__38511),
            .I(N__38508));
    LocalMux I__8722 (
            .O(N__38508),
            .I(\c0.n17_adj_2219 ));
    InMux I__8721 (
            .O(N__38505),
            .I(N__38501));
    InMux I__8720 (
            .O(N__38504),
            .I(N__38498));
    LocalMux I__8719 (
            .O(N__38501),
            .I(\c0.delay_counter_8 ));
    LocalMux I__8718 (
            .O(N__38498),
            .I(\c0.delay_counter_8 ));
    InMux I__8717 (
            .O(N__38493),
            .I(N__38489));
    InMux I__8716 (
            .O(N__38492),
            .I(N__38486));
    LocalMux I__8715 (
            .O(N__38489),
            .I(\c0.delay_counter_3 ));
    LocalMux I__8714 (
            .O(N__38486),
            .I(\c0.delay_counter_3 ));
    InMux I__8713 (
            .O(N__38481),
            .I(N__38478));
    LocalMux I__8712 (
            .O(N__38478),
            .I(\c0.n18_adj_2388 ));
    InMux I__8711 (
            .O(N__38475),
            .I(N__38472));
    LocalMux I__8710 (
            .O(N__38472),
            .I(n17765));
    CascadeMux I__8709 (
            .O(N__38469),
            .I(n17392_cascade_));
    InMux I__8708 (
            .O(N__38466),
            .I(N__38463));
    LocalMux I__8707 (
            .O(N__38463),
            .I(n17416));
    InMux I__8706 (
            .O(N__38460),
            .I(N__38457));
    LocalMux I__8705 (
            .O(N__38457),
            .I(\c0.n20_adj_2255 ));
    InMux I__8704 (
            .O(N__38454),
            .I(N__38450));
    InMux I__8703 (
            .O(N__38453),
            .I(N__38447));
    LocalMux I__8702 (
            .O(N__38450),
            .I(\c0.delay_counter_7 ));
    LocalMux I__8701 (
            .O(N__38447),
            .I(\c0.delay_counter_7 ));
    CascadeMux I__8700 (
            .O(N__38442),
            .I(N__38439));
    InMux I__8699 (
            .O(N__38439),
            .I(N__38435));
    InMux I__8698 (
            .O(N__38438),
            .I(N__38432));
    LocalMux I__8697 (
            .O(N__38435),
            .I(\c0.delay_counter_5 ));
    LocalMux I__8696 (
            .O(N__38432),
            .I(\c0.delay_counter_5 ));
    CascadeMux I__8695 (
            .O(N__38427),
            .I(\c0.n24_adj_2389_cascade_ ));
    InMux I__8694 (
            .O(N__38424),
            .I(N__38421));
    LocalMux I__8693 (
            .O(N__38421),
            .I(N__38418));
    Odrv4 I__8692 (
            .O(N__38418),
            .I(n17327));
    CascadeMux I__8691 (
            .O(N__38415),
            .I(N__38411));
    InMux I__8690 (
            .O(N__38414),
            .I(N__38408));
    InMux I__8689 (
            .O(N__38411),
            .I(N__38405));
    LocalMux I__8688 (
            .O(N__38408),
            .I(N__38402));
    LocalMux I__8687 (
            .O(N__38405),
            .I(\c0.delay_counter_1 ));
    Odrv4 I__8686 (
            .O(N__38402),
            .I(\c0.delay_counter_1 ));
    CascadeMux I__8685 (
            .O(N__38397),
            .I(N__38394));
    InMux I__8684 (
            .O(N__38394),
            .I(N__38390));
    CascadeMux I__8683 (
            .O(N__38393),
            .I(N__38387));
    LocalMux I__8682 (
            .O(N__38390),
            .I(N__38384));
    InMux I__8681 (
            .O(N__38387),
            .I(N__38381));
    Odrv4 I__8680 (
            .O(N__38384),
            .I(\c0.delay_counter_9 ));
    LocalMux I__8679 (
            .O(N__38381),
            .I(\c0.delay_counter_9 ));
    InMux I__8678 (
            .O(N__38376),
            .I(N__38373));
    LocalMux I__8677 (
            .O(N__38373),
            .I(\c0.n26_adj_2391 ));
    CascadeMux I__8676 (
            .O(N__38370),
            .I(N__38366));
    InMux I__8675 (
            .O(N__38369),
            .I(N__38361));
    InMux I__8674 (
            .O(N__38366),
            .I(N__38361));
    LocalMux I__8673 (
            .O(N__38361),
            .I(\c0.delay_counter_4 ));
    CascadeMux I__8672 (
            .O(N__38358),
            .I(\c0.n9453_cascade_ ));
    InMux I__8671 (
            .O(N__38355),
            .I(N__38352));
    LocalMux I__8670 (
            .O(N__38352),
            .I(\c0.n24_adj_2342 ));
    InMux I__8669 (
            .O(N__38349),
            .I(N__38346));
    LocalMux I__8668 (
            .O(N__38346),
            .I(\c0.n453 ));
    InMux I__8667 (
            .O(N__38343),
            .I(N__38337));
    InMux I__8666 (
            .O(N__38342),
            .I(N__38332));
    InMux I__8665 (
            .O(N__38341),
            .I(N__38332));
    InMux I__8664 (
            .O(N__38340),
            .I(N__38329));
    LocalMux I__8663 (
            .O(N__38337),
            .I(n4_adj_2414));
    LocalMux I__8662 (
            .O(N__38332),
            .I(n4_adj_2414));
    LocalMux I__8661 (
            .O(N__38329),
            .I(n4_adj_2414));
    CascadeMux I__8660 (
            .O(N__38322),
            .I(N__38319));
    InMux I__8659 (
            .O(N__38319),
            .I(N__38316));
    LocalMux I__8658 (
            .O(N__38316),
            .I(N__38313));
    Odrv4 I__8657 (
            .O(N__38313),
            .I(\c0.n19 ));
    CascadeMux I__8656 (
            .O(N__38310),
            .I(n9524_cascade_));
    CascadeMux I__8655 (
            .O(N__38307),
            .I(\c0.n16267_cascade_ ));
    InMux I__8654 (
            .O(N__38304),
            .I(N__38301));
    LocalMux I__8653 (
            .O(N__38301),
            .I(\c0.n445 ));
    CascadeMux I__8652 (
            .O(N__38298),
            .I(N__38295));
    InMux I__8651 (
            .O(N__38295),
            .I(N__38292));
    LocalMux I__8650 (
            .O(N__38292),
            .I(\c0.n23_adj_2314 ));
    CascadeMux I__8649 (
            .O(N__38289),
            .I(N__38286));
    InMux I__8648 (
            .O(N__38286),
            .I(N__38283));
    LocalMux I__8647 (
            .O(N__38283),
            .I(\c0.n28 ));
    InMux I__8646 (
            .O(N__38280),
            .I(N__38277));
    LocalMux I__8645 (
            .O(N__38277),
            .I(n5_adj_2407));
    CascadeMux I__8644 (
            .O(N__38274),
            .I(N__38271));
    InMux I__8643 (
            .O(N__38271),
            .I(N__38268));
    LocalMux I__8642 (
            .O(N__38268),
            .I(\c0.n5_adj_2141 ));
    InMux I__8641 (
            .O(N__38265),
            .I(N__38261));
    InMux I__8640 (
            .O(N__38264),
            .I(N__38258));
    LocalMux I__8639 (
            .O(N__38261),
            .I(r_Tx_Data_2));
    LocalMux I__8638 (
            .O(N__38258),
            .I(r_Tx_Data_2));
    InMux I__8637 (
            .O(N__38253),
            .I(N__38250));
    LocalMux I__8636 (
            .O(N__38250),
            .I(N__38246));
    InMux I__8635 (
            .O(N__38249),
            .I(N__38243));
    Span4Mux_v I__8634 (
            .O(N__38246),
            .I(N__38240));
    LocalMux I__8633 (
            .O(N__38243),
            .I(r_Tx_Data_4));
    Odrv4 I__8632 (
            .O(N__38240),
            .I(r_Tx_Data_4));
    CascadeMux I__8631 (
            .O(N__38235),
            .I(n18196_cascade_));
    InMux I__8630 (
            .O(N__38232),
            .I(N__38229));
    LocalMux I__8629 (
            .O(N__38229),
            .I(n18199));
    InMux I__8628 (
            .O(N__38226),
            .I(N__38223));
    LocalMux I__8627 (
            .O(N__38223),
            .I(\c0.tx.n31 ));
    InMux I__8626 (
            .O(N__38220),
            .I(N__38217));
    LocalMux I__8625 (
            .O(N__38217),
            .I(n17759));
    InMux I__8624 (
            .O(N__38214),
            .I(N__38211));
    LocalMux I__8623 (
            .O(N__38211),
            .I(N__38208));
    Odrv4 I__8622 (
            .O(N__38208),
            .I(n17664));
    InMux I__8621 (
            .O(N__38205),
            .I(N__38202));
    LocalMux I__8620 (
            .O(N__38202),
            .I(N__38199));
    Odrv4 I__8619 (
            .O(N__38199),
            .I(\c0.n18166 ));
    InMux I__8618 (
            .O(N__38196),
            .I(N__38193));
    LocalMux I__8617 (
            .O(N__38193),
            .I(N__38190));
    Span4Mux_v I__8616 (
            .O(N__38190),
            .I(N__38187));
    Odrv4 I__8615 (
            .O(N__38187),
            .I(\c0.n2_adj_2145 ));
    CascadeMux I__8614 (
            .O(N__38184),
            .I(N__38181));
    InMux I__8613 (
            .O(N__38181),
            .I(N__38178));
    LocalMux I__8612 (
            .O(N__38178),
            .I(N__38175));
    Span4Mux_v I__8611 (
            .O(N__38175),
            .I(N__38172));
    Span4Mux_h I__8610 (
            .O(N__38172),
            .I(N__38169));
    Odrv4 I__8609 (
            .O(N__38169),
            .I(\c0.n17701 ));
    InMux I__8608 (
            .O(N__38166),
            .I(N__38163));
    LocalMux I__8607 (
            .O(N__38163),
            .I(N__38160));
    Odrv4 I__8606 (
            .O(N__38160),
            .I(n18169));
    InMux I__8605 (
            .O(N__38157),
            .I(N__38154));
    LocalMux I__8604 (
            .O(N__38154),
            .I(N__38150));
    CascadeMux I__8603 (
            .O(N__38153),
            .I(N__38147));
    Span4Mux_v I__8602 (
            .O(N__38150),
            .I(N__38144));
    InMux I__8601 (
            .O(N__38147),
            .I(N__38141));
    Odrv4 I__8600 (
            .O(N__38144),
            .I(rand_setpoint_7));
    LocalMux I__8599 (
            .O(N__38141),
            .I(rand_setpoint_7));
    CascadeMux I__8598 (
            .O(N__38136),
            .I(N__38132));
    InMux I__8597 (
            .O(N__38135),
            .I(N__38127));
    InMux I__8596 (
            .O(N__38132),
            .I(N__38127));
    LocalMux I__8595 (
            .O(N__38127),
            .I(data_out_0_0));
    InMux I__8594 (
            .O(N__38124),
            .I(N__38121));
    LocalMux I__8593 (
            .O(N__38121),
            .I(N__38117));
    CascadeMux I__8592 (
            .O(N__38120),
            .I(N__38114));
    Span4Mux_v I__8591 (
            .O(N__38117),
            .I(N__38111));
    InMux I__8590 (
            .O(N__38114),
            .I(N__38108));
    Odrv4 I__8589 (
            .O(N__38111),
            .I(rand_setpoint_16));
    LocalMux I__8588 (
            .O(N__38108),
            .I(rand_setpoint_16));
    InMux I__8587 (
            .O(N__38103),
            .I(N__38100));
    LocalMux I__8586 (
            .O(N__38100),
            .I(N__38096));
    CascadeMux I__8585 (
            .O(N__38099),
            .I(N__38093));
    Span4Mux_v I__8584 (
            .O(N__38096),
            .I(N__38090));
    InMux I__8583 (
            .O(N__38093),
            .I(N__38087));
    Odrv4 I__8582 (
            .O(N__38090),
            .I(rand_setpoint_15));
    LocalMux I__8581 (
            .O(N__38087),
            .I(rand_setpoint_15));
    CascadeMux I__8580 (
            .O(N__38082),
            .I(N__38079));
    InMux I__8579 (
            .O(N__38079),
            .I(N__38076));
    LocalMux I__8578 (
            .O(N__38076),
            .I(n10_adj_2450));
    CascadeMux I__8577 (
            .O(N__38073),
            .I(n10_adj_2411_cascade_));
    CascadeMux I__8576 (
            .O(N__38070),
            .I(N__38066));
    InMux I__8575 (
            .O(N__38069),
            .I(N__38062));
    InMux I__8574 (
            .O(N__38066),
            .I(N__38059));
    InMux I__8573 (
            .O(N__38065),
            .I(N__38056));
    LocalMux I__8572 (
            .O(N__38062),
            .I(N__38053));
    LocalMux I__8571 (
            .O(N__38059),
            .I(N__38050));
    LocalMux I__8570 (
            .O(N__38056),
            .I(\c0.FRAME_MATCHER_state_27 ));
    Odrv4 I__8569 (
            .O(N__38053),
            .I(\c0.FRAME_MATCHER_state_27 ));
    Odrv12 I__8568 (
            .O(N__38050),
            .I(\c0.FRAME_MATCHER_state_27 ));
    SRMux I__8567 (
            .O(N__38043),
            .I(N__38040));
    LocalMux I__8566 (
            .O(N__38040),
            .I(N__38037));
    Span4Mux_h I__8565 (
            .O(N__38037),
            .I(N__38034));
    Odrv4 I__8564 (
            .O(N__38034),
            .I(\c0.n16718 ));
    InMux I__8563 (
            .O(N__38031),
            .I(N__38028));
    LocalMux I__8562 (
            .O(N__38028),
            .I(N__38025));
    Span4Mux_h I__8561 (
            .O(N__38025),
            .I(N__38022));
    Span4Mux_h I__8560 (
            .O(N__38022),
            .I(N__38019));
    Span4Mux_h I__8559 (
            .O(N__38019),
            .I(N__38015));
    CascadeMux I__8558 (
            .O(N__38018),
            .I(N__38012));
    Span4Mux_h I__8557 (
            .O(N__38015),
            .I(N__38009));
    InMux I__8556 (
            .O(N__38012),
            .I(N__38006));
    Odrv4 I__8555 (
            .O(N__38009),
            .I(rand_setpoint_0));
    LocalMux I__8554 (
            .O(N__38006),
            .I(rand_setpoint_0));
    InMux I__8553 (
            .O(N__38001),
            .I(N__37998));
    LocalMux I__8552 (
            .O(N__37998),
            .I(n2));
    InMux I__8551 (
            .O(N__37995),
            .I(N__37991));
    InMux I__8550 (
            .O(N__37994),
            .I(N__37988));
    LocalMux I__8549 (
            .O(N__37991),
            .I(data_out_2_0));
    LocalMux I__8548 (
            .O(N__37988),
            .I(data_out_2_0));
    InMux I__8547 (
            .O(N__37983),
            .I(N__37980));
    LocalMux I__8546 (
            .O(N__37980),
            .I(N__37977));
    Span4Mux_v I__8545 (
            .O(N__37977),
            .I(N__37974));
    Span4Mux_v I__8544 (
            .O(N__37974),
            .I(N__37970));
    InMux I__8543 (
            .O(N__37973),
            .I(N__37967));
    Odrv4 I__8542 (
            .O(N__37970),
            .I(n4_adj_2427));
    LocalMux I__8541 (
            .O(N__37967),
            .I(n4_adj_2427));
    InMux I__8540 (
            .O(N__37962),
            .I(N__37956));
    InMux I__8539 (
            .O(N__37961),
            .I(N__37956));
    LocalMux I__8538 (
            .O(N__37956),
            .I(N__37953));
    Odrv12 I__8537 (
            .O(N__37953),
            .I(n4_adj_2416));
    InMux I__8536 (
            .O(N__37950),
            .I(N__37938));
    InMux I__8535 (
            .O(N__37949),
            .I(N__37938));
    InMux I__8534 (
            .O(N__37948),
            .I(N__37938));
    InMux I__8533 (
            .O(N__37947),
            .I(N__37938));
    LocalMux I__8532 (
            .O(N__37938),
            .I(N__37935));
    Span12Mux_h I__8531 (
            .O(N__37935),
            .I(N__37930));
    InMux I__8530 (
            .O(N__37934),
            .I(N__37925));
    InMux I__8529 (
            .O(N__37933),
            .I(N__37925));
    Odrv12 I__8528 (
            .O(N__37930),
            .I(r_Bit_Index_1_adj_2436));
    LocalMux I__8527 (
            .O(N__37925),
            .I(r_Bit_Index_1_adj_2436));
    InMux I__8526 (
            .O(N__37920),
            .I(N__37908));
    InMux I__8525 (
            .O(N__37919),
            .I(N__37908));
    InMux I__8524 (
            .O(N__37918),
            .I(N__37908));
    InMux I__8523 (
            .O(N__37917),
            .I(N__37908));
    LocalMux I__8522 (
            .O(N__37908),
            .I(N__37904));
    CascadeMux I__8521 (
            .O(N__37907),
            .I(N__37899));
    Sp12to4 I__8520 (
            .O(N__37904),
            .I(N__37896));
    InMux I__8519 (
            .O(N__37903),
            .I(N__37891));
    InMux I__8518 (
            .O(N__37902),
            .I(N__37891));
    InMux I__8517 (
            .O(N__37899),
            .I(N__37888));
    Span12Mux_v I__8516 (
            .O(N__37896),
            .I(N__37885));
    LocalMux I__8515 (
            .O(N__37891),
            .I(N__37882));
    LocalMux I__8514 (
            .O(N__37888),
            .I(r_Bit_Index_2_adj_2435));
    Odrv12 I__8513 (
            .O(N__37885),
            .I(r_Bit_Index_2_adj_2435));
    Odrv4 I__8512 (
            .O(N__37882),
            .I(r_Bit_Index_2_adj_2435));
    InMux I__8511 (
            .O(N__37875),
            .I(N__37872));
    LocalMux I__8510 (
            .O(N__37872),
            .I(N__37869));
    Span4Mux_v I__8509 (
            .O(N__37869),
            .I(N__37865));
    InMux I__8508 (
            .O(N__37868),
            .I(N__37862));
    Span4Mux_h I__8507 (
            .O(N__37865),
            .I(N__37857));
    LocalMux I__8506 (
            .O(N__37862),
            .I(N__37857));
    Span4Mux_v I__8505 (
            .O(N__37857),
            .I(N__37854));
    Span4Mux_h I__8504 (
            .O(N__37854),
            .I(N__37848));
    InMux I__8503 (
            .O(N__37853),
            .I(N__37841));
    InMux I__8502 (
            .O(N__37852),
            .I(N__37841));
    InMux I__8501 (
            .O(N__37851),
            .I(N__37841));
    Odrv4 I__8500 (
            .O(N__37848),
            .I(r_Bit_Index_0));
    LocalMux I__8499 (
            .O(N__37841),
            .I(r_Bit_Index_0));
    InMux I__8498 (
            .O(N__37836),
            .I(N__37833));
    LocalMux I__8497 (
            .O(N__37833),
            .I(N__37830));
    Span4Mux_h I__8496 (
            .O(N__37830),
            .I(N__37826));
    InMux I__8495 (
            .O(N__37829),
            .I(N__37823));
    Span4Mux_v I__8494 (
            .O(N__37826),
            .I(N__37818));
    LocalMux I__8493 (
            .O(N__37823),
            .I(N__37818));
    Span4Mux_h I__8492 (
            .O(N__37818),
            .I(N__37815));
    Span4Mux_v I__8491 (
            .O(N__37815),
            .I(N__37812));
    Odrv4 I__8490 (
            .O(N__37812),
            .I(\c0.rx.n10158 ));
    InMux I__8489 (
            .O(N__37809),
            .I(N__37805));
    InMux I__8488 (
            .O(N__37808),
            .I(N__37802));
    LocalMux I__8487 (
            .O(N__37805),
            .I(N__37797));
    LocalMux I__8486 (
            .O(N__37802),
            .I(N__37797));
    Span4Mux_h I__8485 (
            .O(N__37797),
            .I(N__37794));
    Span4Mux_h I__8484 (
            .O(N__37794),
            .I(N__37790));
    CascadeMux I__8483 (
            .O(N__37793),
            .I(N__37787));
    Span4Mux_v I__8482 (
            .O(N__37790),
            .I(N__37784));
    InMux I__8481 (
            .O(N__37787),
            .I(N__37781));
    Span4Mux_h I__8480 (
            .O(N__37784),
            .I(N__37778));
    LocalMux I__8479 (
            .O(N__37781),
            .I(\c0.FRAME_MATCHER_state_16 ));
    Odrv4 I__8478 (
            .O(N__37778),
            .I(\c0.FRAME_MATCHER_state_16 ));
    InMux I__8477 (
            .O(N__37773),
            .I(N__37770));
    LocalMux I__8476 (
            .O(N__37770),
            .I(\c0.n48 ));
    InMux I__8475 (
            .O(N__37767),
            .I(N__37758));
    InMux I__8474 (
            .O(N__37766),
            .I(N__37758));
    InMux I__8473 (
            .O(N__37765),
            .I(N__37758));
    LocalMux I__8472 (
            .O(N__37758),
            .I(\c0.FRAME_MATCHER_state_30 ));
    SRMux I__8471 (
            .O(N__37755),
            .I(N__37752));
    LocalMux I__8470 (
            .O(N__37752),
            .I(N__37749));
    Odrv4 I__8469 (
            .O(N__37749),
            .I(\c0.n16698 ));
    CascadeMux I__8468 (
            .O(N__37746),
            .I(N__37742));
    InMux I__8467 (
            .O(N__37745),
            .I(N__37737));
    InMux I__8466 (
            .O(N__37742),
            .I(N__37721));
    InMux I__8465 (
            .O(N__37741),
            .I(N__37721));
    InMux I__8464 (
            .O(N__37740),
            .I(N__37721));
    LocalMux I__8463 (
            .O(N__37737),
            .I(N__37718));
    InMux I__8462 (
            .O(N__37736),
            .I(N__37715));
    InMux I__8461 (
            .O(N__37735),
            .I(N__37710));
    InMux I__8460 (
            .O(N__37734),
            .I(N__37710));
    InMux I__8459 (
            .O(N__37733),
            .I(N__37707));
    InMux I__8458 (
            .O(N__37732),
            .I(N__37704));
    InMux I__8457 (
            .O(N__37731),
            .I(N__37701));
    InMux I__8456 (
            .O(N__37730),
            .I(N__37696));
    InMux I__8455 (
            .O(N__37729),
            .I(N__37696));
    InMux I__8454 (
            .O(N__37728),
            .I(N__37693));
    LocalMux I__8453 (
            .O(N__37721),
            .I(N__37687));
    Span4Mux_h I__8452 (
            .O(N__37718),
            .I(N__37682));
    LocalMux I__8451 (
            .O(N__37715),
            .I(N__37682));
    LocalMux I__8450 (
            .O(N__37710),
            .I(N__37671));
    LocalMux I__8449 (
            .O(N__37707),
            .I(N__37671));
    LocalMux I__8448 (
            .O(N__37704),
            .I(N__37671));
    LocalMux I__8447 (
            .O(N__37701),
            .I(N__37671));
    LocalMux I__8446 (
            .O(N__37696),
            .I(N__37671));
    LocalMux I__8445 (
            .O(N__37693),
            .I(N__37668));
    InMux I__8444 (
            .O(N__37692),
            .I(N__37661));
    InMux I__8443 (
            .O(N__37691),
            .I(N__37661));
    InMux I__8442 (
            .O(N__37690),
            .I(N__37661));
    Span4Mux_v I__8441 (
            .O(N__37687),
            .I(N__37658));
    Span4Mux_v I__8440 (
            .O(N__37682),
            .I(N__37649));
    Span4Mux_v I__8439 (
            .O(N__37671),
            .I(N__37649));
    Span4Mux_h I__8438 (
            .O(N__37668),
            .I(N__37649));
    LocalMux I__8437 (
            .O(N__37661),
            .I(N__37649));
    Odrv4 I__8436 (
            .O(N__37658),
            .I(\c0.n15179 ));
    Odrv4 I__8435 (
            .O(N__37649),
            .I(\c0.n15179 ));
    InMux I__8434 (
            .O(N__37644),
            .I(N__37641));
    LocalMux I__8433 (
            .O(N__37641),
            .I(\c0.n17686 ));
    InMux I__8432 (
            .O(N__37638),
            .I(N__37633));
    InMux I__8431 (
            .O(N__37637),
            .I(N__37630));
    InMux I__8430 (
            .O(N__37636),
            .I(N__37627));
    LocalMux I__8429 (
            .O(N__37633),
            .I(N__37624));
    LocalMux I__8428 (
            .O(N__37630),
            .I(N__37619));
    LocalMux I__8427 (
            .O(N__37627),
            .I(N__37616));
    Span4Mux_v I__8426 (
            .O(N__37624),
            .I(N__37613));
    InMux I__8425 (
            .O(N__37623),
            .I(N__37610));
    InMux I__8424 (
            .O(N__37622),
            .I(N__37607));
    Span12Mux_s4_h I__8423 (
            .O(N__37619),
            .I(N__37600));
    Span12Mux_v I__8422 (
            .O(N__37616),
            .I(N__37600));
    Sp12to4 I__8421 (
            .O(N__37613),
            .I(N__37600));
    LocalMux I__8420 (
            .O(N__37610),
            .I(\c0.data_out_frame2_0_4 ));
    LocalMux I__8419 (
            .O(N__37607),
            .I(\c0.data_out_frame2_0_4 ));
    Odrv12 I__8418 (
            .O(N__37600),
            .I(\c0.data_out_frame2_0_4 ));
    InMux I__8417 (
            .O(N__37593),
            .I(N__37590));
    LocalMux I__8416 (
            .O(N__37590),
            .I(\c0.n17688 ));
    InMux I__8415 (
            .O(N__37587),
            .I(N__37584));
    LocalMux I__8414 (
            .O(N__37584),
            .I(N__37577));
    CascadeMux I__8413 (
            .O(N__37583),
            .I(N__37574));
    InMux I__8412 (
            .O(N__37582),
            .I(N__37569));
    InMux I__8411 (
            .O(N__37581),
            .I(N__37569));
    InMux I__8410 (
            .O(N__37580),
            .I(N__37565));
    Span4Mux_h I__8409 (
            .O(N__37577),
            .I(N__37562));
    InMux I__8408 (
            .O(N__37574),
            .I(N__37559));
    LocalMux I__8407 (
            .O(N__37569),
            .I(N__37556));
    InMux I__8406 (
            .O(N__37568),
            .I(N__37553));
    LocalMux I__8405 (
            .O(N__37565),
            .I(N__37550));
    Span4Mux_h I__8404 (
            .O(N__37562),
            .I(N__37547));
    LocalMux I__8403 (
            .O(N__37559),
            .I(N__37542));
    Span12Mux_s11_h I__8402 (
            .O(N__37556),
            .I(N__37542));
    LocalMux I__8401 (
            .O(N__37553),
            .I(N__37539));
    Span4Mux_v I__8400 (
            .O(N__37550),
            .I(N__37536));
    Span4Mux_h I__8399 (
            .O(N__37547),
            .I(N__37533));
    Odrv12 I__8398 (
            .O(N__37542),
            .I(\c0.data_out_frame2_0_3 ));
    Odrv4 I__8397 (
            .O(N__37539),
            .I(\c0.data_out_frame2_0_3 ));
    Odrv4 I__8396 (
            .O(N__37536),
            .I(\c0.data_out_frame2_0_3 ));
    Odrv4 I__8395 (
            .O(N__37533),
            .I(\c0.data_out_frame2_0_3 ));
    InMux I__8394 (
            .O(N__37524),
            .I(N__37520));
    CascadeMux I__8393 (
            .O(N__37523),
            .I(N__37517));
    LocalMux I__8392 (
            .O(N__37520),
            .I(N__37514));
    InMux I__8391 (
            .O(N__37517),
            .I(N__37511));
    Span4Mux_h I__8390 (
            .O(N__37514),
            .I(N__37508));
    LocalMux I__8389 (
            .O(N__37511),
            .I(\c0.data_in_frame_3_7 ));
    Odrv4 I__8388 (
            .O(N__37508),
            .I(\c0.data_in_frame_3_7 ));
    InMux I__8387 (
            .O(N__37503),
            .I(N__37499));
    InMux I__8386 (
            .O(N__37502),
            .I(N__37496));
    LocalMux I__8385 (
            .O(N__37499),
            .I(\c0.n2126 ));
    LocalMux I__8384 (
            .O(N__37496),
            .I(\c0.n2126 ));
    CascadeMux I__8383 (
            .O(N__37491),
            .I(N__37488));
    InMux I__8382 (
            .O(N__37488),
            .I(N__37484));
    InMux I__8381 (
            .O(N__37487),
            .I(N__37481));
    LocalMux I__8380 (
            .O(N__37484),
            .I(N__37478));
    LocalMux I__8379 (
            .O(N__37481),
            .I(\c0.data_in_frame_3_0 ));
    Odrv4 I__8378 (
            .O(N__37478),
            .I(\c0.data_in_frame_3_0 ));
    InMux I__8377 (
            .O(N__37473),
            .I(N__37468));
    InMux I__8376 (
            .O(N__37472),
            .I(N__37465));
    InMux I__8375 (
            .O(N__37471),
            .I(N__37461));
    LocalMux I__8374 (
            .O(N__37468),
            .I(N__37458));
    LocalMux I__8373 (
            .O(N__37465),
            .I(N__37455));
    InMux I__8372 (
            .O(N__37464),
            .I(N__37452));
    LocalMux I__8371 (
            .O(N__37461),
            .I(\c0.n2138 ));
    Odrv4 I__8370 (
            .O(N__37458),
            .I(\c0.n2138 ));
    Odrv4 I__8369 (
            .O(N__37455),
            .I(\c0.n2138 ));
    LocalMux I__8368 (
            .O(N__37452),
            .I(\c0.n2138 ));
    InMux I__8367 (
            .O(N__37443),
            .I(N__37440));
    LocalMux I__8366 (
            .O(N__37440),
            .I(N__37435));
    InMux I__8365 (
            .O(N__37439),
            .I(N__37430));
    InMux I__8364 (
            .O(N__37438),
            .I(N__37430));
    Span4Mux_h I__8363 (
            .O(N__37435),
            .I(N__37427));
    LocalMux I__8362 (
            .O(N__37430),
            .I(\c0.data_in_frame_2_1 ));
    Odrv4 I__8361 (
            .O(N__37427),
            .I(\c0.data_in_frame_2_1 ));
    CascadeMux I__8360 (
            .O(N__37422),
            .I(N__37419));
    InMux I__8359 (
            .O(N__37419),
            .I(N__37414));
    InMux I__8358 (
            .O(N__37418),
            .I(N__37411));
    InMux I__8357 (
            .O(N__37417),
            .I(N__37408));
    LocalMux I__8356 (
            .O(N__37414),
            .I(\c0.data_in_frame_2_2 ));
    LocalMux I__8355 (
            .O(N__37411),
            .I(\c0.data_in_frame_2_2 ));
    LocalMux I__8354 (
            .O(N__37408),
            .I(\c0.data_in_frame_2_2 ));
    CascadeMux I__8353 (
            .O(N__37401),
            .I(\c0.n18_adj_2316_cascade_ ));
    InMux I__8352 (
            .O(N__37398),
            .I(N__37393));
    InMux I__8351 (
            .O(N__37397),
            .I(N__37390));
    InMux I__8350 (
            .O(N__37396),
            .I(N__37386));
    LocalMux I__8349 (
            .O(N__37393),
            .I(N__37381));
    LocalMux I__8348 (
            .O(N__37390),
            .I(N__37381));
    InMux I__8347 (
            .O(N__37389),
            .I(N__37373));
    LocalMux I__8346 (
            .O(N__37386),
            .I(N__37370));
    Span4Mux_h I__8345 (
            .O(N__37381),
            .I(N__37367));
    InMux I__8344 (
            .O(N__37380),
            .I(N__37364));
    InMux I__8343 (
            .O(N__37379),
            .I(N__37357));
    InMux I__8342 (
            .O(N__37378),
            .I(N__37357));
    InMux I__8341 (
            .O(N__37377),
            .I(N__37357));
    InMux I__8340 (
            .O(N__37376),
            .I(N__37354));
    LocalMux I__8339 (
            .O(N__37373),
            .I(\c0.data_in_frame_0_7 ));
    Odrv4 I__8338 (
            .O(N__37370),
            .I(\c0.data_in_frame_0_7 ));
    Odrv4 I__8337 (
            .O(N__37367),
            .I(\c0.data_in_frame_0_7 ));
    LocalMux I__8336 (
            .O(N__37364),
            .I(\c0.data_in_frame_0_7 ));
    LocalMux I__8335 (
            .O(N__37357),
            .I(\c0.data_in_frame_0_7 ));
    LocalMux I__8334 (
            .O(N__37354),
            .I(\c0.data_in_frame_0_7 ));
    InMux I__8333 (
            .O(N__37341),
            .I(N__37338));
    LocalMux I__8332 (
            .O(N__37338),
            .I(\c0.n23_adj_2322 ));
    InMux I__8331 (
            .O(N__37335),
            .I(N__37331));
    CascadeMux I__8330 (
            .O(N__37334),
            .I(N__37328));
    LocalMux I__8329 (
            .O(N__37331),
            .I(N__37324));
    InMux I__8328 (
            .O(N__37328),
            .I(N__37321));
    InMux I__8327 (
            .O(N__37327),
            .I(N__37318));
    Span4Mux_h I__8326 (
            .O(N__37324),
            .I(N__37315));
    LocalMux I__8325 (
            .O(N__37321),
            .I(\c0.FRAME_MATCHER_state_23 ));
    LocalMux I__8324 (
            .O(N__37318),
            .I(\c0.FRAME_MATCHER_state_23 ));
    Odrv4 I__8323 (
            .O(N__37315),
            .I(\c0.FRAME_MATCHER_state_23 ));
    SRMux I__8322 (
            .O(N__37308),
            .I(N__37305));
    LocalMux I__8321 (
            .O(N__37305),
            .I(N__37302));
    Odrv4 I__8320 (
            .O(N__37302),
            .I(\c0.n13381 ));
    InMux I__8319 (
            .O(N__37299),
            .I(N__37296));
    LocalMux I__8318 (
            .O(N__37296),
            .I(N__37292));
    CascadeMux I__8317 (
            .O(N__37295),
            .I(N__37289));
    Span4Mux_v I__8316 (
            .O(N__37292),
            .I(N__37286));
    InMux I__8315 (
            .O(N__37289),
            .I(N__37282));
    Span4Mux_h I__8314 (
            .O(N__37286),
            .I(N__37279));
    InMux I__8313 (
            .O(N__37285),
            .I(N__37276));
    LocalMux I__8312 (
            .O(N__37282),
            .I(\c0.FRAME_MATCHER_state_11 ));
    Odrv4 I__8311 (
            .O(N__37279),
            .I(\c0.FRAME_MATCHER_state_11 ));
    LocalMux I__8310 (
            .O(N__37276),
            .I(\c0.FRAME_MATCHER_state_11 ));
    SRMux I__8309 (
            .O(N__37269),
            .I(N__37266));
    LocalMux I__8308 (
            .O(N__37266),
            .I(N__37263));
    Span4Mux_v I__8307 (
            .O(N__37263),
            .I(N__37260));
    Span4Mux_h I__8306 (
            .O(N__37260),
            .I(N__37257));
    Odrv4 I__8305 (
            .O(N__37257),
            .I(\c0.n8_adj_2333 ));
    CascadeMux I__8304 (
            .O(N__37254),
            .I(N__37249));
    InMux I__8303 (
            .O(N__37253),
            .I(N__37246));
    CascadeMux I__8302 (
            .O(N__37252),
            .I(N__37242));
    InMux I__8301 (
            .O(N__37249),
            .I(N__37239));
    LocalMux I__8300 (
            .O(N__37246),
            .I(N__37235));
    InMux I__8299 (
            .O(N__37245),
            .I(N__37232));
    InMux I__8298 (
            .O(N__37242),
            .I(N__37229));
    LocalMux I__8297 (
            .O(N__37239),
            .I(N__37226));
    InMux I__8296 (
            .O(N__37238),
            .I(N__37223));
    Span12Mux_h I__8295 (
            .O(N__37235),
            .I(N__37220));
    LocalMux I__8294 (
            .O(N__37232),
            .I(N__37215));
    LocalMux I__8293 (
            .O(N__37229),
            .I(N__37215));
    Span4Mux_v I__8292 (
            .O(N__37226),
            .I(N__37212));
    LocalMux I__8291 (
            .O(N__37223),
            .I(data_out_frame2_8_2));
    Odrv12 I__8290 (
            .O(N__37220),
            .I(data_out_frame2_8_2));
    Odrv4 I__8289 (
            .O(N__37215),
            .I(data_out_frame2_8_2));
    Odrv4 I__8288 (
            .O(N__37212),
            .I(data_out_frame2_8_2));
    InMux I__8287 (
            .O(N__37203),
            .I(N__37200));
    LocalMux I__8286 (
            .O(N__37200),
            .I(N__37197));
    Span12Mux_s6_h I__8285 (
            .O(N__37197),
            .I(N__37194));
    Odrv12 I__8284 (
            .O(N__37194),
            .I(\c0.n16 ));
    InMux I__8283 (
            .O(N__37191),
            .I(N__37188));
    LocalMux I__8282 (
            .O(N__37188),
            .I(N__37182));
    InMux I__8281 (
            .O(N__37187),
            .I(N__37179));
    InMux I__8280 (
            .O(N__37186),
            .I(N__37176));
    InMux I__8279 (
            .O(N__37185),
            .I(N__37171));
    Span4Mux_v I__8278 (
            .O(N__37182),
            .I(N__37168));
    LocalMux I__8277 (
            .O(N__37179),
            .I(N__37163));
    LocalMux I__8276 (
            .O(N__37176),
            .I(N__37163));
    InMux I__8275 (
            .O(N__37175),
            .I(N__37160));
    InMux I__8274 (
            .O(N__37174),
            .I(N__37157));
    LocalMux I__8273 (
            .O(N__37171),
            .I(N__37152));
    Span4Mux_h I__8272 (
            .O(N__37168),
            .I(N__37143));
    Span4Mux_v I__8271 (
            .O(N__37163),
            .I(N__37143));
    LocalMux I__8270 (
            .O(N__37160),
            .I(N__37143));
    LocalMux I__8269 (
            .O(N__37157),
            .I(N__37143));
    InMux I__8268 (
            .O(N__37156),
            .I(N__37140));
    InMux I__8267 (
            .O(N__37155),
            .I(N__37137));
    Span4Mux_v I__8266 (
            .O(N__37152),
            .I(N__37132));
    Span4Mux_v I__8265 (
            .O(N__37143),
            .I(N__37132));
    LocalMux I__8264 (
            .O(N__37140),
            .I(N__37129));
    LocalMux I__8263 (
            .O(N__37137),
            .I(N__37126));
    Span4Mux_h I__8262 (
            .O(N__37132),
            .I(N__37123));
    Span4Mux_h I__8261 (
            .O(N__37129),
            .I(N__37120));
    Odrv4 I__8260 (
            .O(N__37126),
            .I(\c0.FRAME_MATCHER_i_0 ));
    Odrv4 I__8259 (
            .O(N__37123),
            .I(\c0.FRAME_MATCHER_i_0 ));
    Odrv4 I__8258 (
            .O(N__37120),
            .I(\c0.FRAME_MATCHER_i_0 ));
    InMux I__8257 (
            .O(N__37113),
            .I(N__37109));
    InMux I__8256 (
            .O(N__37112),
            .I(N__37106));
    LocalMux I__8255 (
            .O(N__37109),
            .I(N__37102));
    LocalMux I__8254 (
            .O(N__37106),
            .I(N__37099));
    InMux I__8253 (
            .O(N__37105),
            .I(N__37096));
    Span4Mux_v I__8252 (
            .O(N__37102),
            .I(N__37089));
    Span4Mux_h I__8251 (
            .O(N__37099),
            .I(N__37089));
    LocalMux I__8250 (
            .O(N__37096),
            .I(N__37089));
    Span4Mux_h I__8249 (
            .O(N__37089),
            .I(N__37085));
    InMux I__8248 (
            .O(N__37088),
            .I(N__37082));
    Span4Mux_v I__8247 (
            .O(N__37085),
            .I(N__37074));
    LocalMux I__8246 (
            .O(N__37082),
            .I(N__37071));
    InMux I__8245 (
            .O(N__37081),
            .I(N__37062));
    InMux I__8244 (
            .O(N__37080),
            .I(N__37062));
    InMux I__8243 (
            .O(N__37079),
            .I(N__37062));
    InMux I__8242 (
            .O(N__37078),
            .I(N__37062));
    InMux I__8241 (
            .O(N__37077),
            .I(N__37059));
    Odrv4 I__8240 (
            .O(N__37074),
            .I(\c0.FRAME_MATCHER_i_2 ));
    Odrv4 I__8239 (
            .O(N__37071),
            .I(\c0.FRAME_MATCHER_i_2 ));
    LocalMux I__8238 (
            .O(N__37062),
            .I(\c0.FRAME_MATCHER_i_2 ));
    LocalMux I__8237 (
            .O(N__37059),
            .I(\c0.FRAME_MATCHER_i_2 ));
    CascadeMux I__8236 (
            .O(N__37050),
            .I(\c0.n15171_cascade_ ));
    CascadeMux I__8235 (
            .O(N__37047),
            .I(N__37040));
    InMux I__8234 (
            .O(N__37046),
            .I(N__37037));
    InMux I__8233 (
            .O(N__37045),
            .I(N__37034));
    InMux I__8232 (
            .O(N__37044),
            .I(N__37029));
    InMux I__8231 (
            .O(N__37043),
            .I(N__37029));
    InMux I__8230 (
            .O(N__37040),
            .I(N__37026));
    LocalMux I__8229 (
            .O(N__37037),
            .I(\c0.data_in_frame_1_6 ));
    LocalMux I__8228 (
            .O(N__37034),
            .I(\c0.data_in_frame_1_6 ));
    LocalMux I__8227 (
            .O(N__37029),
            .I(\c0.data_in_frame_1_6 ));
    LocalMux I__8226 (
            .O(N__37026),
            .I(\c0.data_in_frame_1_6 ));
    InMux I__8225 (
            .O(N__37017),
            .I(N__37014));
    LocalMux I__8224 (
            .O(N__37014),
            .I(N__37011));
    Span4Mux_h I__8223 (
            .O(N__37011),
            .I(N__37007));
    InMux I__8222 (
            .O(N__37010),
            .I(N__37004));
    Odrv4 I__8221 (
            .O(N__37007),
            .I(\c0.n2124 ));
    LocalMux I__8220 (
            .O(N__37004),
            .I(\c0.n2124 ));
    CascadeMux I__8219 (
            .O(N__36999),
            .I(N__36996));
    InMux I__8218 (
            .O(N__36996),
            .I(N__36993));
    LocalMux I__8217 (
            .O(N__36993),
            .I(N__36989));
    InMux I__8216 (
            .O(N__36992),
            .I(N__36986));
    Span4Mux_v I__8215 (
            .O(N__36989),
            .I(N__36983));
    LocalMux I__8214 (
            .O(N__36986),
            .I(data_in_frame_6_6));
    Odrv4 I__8213 (
            .O(N__36983),
            .I(data_in_frame_6_6));
    InMux I__8212 (
            .O(N__36978),
            .I(N__36975));
    LocalMux I__8211 (
            .O(N__36975),
            .I(\c0.n17214 ));
    InMux I__8210 (
            .O(N__36972),
            .I(N__36969));
    LocalMux I__8209 (
            .O(N__36969),
            .I(\c0.n28_adj_2374 ));
    CascadeMux I__8208 (
            .O(N__36966),
            .I(\c0.n27_adj_2381_cascade_ ));
    InMux I__8207 (
            .O(N__36963),
            .I(N__36960));
    LocalMux I__8206 (
            .O(N__36960),
            .I(\c0.n29 ));
    CascadeMux I__8205 (
            .O(N__36957),
            .I(\c0.n12491_cascade_ ));
    InMux I__8204 (
            .O(N__36954),
            .I(N__36950));
    InMux I__8203 (
            .O(N__36953),
            .I(N__36944));
    LocalMux I__8202 (
            .O(N__36950),
            .I(N__36941));
    InMux I__8201 (
            .O(N__36949),
            .I(N__36938));
    InMux I__8200 (
            .O(N__36948),
            .I(N__36935));
    InMux I__8199 (
            .O(N__36947),
            .I(N__36932));
    LocalMux I__8198 (
            .O(N__36944),
            .I(\c0.data_in_frame_0_1 ));
    Odrv4 I__8197 (
            .O(N__36941),
            .I(\c0.data_in_frame_0_1 ));
    LocalMux I__8196 (
            .O(N__36938),
            .I(\c0.data_in_frame_0_1 ));
    LocalMux I__8195 (
            .O(N__36935),
            .I(\c0.data_in_frame_0_1 ));
    LocalMux I__8194 (
            .O(N__36932),
            .I(\c0.data_in_frame_0_1 ));
    InMux I__8193 (
            .O(N__36921),
            .I(N__36918));
    LocalMux I__8192 (
            .O(N__36918),
            .I(N__36914));
    InMux I__8191 (
            .O(N__36917),
            .I(N__36911));
    Odrv4 I__8190 (
            .O(N__36914),
            .I(\c0.n10259 ));
    LocalMux I__8189 (
            .O(N__36911),
            .I(\c0.n10259 ));
    InMux I__8188 (
            .O(N__36906),
            .I(N__36903));
    LocalMux I__8187 (
            .O(N__36903),
            .I(N__36899));
    InMux I__8186 (
            .O(N__36902),
            .I(N__36895));
    Span4Mux_h I__8185 (
            .O(N__36899),
            .I(N__36892));
    InMux I__8184 (
            .O(N__36898),
            .I(N__36889));
    LocalMux I__8183 (
            .O(N__36895),
            .I(\c0.data_in_frame_2_7 ));
    Odrv4 I__8182 (
            .O(N__36892),
            .I(\c0.data_in_frame_2_7 ));
    LocalMux I__8181 (
            .O(N__36889),
            .I(\c0.data_in_frame_2_7 ));
    CascadeMux I__8180 (
            .O(N__36882),
            .I(N__36878));
    InMux I__8179 (
            .O(N__36881),
            .I(N__36873));
    InMux I__8178 (
            .O(N__36878),
            .I(N__36870));
    InMux I__8177 (
            .O(N__36877),
            .I(N__36867));
    InMux I__8176 (
            .O(N__36876),
            .I(N__36864));
    LocalMux I__8175 (
            .O(N__36873),
            .I(N__36858));
    LocalMux I__8174 (
            .O(N__36870),
            .I(N__36853));
    LocalMux I__8173 (
            .O(N__36867),
            .I(N__36853));
    LocalMux I__8172 (
            .O(N__36864),
            .I(N__36850));
    InMux I__8171 (
            .O(N__36863),
            .I(N__36847));
    CascadeMux I__8170 (
            .O(N__36862),
            .I(N__36844));
    CascadeMux I__8169 (
            .O(N__36861),
            .I(N__36841));
    Span4Mux_v I__8168 (
            .O(N__36858),
            .I(N__36835));
    Span4Mux_v I__8167 (
            .O(N__36853),
            .I(N__36835));
    Span4Mux_v I__8166 (
            .O(N__36850),
            .I(N__36830));
    LocalMux I__8165 (
            .O(N__36847),
            .I(N__36830));
    InMux I__8164 (
            .O(N__36844),
            .I(N__36827));
    InMux I__8163 (
            .O(N__36841),
            .I(N__36824));
    InMux I__8162 (
            .O(N__36840),
            .I(N__36821));
    Span4Mux_h I__8161 (
            .O(N__36835),
            .I(N__36818));
    Span4Mux_v I__8160 (
            .O(N__36830),
            .I(N__36815));
    LocalMux I__8159 (
            .O(N__36827),
            .I(rx_data_2));
    LocalMux I__8158 (
            .O(N__36824),
            .I(rx_data_2));
    LocalMux I__8157 (
            .O(N__36821),
            .I(rx_data_2));
    Odrv4 I__8156 (
            .O(N__36818),
            .I(rx_data_2));
    Odrv4 I__8155 (
            .O(N__36815),
            .I(rx_data_2));
    InMux I__8154 (
            .O(N__36804),
            .I(N__36795));
    InMux I__8153 (
            .O(N__36803),
            .I(N__36790));
    InMux I__8152 (
            .O(N__36802),
            .I(N__36790));
    InMux I__8151 (
            .O(N__36801),
            .I(N__36787));
    InMux I__8150 (
            .O(N__36800),
            .I(N__36782));
    InMux I__8149 (
            .O(N__36799),
            .I(N__36782));
    InMux I__8148 (
            .O(N__36798),
            .I(N__36779));
    LocalMux I__8147 (
            .O(N__36795),
            .I(N__36775));
    LocalMux I__8146 (
            .O(N__36790),
            .I(N__36770));
    LocalMux I__8145 (
            .O(N__36787),
            .I(N__36770));
    LocalMux I__8144 (
            .O(N__36782),
            .I(N__36765));
    LocalMux I__8143 (
            .O(N__36779),
            .I(N__36765));
    CascadeMux I__8142 (
            .O(N__36778),
            .I(N__36762));
    Span4Mux_h I__8141 (
            .O(N__36775),
            .I(N__36757));
    Span4Mux_h I__8140 (
            .O(N__36770),
            .I(N__36757));
    Span4Mux_v I__8139 (
            .O(N__36765),
            .I(N__36754));
    InMux I__8138 (
            .O(N__36762),
            .I(N__36751));
    Span4Mux_h I__8137 (
            .O(N__36757),
            .I(N__36748));
    Span4Mux_h I__8136 (
            .O(N__36754),
            .I(N__36745));
    LocalMux I__8135 (
            .O(N__36751),
            .I(rx_data_0));
    Odrv4 I__8134 (
            .O(N__36748),
            .I(rx_data_0));
    Odrv4 I__8133 (
            .O(N__36745),
            .I(rx_data_0));
    InMux I__8132 (
            .O(N__36738),
            .I(N__36735));
    LocalMux I__8131 (
            .O(N__36735),
            .I(N__36732));
    Sp12to4 I__8130 (
            .O(N__36732),
            .I(N__36729));
    Span12Mux_v I__8129 (
            .O(N__36729),
            .I(N__36726));
    Span12Mux_h I__8128 (
            .O(N__36726),
            .I(N__36723));
    Odrv12 I__8127 (
            .O(N__36723),
            .I(\c0.rx.r_Rx_Data_R ));
    InMux I__8126 (
            .O(N__36720),
            .I(N__36711));
    InMux I__8125 (
            .O(N__36719),
            .I(N__36711));
    InMux I__8124 (
            .O(N__36718),
            .I(N__36711));
    LocalMux I__8123 (
            .O(N__36711),
            .I(N__36707));
    InMux I__8122 (
            .O(N__36710),
            .I(N__36704));
    Span4Mux_v I__8121 (
            .O(N__36707),
            .I(N__36699));
    LocalMux I__8120 (
            .O(N__36704),
            .I(N__36699));
    Span4Mux_h I__8119 (
            .O(N__36699),
            .I(N__36696));
    Span4Mux_v I__8118 (
            .O(N__36696),
            .I(N__36693));
    Odrv4 I__8117 (
            .O(N__36693),
            .I(n10010));
    CascadeMux I__8116 (
            .O(N__36690),
            .I(N__36684));
    CascadeMux I__8115 (
            .O(N__36689),
            .I(N__36681));
    CascadeMux I__8114 (
            .O(N__36688),
            .I(N__36676));
    InMux I__8113 (
            .O(N__36687),
            .I(N__36670));
    InMux I__8112 (
            .O(N__36684),
            .I(N__36670));
    InMux I__8111 (
            .O(N__36681),
            .I(N__36665));
    InMux I__8110 (
            .O(N__36680),
            .I(N__36665));
    InMux I__8109 (
            .O(N__36679),
            .I(N__36662));
    InMux I__8108 (
            .O(N__36676),
            .I(N__36659));
    InMux I__8107 (
            .O(N__36675),
            .I(N__36656));
    LocalMux I__8106 (
            .O(N__36670),
            .I(N__36652));
    LocalMux I__8105 (
            .O(N__36665),
            .I(N__36649));
    LocalMux I__8104 (
            .O(N__36662),
            .I(N__36646));
    LocalMux I__8103 (
            .O(N__36659),
            .I(N__36641));
    LocalMux I__8102 (
            .O(N__36656),
            .I(N__36641));
    InMux I__8101 (
            .O(N__36655),
            .I(N__36638));
    Span4Mux_h I__8100 (
            .O(N__36652),
            .I(N__36635));
    Span4Mux_h I__8099 (
            .O(N__36649),
            .I(N__36632));
    Span4Mux_v I__8098 (
            .O(N__36646),
            .I(N__36627));
    Span4Mux_h I__8097 (
            .O(N__36641),
            .I(N__36627));
    LocalMux I__8096 (
            .O(N__36638),
            .I(rx_data_5));
    Odrv4 I__8095 (
            .O(N__36635),
            .I(rx_data_5));
    Odrv4 I__8094 (
            .O(N__36632),
            .I(rx_data_5));
    Odrv4 I__8093 (
            .O(N__36627),
            .I(rx_data_5));
    InMux I__8092 (
            .O(N__36618),
            .I(N__36615));
    LocalMux I__8091 (
            .O(N__36615),
            .I(N__36612));
    Odrv12 I__8090 (
            .O(N__36612),
            .I(\c0.n24_adj_2317 ));
    CascadeMux I__8089 (
            .O(N__36609),
            .I(N__36606));
    InMux I__8088 (
            .O(N__36606),
            .I(N__36603));
    LocalMux I__8087 (
            .O(N__36603),
            .I(N__36600));
    Odrv4 I__8086 (
            .O(N__36600),
            .I(\c0.n22_adj_2319 ));
    InMux I__8085 (
            .O(N__36597),
            .I(N__36594));
    LocalMux I__8084 (
            .O(N__36594),
            .I(\c0.n21_adj_2323 ));
    CascadeMux I__8083 (
            .O(N__36591),
            .I(N__36588));
    InMux I__8082 (
            .O(N__36588),
            .I(N__36585));
    LocalMux I__8081 (
            .O(N__36585),
            .I(\c0.n22_adj_2313 ));
    InMux I__8080 (
            .O(N__36582),
            .I(\c0.n16071 ));
    InMux I__8079 (
            .O(N__36579),
            .I(N__36576));
    LocalMux I__8078 (
            .O(N__36576),
            .I(\c0.n21_adj_2262 ));
    InMux I__8077 (
            .O(N__36573),
            .I(\c0.n16072 ));
    InMux I__8076 (
            .O(N__36570),
            .I(bfn_12_32_0_));
    InMux I__8075 (
            .O(N__36567),
            .I(\c0.n16074 ));
    InMux I__8074 (
            .O(N__36564),
            .I(\c0.n16075 ));
    InMux I__8073 (
            .O(N__36561),
            .I(\c0.n16076 ));
    InMux I__8072 (
            .O(N__36558),
            .I(\c0.n16077 ));
    InMux I__8071 (
            .O(N__36555),
            .I(\c0.n16078 ));
    CEMux I__8070 (
            .O(N__36552),
            .I(N__36548));
    CEMux I__8069 (
            .O(N__36551),
            .I(N__36545));
    LocalMux I__8068 (
            .O(N__36548),
            .I(N__36542));
    LocalMux I__8067 (
            .O(N__36545),
            .I(N__36539));
    Span4Mux_h I__8066 (
            .O(N__36542),
            .I(N__36536));
    Span4Mux_s2_v I__8065 (
            .O(N__36539),
            .I(N__36533));
    Odrv4 I__8064 (
            .O(N__36536),
            .I(\c0.n10594 ));
    Odrv4 I__8063 (
            .O(N__36533),
            .I(\c0.n10594 ));
    InMux I__8062 (
            .O(N__36528),
            .I(N__36525));
    LocalMux I__8061 (
            .O(N__36525),
            .I(\c0.n16353 ));
    InMux I__8060 (
            .O(N__36522),
            .I(N__36519));
    LocalMux I__8059 (
            .O(N__36519),
            .I(N__36516));
    Odrv4 I__8058 (
            .O(N__36516),
            .I(\c0.n26_adj_2368 ));
    CascadeMux I__8057 (
            .O(N__36513),
            .I(N__36510));
    InMux I__8056 (
            .O(N__36510),
            .I(N__36507));
    LocalMux I__8055 (
            .O(N__36507),
            .I(N__36504));
    Odrv12 I__8054 (
            .O(N__36504),
            .I(\c0.n16474 ));
    InMux I__8053 (
            .O(N__36501),
            .I(N__36498));
    LocalMux I__8052 (
            .O(N__36498),
            .I(\c0.n18_adj_2360 ));
    InMux I__8051 (
            .O(N__36495),
            .I(N__36492));
    LocalMux I__8050 (
            .O(N__36492),
            .I(\c0.n27 ));
    InMux I__8049 (
            .O(N__36489),
            .I(\c0.n16066 ));
    InMux I__8048 (
            .O(N__36486),
            .I(\c0.n16067 ));
    CascadeMux I__8047 (
            .O(N__36483),
            .I(N__36480));
    InMux I__8046 (
            .O(N__36480),
            .I(N__36477));
    LocalMux I__8045 (
            .O(N__36477),
            .I(\c0.n25_adj_2386 ));
    InMux I__8044 (
            .O(N__36474),
            .I(\c0.n16068 ));
    InMux I__8043 (
            .O(N__36471),
            .I(\c0.n16069 ));
    InMux I__8042 (
            .O(N__36468),
            .I(\c0.n16070 ));
    CascadeMux I__8041 (
            .O(N__36465),
            .I(n4_adj_2419_cascade_));
    CascadeMux I__8040 (
            .O(N__36462),
            .I(n5_adj_2407_cascade_));
    CascadeMux I__8039 (
            .O(N__36459),
            .I(n10_adj_2444_cascade_));
    InMux I__8038 (
            .O(N__36456),
            .I(N__36453));
    LocalMux I__8037 (
            .O(N__36453),
            .I(n8_adj_2447));
    InMux I__8036 (
            .O(N__36450),
            .I(N__36447));
    LocalMux I__8035 (
            .O(N__36447),
            .I(n4_adj_2419));
    InMux I__8034 (
            .O(N__36444),
            .I(N__36441));
    LocalMux I__8033 (
            .O(N__36441),
            .I(N__36438));
    Span4Mux_v I__8032 (
            .O(N__36438),
            .I(N__36435));
    Odrv4 I__8031 (
            .O(N__36435),
            .I(\c0.n17696 ));
    CascadeMux I__8030 (
            .O(N__36432),
            .I(n18073_cascade_));
    CascadeMux I__8029 (
            .O(N__36429),
            .I(\c0.tx.n10688_cascade_ ));
    CascadeMux I__8028 (
            .O(N__36426),
            .I(N__36422));
    InMux I__8027 (
            .O(N__36425),
            .I(N__36417));
    InMux I__8026 (
            .O(N__36422),
            .I(N__36417));
    LocalMux I__8025 (
            .O(N__36417),
            .I(r_Tx_Data_1));
    InMux I__8024 (
            .O(N__36414),
            .I(N__36411));
    LocalMux I__8023 (
            .O(N__36411),
            .I(N__36407));
    CascadeMux I__8022 (
            .O(N__36410),
            .I(N__36404));
    Span4Mux_v I__8021 (
            .O(N__36407),
            .I(N__36401));
    InMux I__8020 (
            .O(N__36404),
            .I(N__36398));
    Odrv4 I__8019 (
            .O(N__36401),
            .I(rand_setpoint_1));
    LocalMux I__8018 (
            .O(N__36398),
            .I(rand_setpoint_1));
    InMux I__8017 (
            .O(N__36393),
            .I(N__36389));
    InMux I__8016 (
            .O(N__36392),
            .I(N__36386));
    LocalMux I__8015 (
            .O(N__36389),
            .I(N__36383));
    LocalMux I__8014 (
            .O(N__36386),
            .I(r_Tx_Data_3));
    Odrv4 I__8013 (
            .O(N__36383),
            .I(r_Tx_Data_3));
    InMux I__8012 (
            .O(N__36378),
            .I(N__36375));
    LocalMux I__8011 (
            .O(N__36375),
            .I(n18070));
    InMux I__8010 (
            .O(N__36372),
            .I(N__36367));
    InMux I__8009 (
            .O(N__36371),
            .I(N__36362));
    InMux I__8008 (
            .O(N__36370),
            .I(N__36362));
    LocalMux I__8007 (
            .O(N__36367),
            .I(\c0.tx.n10688 ));
    LocalMux I__8006 (
            .O(N__36362),
            .I(\c0.tx.n10688 ));
    CascadeMux I__8005 (
            .O(N__36357),
            .I(n10_adj_2409_cascade_));
    CascadeMux I__8004 (
            .O(N__36354),
            .I(\c0.n8_adj_2183_cascade_ ));
    InMux I__8003 (
            .O(N__36351),
            .I(N__36348));
    LocalMux I__8002 (
            .O(N__36348),
            .I(\c0.n17671 ));
    InMux I__8001 (
            .O(N__36345),
            .I(N__36342));
    LocalMux I__8000 (
            .O(N__36342),
            .I(N__36339));
    Span4Mux_h I__7999 (
            .O(N__36339),
            .I(N__36335));
    CascadeMux I__7998 (
            .O(N__36338),
            .I(N__36332));
    Sp12to4 I__7997 (
            .O(N__36335),
            .I(N__36329));
    InMux I__7996 (
            .O(N__36332),
            .I(N__36326));
    Odrv12 I__7995 (
            .O(N__36329),
            .I(rand_setpoint_4));
    LocalMux I__7994 (
            .O(N__36326),
            .I(rand_setpoint_4));
    CascadeMux I__7993 (
            .O(N__36321),
            .I(data_out_10__7__N_110_cascade_));
    InMux I__7992 (
            .O(N__36318),
            .I(N__36315));
    LocalMux I__7991 (
            .O(N__36315),
            .I(N__36311));
    CascadeMux I__7990 (
            .O(N__36314),
            .I(N__36308));
    Span4Mux_h I__7989 (
            .O(N__36311),
            .I(N__36305));
    InMux I__7988 (
            .O(N__36308),
            .I(N__36302));
    Odrv4 I__7987 (
            .O(N__36305),
            .I(rand_setpoint_6));
    LocalMux I__7986 (
            .O(N__36302),
            .I(rand_setpoint_6));
    InMux I__7985 (
            .O(N__36297),
            .I(N__36294));
    LocalMux I__7984 (
            .O(N__36294),
            .I(N__36290));
    InMux I__7983 (
            .O(N__36293),
            .I(N__36287));
    Span4Mux_h I__7982 (
            .O(N__36290),
            .I(N__36284));
    LocalMux I__7981 (
            .O(N__36287),
            .I(\c0.data_out_1_2 ));
    Odrv4 I__7980 (
            .O(N__36284),
            .I(\c0.data_out_1_2 ));
    InMux I__7979 (
            .O(N__36279),
            .I(N__36276));
    LocalMux I__7978 (
            .O(N__36276),
            .I(N__36272));
    InMux I__7977 (
            .O(N__36275),
            .I(N__36269));
    Span4Mux_v I__7976 (
            .O(N__36272),
            .I(N__36266));
    LocalMux I__7975 (
            .O(N__36269),
            .I(N__36263));
    Span4Mux_h I__7974 (
            .O(N__36266),
            .I(N__36258));
    Span4Mux_v I__7973 (
            .O(N__36263),
            .I(N__36258));
    Span4Mux_v I__7972 (
            .O(N__36258),
            .I(N__36254));
    InMux I__7971 (
            .O(N__36257),
            .I(N__36251));
    Odrv4 I__7970 (
            .O(N__36254),
            .I(blink_counter_24));
    LocalMux I__7969 (
            .O(N__36251),
            .I(blink_counter_24));
    InMux I__7968 (
            .O(N__36246),
            .I(N__36242));
    InMux I__7967 (
            .O(N__36245),
            .I(N__36239));
    LocalMux I__7966 (
            .O(N__36242),
            .I(N__36236));
    LocalMux I__7965 (
            .O(N__36239),
            .I(N__36233));
    Span4Mux_v I__7964 (
            .O(N__36236),
            .I(N__36230));
    Span4Mux_v I__7963 (
            .O(N__36233),
            .I(N__36227));
    Span4Mux_v I__7962 (
            .O(N__36230),
            .I(N__36223));
    Span4Mux_v I__7961 (
            .O(N__36227),
            .I(N__36220));
    InMux I__7960 (
            .O(N__36226),
            .I(N__36217));
    Odrv4 I__7959 (
            .O(N__36223),
            .I(blink_counter_23));
    Odrv4 I__7958 (
            .O(N__36220),
            .I(blink_counter_23));
    LocalMux I__7957 (
            .O(N__36217),
            .I(blink_counter_23));
    CascadeMux I__7956 (
            .O(N__36210),
            .I(N__36207));
    InMux I__7955 (
            .O(N__36207),
            .I(N__36204));
    LocalMux I__7954 (
            .O(N__36204),
            .I(N__36200));
    InMux I__7953 (
            .O(N__36203),
            .I(N__36197));
    Span4Mux_v I__7952 (
            .O(N__36200),
            .I(N__36194));
    LocalMux I__7951 (
            .O(N__36197),
            .I(N__36191));
    Span4Mux_v I__7950 (
            .O(N__36194),
            .I(N__36187));
    Span12Mux_v I__7949 (
            .O(N__36191),
            .I(N__36184));
    InMux I__7948 (
            .O(N__36190),
            .I(N__36181));
    Odrv4 I__7947 (
            .O(N__36187),
            .I(blink_counter_22));
    Odrv12 I__7946 (
            .O(N__36184),
            .I(blink_counter_22));
    LocalMux I__7945 (
            .O(N__36181),
            .I(blink_counter_22));
    CascadeMux I__7944 (
            .O(N__36174),
            .I(N__36171));
    InMux I__7943 (
            .O(N__36171),
            .I(N__36167));
    InMux I__7942 (
            .O(N__36170),
            .I(N__36164));
    LocalMux I__7941 (
            .O(N__36167),
            .I(N__36161));
    LocalMux I__7940 (
            .O(N__36164),
            .I(N__36158));
    Span4Mux_v I__7939 (
            .O(N__36161),
            .I(N__36155));
    Span12Mux_v I__7938 (
            .O(N__36158),
            .I(N__36151));
    Span4Mux_v I__7937 (
            .O(N__36155),
            .I(N__36148));
    InMux I__7936 (
            .O(N__36154),
            .I(N__36145));
    Odrv12 I__7935 (
            .O(N__36151),
            .I(blink_counter_21));
    Odrv4 I__7934 (
            .O(N__36148),
            .I(blink_counter_21));
    LocalMux I__7933 (
            .O(N__36145),
            .I(blink_counter_21));
    InMux I__7932 (
            .O(N__36138),
            .I(N__36135));
    LocalMux I__7931 (
            .O(N__36135),
            .I(N__36132));
    Odrv4 I__7930 (
            .O(N__36132),
            .I(n10140));
    InMux I__7929 (
            .O(N__36129),
            .I(N__36126));
    LocalMux I__7928 (
            .O(N__36126),
            .I(n8));
    CascadeMux I__7927 (
            .O(N__36123),
            .I(n4_adj_2417_cascade_));
    InMux I__7926 (
            .O(N__36120),
            .I(N__36115));
    InMux I__7925 (
            .O(N__36119),
            .I(N__36110));
    InMux I__7924 (
            .O(N__36118),
            .I(N__36110));
    LocalMux I__7923 (
            .O(N__36115),
            .I(N__36104));
    LocalMux I__7922 (
            .O(N__36110),
            .I(N__36104));
    InMux I__7921 (
            .O(N__36109),
            .I(N__36101));
    Span4Mux_v I__7920 (
            .O(N__36104),
            .I(N__36096));
    LocalMux I__7919 (
            .O(N__36101),
            .I(N__36096));
    Odrv4 I__7918 (
            .O(N__36096),
            .I(FRAME_MATCHER_state_31_N_1406_2));
    CascadeMux I__7917 (
            .O(N__36093),
            .I(N__36087));
    InMux I__7916 (
            .O(N__36092),
            .I(N__36083));
    InMux I__7915 (
            .O(N__36091),
            .I(N__36078));
    InMux I__7914 (
            .O(N__36090),
            .I(N__36078));
    InMux I__7913 (
            .O(N__36087),
            .I(N__36073));
    InMux I__7912 (
            .O(N__36086),
            .I(N__36073));
    LocalMux I__7911 (
            .O(N__36083),
            .I(N__36066));
    LocalMux I__7910 (
            .O(N__36078),
            .I(N__36063));
    LocalMux I__7909 (
            .O(N__36073),
            .I(N__36058));
    InMux I__7908 (
            .O(N__36072),
            .I(N__36055));
    InMux I__7907 (
            .O(N__36071),
            .I(N__36050));
    InMux I__7906 (
            .O(N__36070),
            .I(N__36050));
    InMux I__7905 (
            .O(N__36069),
            .I(N__36047));
    Span12Mux_v I__7904 (
            .O(N__36066),
            .I(N__36044));
    Span4Mux_v I__7903 (
            .O(N__36063),
            .I(N__36041));
    InMux I__7902 (
            .O(N__36062),
            .I(N__36036));
    InMux I__7901 (
            .O(N__36061),
            .I(N__36036));
    Span4Mux_h I__7900 (
            .O(N__36058),
            .I(N__36031));
    LocalMux I__7899 (
            .O(N__36055),
            .I(N__36031));
    LocalMux I__7898 (
            .O(N__36050),
            .I(N__36028));
    LocalMux I__7897 (
            .O(N__36047),
            .I(FRAME_MATCHER_state_2));
    Odrv12 I__7896 (
            .O(N__36044),
            .I(FRAME_MATCHER_state_2));
    Odrv4 I__7895 (
            .O(N__36041),
            .I(FRAME_MATCHER_state_2));
    LocalMux I__7894 (
            .O(N__36036),
            .I(FRAME_MATCHER_state_2));
    Odrv4 I__7893 (
            .O(N__36031),
            .I(FRAME_MATCHER_state_2));
    Odrv4 I__7892 (
            .O(N__36028),
            .I(FRAME_MATCHER_state_2));
    InMux I__7891 (
            .O(N__36015),
            .I(N__36012));
    LocalMux I__7890 (
            .O(N__36012),
            .I(N__36009));
    Span4Mux_v I__7889 (
            .O(N__36009),
            .I(N__36006));
    Span4Mux_v I__7888 (
            .O(N__36006),
            .I(N__36002));
    InMux I__7887 (
            .O(N__36005),
            .I(N__35999));
    Odrv4 I__7886 (
            .O(N__36002),
            .I(blink_counter_25));
    LocalMux I__7885 (
            .O(N__35999),
            .I(blink_counter_25));
    InMux I__7884 (
            .O(N__35994),
            .I(N__35991));
    LocalMux I__7883 (
            .O(N__35991),
            .I(n17428));
    InMux I__7882 (
            .O(N__35988),
            .I(N__35985));
    LocalMux I__7881 (
            .O(N__35985),
            .I(N__35982));
    Span4Mux_v I__7880 (
            .O(N__35982),
            .I(N__35979));
    Odrv4 I__7879 (
            .O(N__35979),
            .I(n17427));
    IoInMux I__7878 (
            .O(N__35976),
            .I(N__35973));
    LocalMux I__7877 (
            .O(N__35973),
            .I(N__35970));
    Span4Mux_s3_v I__7876 (
            .O(N__35970),
            .I(N__35967));
    Span4Mux_v I__7875 (
            .O(N__35967),
            .I(N__35964));
    Sp12to4 I__7874 (
            .O(N__35964),
            .I(N__35961));
    Odrv12 I__7873 (
            .O(N__35961),
            .I(LED_c));
    CascadeMux I__7872 (
            .O(N__35958),
            .I(N__35954));
    CascadeMux I__7871 (
            .O(N__35957),
            .I(N__35951));
    InMux I__7870 (
            .O(N__35954),
            .I(N__35947));
    InMux I__7869 (
            .O(N__35951),
            .I(N__35942));
    InMux I__7868 (
            .O(N__35950),
            .I(N__35942));
    LocalMux I__7867 (
            .O(N__35947),
            .I(N__35937));
    LocalMux I__7866 (
            .O(N__35942),
            .I(N__35934));
    InMux I__7865 (
            .O(N__35941),
            .I(N__35929));
    InMux I__7864 (
            .O(N__35940),
            .I(N__35929));
    Span4Mux_h I__7863 (
            .O(N__35937),
            .I(N__35926));
    Span4Mux_h I__7862 (
            .O(N__35934),
            .I(N__35923));
    LocalMux I__7861 (
            .O(N__35929),
            .I(N__35920));
    Span4Mux_h I__7860 (
            .O(N__35926),
            .I(N__35917));
    Span4Mux_h I__7859 (
            .O(N__35923),
            .I(N__35914));
    Span4Mux_v I__7858 (
            .O(N__35920),
            .I(N__35911));
    Odrv4 I__7857 (
            .O(N__35917),
            .I(n3779));
    Odrv4 I__7856 (
            .O(N__35914),
            .I(n3779));
    Odrv4 I__7855 (
            .O(N__35911),
            .I(n3779));
    InMux I__7854 (
            .O(N__35904),
            .I(N__35899));
    InMux I__7853 (
            .O(N__35903),
            .I(N__35896));
    InMux I__7852 (
            .O(N__35902),
            .I(N__35893));
    LocalMux I__7851 (
            .O(N__35899),
            .I(N__35888));
    LocalMux I__7850 (
            .O(N__35896),
            .I(N__35883));
    LocalMux I__7849 (
            .O(N__35893),
            .I(N__35883));
    InMux I__7848 (
            .O(N__35892),
            .I(N__35878));
    InMux I__7847 (
            .O(N__35891),
            .I(N__35878));
    Odrv4 I__7846 (
            .O(N__35888),
            .I(FRAME_MATCHER_i_31__N_1273));
    Odrv4 I__7845 (
            .O(N__35883),
            .I(FRAME_MATCHER_i_31__N_1273));
    LocalMux I__7844 (
            .O(N__35878),
            .I(FRAME_MATCHER_i_31__N_1273));
    CascadeMux I__7843 (
            .O(N__35871),
            .I(N__35868));
    InMux I__7842 (
            .O(N__35868),
            .I(N__35865));
    LocalMux I__7841 (
            .O(N__35865),
            .I(n6_adj_2488));
    InMux I__7840 (
            .O(N__35862),
            .I(N__35859));
    LocalMux I__7839 (
            .O(N__35859),
            .I(N__35855));
    InMux I__7838 (
            .O(N__35858),
            .I(N__35852));
    Span4Mux_v I__7837 (
            .O(N__35855),
            .I(N__35849));
    LocalMux I__7836 (
            .O(N__35852),
            .I(data_out_3_0));
    Odrv4 I__7835 (
            .O(N__35849),
            .I(data_out_3_0));
    InMux I__7834 (
            .O(N__35844),
            .I(N__35841));
    LocalMux I__7833 (
            .O(N__35841),
            .I(N__35838));
    Span4Mux_h I__7832 (
            .O(N__35838),
            .I(N__35835));
    Odrv4 I__7831 (
            .O(N__35835),
            .I(n18175));
    InMux I__7830 (
            .O(N__35832),
            .I(N__35829));
    LocalMux I__7829 (
            .O(N__35829),
            .I(N__35825));
    InMux I__7828 (
            .O(N__35828),
            .I(N__35822));
    Span12Mux_s11_h I__7827 (
            .O(N__35825),
            .I(N__35814));
    LocalMux I__7826 (
            .O(N__35822),
            .I(N__35811));
    InMux I__7825 (
            .O(N__35821),
            .I(N__35806));
    InMux I__7824 (
            .O(N__35820),
            .I(N__35806));
    InMux I__7823 (
            .O(N__35819),
            .I(N__35799));
    InMux I__7822 (
            .O(N__35818),
            .I(N__35799));
    InMux I__7821 (
            .O(N__35817),
            .I(N__35799));
    Odrv12 I__7820 (
            .O(N__35814),
            .I(n5));
    Odrv4 I__7819 (
            .O(N__35811),
            .I(n5));
    LocalMux I__7818 (
            .O(N__35806),
            .I(n5));
    LocalMux I__7817 (
            .O(N__35799),
            .I(n5));
    InMux I__7816 (
            .O(N__35790),
            .I(N__35787));
    LocalMux I__7815 (
            .O(N__35787),
            .I(N__35783));
    InMux I__7814 (
            .O(N__35786),
            .I(N__35780));
    Odrv4 I__7813 (
            .O(N__35783),
            .I(n1_adj_2486));
    LocalMux I__7812 (
            .O(N__35780),
            .I(n1_adj_2486));
    InMux I__7811 (
            .O(N__35775),
            .I(N__35772));
    LocalMux I__7810 (
            .O(N__35772),
            .I(N__35769));
    Odrv4 I__7809 (
            .O(N__35769),
            .I(n9378));
    CascadeMux I__7808 (
            .O(N__35766),
            .I(N__35762));
    CascadeMux I__7807 (
            .O(N__35765),
            .I(N__35759));
    InMux I__7806 (
            .O(N__35762),
            .I(N__35754));
    InMux I__7805 (
            .O(N__35759),
            .I(N__35751));
    CascadeMux I__7804 (
            .O(N__35758),
            .I(N__35747));
    InMux I__7803 (
            .O(N__35757),
            .I(N__35740));
    LocalMux I__7802 (
            .O(N__35754),
            .I(N__35737));
    LocalMux I__7801 (
            .O(N__35751),
            .I(N__35734));
    InMux I__7800 (
            .O(N__35750),
            .I(N__35729));
    InMux I__7799 (
            .O(N__35747),
            .I(N__35729));
    CascadeMux I__7798 (
            .O(N__35746),
            .I(N__35726));
    CascadeMux I__7797 (
            .O(N__35745),
            .I(N__35720));
    CascadeMux I__7796 (
            .O(N__35744),
            .I(N__35716));
    InMux I__7795 (
            .O(N__35743),
            .I(N__35713));
    LocalMux I__7794 (
            .O(N__35740),
            .I(N__35708));
    Span4Mux_h I__7793 (
            .O(N__35737),
            .I(N__35705));
    Span4Mux_h I__7792 (
            .O(N__35734),
            .I(N__35699));
    LocalMux I__7791 (
            .O(N__35729),
            .I(N__35696));
    InMux I__7790 (
            .O(N__35726),
            .I(N__35693));
    InMux I__7789 (
            .O(N__35725),
            .I(N__35690));
    InMux I__7788 (
            .O(N__35724),
            .I(N__35683));
    InMux I__7787 (
            .O(N__35723),
            .I(N__35683));
    InMux I__7786 (
            .O(N__35720),
            .I(N__35683));
    InMux I__7785 (
            .O(N__35719),
            .I(N__35679));
    InMux I__7784 (
            .O(N__35716),
            .I(N__35676));
    LocalMux I__7783 (
            .O(N__35713),
            .I(N__35673));
    InMux I__7782 (
            .O(N__35712),
            .I(N__35668));
    InMux I__7781 (
            .O(N__35711),
            .I(N__35668));
    Span4Mux_v I__7780 (
            .O(N__35708),
            .I(N__35663));
    Span4Mux_v I__7779 (
            .O(N__35705),
            .I(N__35663));
    InMux I__7778 (
            .O(N__35704),
            .I(N__35660));
    InMux I__7777 (
            .O(N__35703),
            .I(N__35655));
    InMux I__7776 (
            .O(N__35702),
            .I(N__35655));
    Span4Mux_v I__7775 (
            .O(N__35699),
            .I(N__35644));
    Span4Mux_h I__7774 (
            .O(N__35696),
            .I(N__35644));
    LocalMux I__7773 (
            .O(N__35693),
            .I(N__35644));
    LocalMux I__7772 (
            .O(N__35690),
            .I(N__35644));
    LocalMux I__7771 (
            .O(N__35683),
            .I(N__35644));
    InMux I__7770 (
            .O(N__35682),
            .I(N__35641));
    LocalMux I__7769 (
            .O(N__35679),
            .I(FRAME_MATCHER_state_1));
    LocalMux I__7768 (
            .O(N__35676),
            .I(FRAME_MATCHER_state_1));
    Odrv12 I__7767 (
            .O(N__35673),
            .I(FRAME_MATCHER_state_1));
    LocalMux I__7766 (
            .O(N__35668),
            .I(FRAME_MATCHER_state_1));
    Odrv4 I__7765 (
            .O(N__35663),
            .I(FRAME_MATCHER_state_1));
    LocalMux I__7764 (
            .O(N__35660),
            .I(FRAME_MATCHER_state_1));
    LocalMux I__7763 (
            .O(N__35655),
            .I(FRAME_MATCHER_state_1));
    Odrv4 I__7762 (
            .O(N__35644),
            .I(FRAME_MATCHER_state_1));
    LocalMux I__7761 (
            .O(N__35641),
            .I(FRAME_MATCHER_state_1));
    CascadeMux I__7760 (
            .O(N__35622),
            .I(N__35619));
    InMux I__7759 (
            .O(N__35619),
            .I(N__35616));
    LocalMux I__7758 (
            .O(N__35616),
            .I(N__35613));
    Odrv12 I__7757 (
            .O(N__35613),
            .I(\c0.n16261 ));
    InMux I__7756 (
            .O(N__35610),
            .I(N__35607));
    LocalMux I__7755 (
            .O(N__35607),
            .I(N__35602));
    InMux I__7754 (
            .O(N__35606),
            .I(N__35599));
    CascadeMux I__7753 (
            .O(N__35605),
            .I(N__35596));
    Span4Mux_h I__7752 (
            .O(N__35602),
            .I(N__35590));
    LocalMux I__7751 (
            .O(N__35599),
            .I(N__35590));
    InMux I__7750 (
            .O(N__35596),
            .I(N__35587));
    InMux I__7749 (
            .O(N__35595),
            .I(N__35584));
    Span4Mux_h I__7748 (
            .O(N__35590),
            .I(N__35579));
    LocalMux I__7747 (
            .O(N__35587),
            .I(N__35574));
    LocalMux I__7746 (
            .O(N__35584),
            .I(N__35574));
    InMux I__7745 (
            .O(N__35583),
            .I(N__35569));
    InMux I__7744 (
            .O(N__35582),
            .I(N__35569));
    Span4Mux_v I__7743 (
            .O(N__35579),
            .I(N__35566));
    Span12Mux_s11_h I__7742 (
            .O(N__35574),
            .I(N__35563));
    LocalMux I__7741 (
            .O(N__35569),
            .I(N__35560));
    Odrv4 I__7740 (
            .O(N__35566),
            .I(\c0.r_SM_Main_2_N_2034_0_adj_2167 ));
    Odrv12 I__7739 (
            .O(N__35563),
            .I(\c0.r_SM_Main_2_N_2034_0_adj_2167 ));
    Odrv12 I__7738 (
            .O(N__35560),
            .I(\c0.r_SM_Main_2_N_2034_0_adj_2167 ));
    SRMux I__7737 (
            .O(N__35553),
            .I(N__35546));
    InMux I__7736 (
            .O(N__35552),
            .I(N__35541));
    InMux I__7735 (
            .O(N__35551),
            .I(N__35541));
    InMux I__7734 (
            .O(N__35550),
            .I(N__35536));
    InMux I__7733 (
            .O(N__35549),
            .I(N__35536));
    LocalMux I__7732 (
            .O(N__35546),
            .I(N__35529));
    LocalMux I__7731 (
            .O(N__35541),
            .I(N__35526));
    LocalMux I__7730 (
            .O(N__35536),
            .I(N__35523));
    InMux I__7729 (
            .O(N__35535),
            .I(N__35518));
    InMux I__7728 (
            .O(N__35534),
            .I(N__35518));
    InMux I__7727 (
            .O(N__35533),
            .I(N__35515));
    InMux I__7726 (
            .O(N__35532),
            .I(N__35512));
    Odrv12 I__7725 (
            .O(N__35529),
            .I(\c0.n10018 ));
    Odrv4 I__7724 (
            .O(N__35526),
            .I(\c0.n10018 ));
    Odrv4 I__7723 (
            .O(N__35523),
            .I(\c0.n10018 ));
    LocalMux I__7722 (
            .O(N__35518),
            .I(\c0.n10018 ));
    LocalMux I__7721 (
            .O(N__35515),
            .I(\c0.n10018 ));
    LocalMux I__7720 (
            .O(N__35512),
            .I(\c0.n10018 ));
    InMux I__7719 (
            .O(N__35499),
            .I(N__35496));
    LocalMux I__7718 (
            .O(N__35496),
            .I(n10088));
    CascadeMux I__7717 (
            .O(N__35493),
            .I(N__35489));
    InMux I__7716 (
            .O(N__35492),
            .I(N__35486));
    InMux I__7715 (
            .O(N__35489),
            .I(N__35483));
    LocalMux I__7714 (
            .O(N__35486),
            .I(N__35480));
    LocalMux I__7713 (
            .O(N__35483),
            .I(N__35477));
    Span4Mux_v I__7712 (
            .O(N__35480),
            .I(N__35474));
    Span4Mux_h I__7711 (
            .O(N__35477),
            .I(N__35471));
    Span4Mux_h I__7710 (
            .O(N__35474),
            .I(N__35468));
    Odrv4 I__7709 (
            .O(N__35471),
            .I(n17086));
    Odrv4 I__7708 (
            .O(N__35468),
            .I(n17086));
    InMux I__7707 (
            .O(N__35463),
            .I(N__35457));
    InMux I__7706 (
            .O(N__35462),
            .I(N__35457));
    LocalMux I__7705 (
            .O(N__35457),
            .I(n17063));
    InMux I__7704 (
            .O(N__35454),
            .I(N__35448));
    InMux I__7703 (
            .O(N__35453),
            .I(N__35448));
    LocalMux I__7702 (
            .O(N__35448),
            .I(n17089));
    InMux I__7701 (
            .O(N__35445),
            .I(N__35442));
    LocalMux I__7700 (
            .O(N__35442),
            .I(n17090));
    InMux I__7699 (
            .O(N__35439),
            .I(N__35433));
    InMux I__7698 (
            .O(N__35438),
            .I(N__35433));
    LocalMux I__7697 (
            .O(N__35433),
            .I(n3_adj_2485));
    InMux I__7696 (
            .O(N__35430),
            .I(N__35427));
    LocalMux I__7695 (
            .O(N__35427),
            .I(N__35424));
    Odrv4 I__7694 (
            .O(N__35424),
            .I(n6));
    InMux I__7693 (
            .O(N__35421),
            .I(N__35415));
    InMux I__7692 (
            .O(N__35420),
            .I(N__35415));
    LocalMux I__7691 (
            .O(N__35415),
            .I(n17349));
    CascadeMux I__7690 (
            .O(N__35412),
            .I(n3_adj_2485_cascade_));
    InMux I__7689 (
            .O(N__35409),
            .I(N__35406));
    LocalMux I__7688 (
            .O(N__35406),
            .I(N__35402));
    CascadeMux I__7687 (
            .O(N__35405),
            .I(N__35398));
    Span4Mux_h I__7686 (
            .O(N__35402),
            .I(N__35395));
    InMux I__7685 (
            .O(N__35401),
            .I(N__35390));
    InMux I__7684 (
            .O(N__35398),
            .I(N__35390));
    Odrv4 I__7683 (
            .O(N__35395),
            .I(data_in_2_1));
    LocalMux I__7682 (
            .O(N__35390),
            .I(data_in_2_1));
    InMux I__7681 (
            .O(N__35385),
            .I(N__35381));
    InMux I__7680 (
            .O(N__35384),
            .I(N__35378));
    LocalMux I__7679 (
            .O(N__35381),
            .I(N__35374));
    LocalMux I__7678 (
            .O(N__35378),
            .I(N__35371));
    InMux I__7677 (
            .O(N__35377),
            .I(N__35367));
    Span4Mux_v I__7676 (
            .O(N__35374),
            .I(N__35364));
    Span4Mux_h I__7675 (
            .O(N__35371),
            .I(N__35361));
    InMux I__7674 (
            .O(N__35370),
            .I(N__35358));
    LocalMux I__7673 (
            .O(N__35367),
            .I(N__35353));
    Span4Mux_v I__7672 (
            .O(N__35364),
            .I(N__35353));
    Odrv4 I__7671 (
            .O(N__35361),
            .I(data_in_1_1));
    LocalMux I__7670 (
            .O(N__35358),
            .I(data_in_1_1));
    Odrv4 I__7669 (
            .O(N__35353),
            .I(data_in_1_1));
    CascadeMux I__7668 (
            .O(N__35346),
            .I(N__35342));
    CascadeMux I__7667 (
            .O(N__35345),
            .I(N__35339));
    InMux I__7666 (
            .O(N__35342),
            .I(N__35336));
    InMux I__7665 (
            .O(N__35339),
            .I(N__35333));
    LocalMux I__7664 (
            .O(N__35336),
            .I(N__35330));
    LocalMux I__7663 (
            .O(N__35333),
            .I(\c0.data_in_frame_3_5 ));
    Odrv12 I__7662 (
            .O(N__35330),
            .I(\c0.data_in_frame_3_5 ));
    InMux I__7661 (
            .O(N__35325),
            .I(N__35321));
    InMux I__7660 (
            .O(N__35324),
            .I(N__35318));
    LocalMux I__7659 (
            .O(N__35321),
            .I(N__35314));
    LocalMux I__7658 (
            .O(N__35318),
            .I(N__35311));
    InMux I__7657 (
            .O(N__35317),
            .I(N__35308));
    Sp12to4 I__7656 (
            .O(N__35314),
            .I(N__35303));
    Sp12to4 I__7655 (
            .O(N__35311),
            .I(N__35303));
    LocalMux I__7654 (
            .O(N__35308),
            .I(\c0.data_in_frame_2_3 ));
    Odrv12 I__7653 (
            .O(N__35303),
            .I(\c0.data_in_frame_2_3 ));
    CascadeMux I__7652 (
            .O(N__35298),
            .I(N__35294));
    CascadeMux I__7651 (
            .O(N__35297),
            .I(N__35289));
    InMux I__7650 (
            .O(N__35294),
            .I(N__35284));
    InMux I__7649 (
            .O(N__35293),
            .I(N__35281));
    CascadeMux I__7648 (
            .O(N__35292),
            .I(N__35278));
    InMux I__7647 (
            .O(N__35289),
            .I(N__35269));
    InMux I__7646 (
            .O(N__35288),
            .I(N__35269));
    InMux I__7645 (
            .O(N__35287),
            .I(N__35269));
    LocalMux I__7644 (
            .O(N__35284),
            .I(N__35264));
    LocalMux I__7643 (
            .O(N__35281),
            .I(N__35264));
    InMux I__7642 (
            .O(N__35278),
            .I(N__35261));
    InMux I__7641 (
            .O(N__35277),
            .I(N__35258));
    InMux I__7640 (
            .O(N__35276),
            .I(N__35255));
    LocalMux I__7639 (
            .O(N__35269),
            .I(N__35250));
    Span4Mux_v I__7638 (
            .O(N__35264),
            .I(N__35250));
    LocalMux I__7637 (
            .O(N__35261),
            .I(rx_data_3));
    LocalMux I__7636 (
            .O(N__35258),
            .I(rx_data_3));
    LocalMux I__7635 (
            .O(N__35255),
            .I(rx_data_3));
    Odrv4 I__7634 (
            .O(N__35250),
            .I(rx_data_3));
    InMux I__7633 (
            .O(N__35241),
            .I(N__35238));
    LocalMux I__7632 (
            .O(N__35238),
            .I(N__35234));
    InMux I__7631 (
            .O(N__35237),
            .I(N__35230));
    Span4Mux_h I__7630 (
            .O(N__35234),
            .I(N__35227));
    InMux I__7629 (
            .O(N__35233),
            .I(N__35224));
    LocalMux I__7628 (
            .O(N__35230),
            .I(N__35221));
    Odrv4 I__7627 (
            .O(N__35227),
            .I(data_in_3_3));
    LocalMux I__7626 (
            .O(N__35224),
            .I(data_in_3_3));
    Odrv12 I__7625 (
            .O(N__35221),
            .I(data_in_3_3));
    InMux I__7624 (
            .O(N__35214),
            .I(N__35211));
    LocalMux I__7623 (
            .O(N__35211),
            .I(N__35207));
    InMux I__7622 (
            .O(N__35210),
            .I(N__35204));
    Span4Mux_h I__7621 (
            .O(N__35207),
            .I(N__35201));
    LocalMux I__7620 (
            .O(N__35204),
            .I(N__35197));
    Span4Mux_h I__7619 (
            .O(N__35201),
            .I(N__35194));
    InMux I__7618 (
            .O(N__35200),
            .I(N__35191));
    Span12Mux_h I__7617 (
            .O(N__35197),
            .I(N__35188));
    Span4Mux_h I__7616 (
            .O(N__35194),
            .I(N__35185));
    LocalMux I__7615 (
            .O(N__35191),
            .I(\c0.FRAME_MATCHER_state_28 ));
    Odrv12 I__7614 (
            .O(N__35188),
            .I(\c0.FRAME_MATCHER_state_28 ));
    Odrv4 I__7613 (
            .O(N__35185),
            .I(\c0.FRAME_MATCHER_state_28 ));
    InMux I__7612 (
            .O(N__35178),
            .I(N__35175));
    LocalMux I__7611 (
            .O(N__35175),
            .I(N__35172));
    Span4Mux_h I__7610 (
            .O(N__35172),
            .I(N__35169));
    Odrv4 I__7609 (
            .O(N__35169),
            .I(\c0.n50 ));
    CascadeMux I__7608 (
            .O(N__35166),
            .I(\c0.n47_cascade_ ));
    InMux I__7607 (
            .O(N__35163),
            .I(N__35160));
    LocalMux I__7606 (
            .O(N__35160),
            .I(\c0.n49 ));
    InMux I__7605 (
            .O(N__35157),
            .I(N__35154));
    LocalMux I__7604 (
            .O(N__35154),
            .I(N__35151));
    Span12Mux_h I__7603 (
            .O(N__35151),
            .I(N__35148));
    Odrv12 I__7602 (
            .O(N__35148),
            .I(\c0.n51 ));
    CascadeMux I__7601 (
            .O(N__35145),
            .I(\c0.n56_cascade_ ));
    InMux I__7600 (
            .O(N__35142),
            .I(N__35139));
    LocalMux I__7599 (
            .O(N__35139),
            .I(N__35136));
    Span4Mux_h I__7598 (
            .O(N__35136),
            .I(N__35133));
    Odrv4 I__7597 (
            .O(N__35133),
            .I(\c0.n45 ));
    CascadeMux I__7596 (
            .O(N__35130),
            .I(\c0.n10018_cascade_ ));
    CascadeMux I__7595 (
            .O(N__35127),
            .I(N__35124));
    InMux I__7594 (
            .O(N__35124),
            .I(N__35121));
    LocalMux I__7593 (
            .O(N__35121),
            .I(N__35116));
    InMux I__7592 (
            .O(N__35120),
            .I(N__35113));
    CascadeMux I__7591 (
            .O(N__35119),
            .I(N__35110));
    Span4Mux_v I__7590 (
            .O(N__35116),
            .I(N__35105));
    LocalMux I__7589 (
            .O(N__35113),
            .I(N__35105));
    InMux I__7588 (
            .O(N__35110),
            .I(N__35102));
    Span4Mux_h I__7587 (
            .O(N__35105),
            .I(N__35099));
    LocalMux I__7586 (
            .O(N__35102),
            .I(\c0.data_in_frame_2_0 ));
    Odrv4 I__7585 (
            .O(N__35099),
            .I(\c0.data_in_frame_2_0 ));
    InMux I__7584 (
            .O(N__35094),
            .I(N__35089));
    InMux I__7583 (
            .O(N__35093),
            .I(N__35084));
    InMux I__7582 (
            .O(N__35092),
            .I(N__35084));
    LocalMux I__7581 (
            .O(N__35089),
            .I(N__35081));
    LocalMux I__7580 (
            .O(N__35084),
            .I(N__35078));
    Span4Mux_h I__7579 (
            .O(N__35081),
            .I(N__35075));
    Span4Mux_h I__7578 (
            .O(N__35078),
            .I(N__35071));
    Span4Mux_h I__7577 (
            .O(N__35075),
            .I(N__35068));
    InMux I__7576 (
            .O(N__35074),
            .I(N__35065));
    Span4Mux_v I__7575 (
            .O(N__35071),
            .I(N__35062));
    Odrv4 I__7574 (
            .O(N__35068),
            .I(data_in_3_6));
    LocalMux I__7573 (
            .O(N__35065),
            .I(data_in_3_6));
    Odrv4 I__7572 (
            .O(N__35062),
            .I(data_in_3_6));
    InMux I__7571 (
            .O(N__35055),
            .I(N__35052));
    LocalMux I__7570 (
            .O(N__35052),
            .I(N__35047));
    InMux I__7569 (
            .O(N__35051),
            .I(N__35044));
    InMux I__7568 (
            .O(N__35050),
            .I(N__35041));
    Odrv12 I__7567 (
            .O(N__35047),
            .I(data_in_1_0));
    LocalMux I__7566 (
            .O(N__35044),
            .I(data_in_1_0));
    LocalMux I__7565 (
            .O(N__35041),
            .I(data_in_1_0));
    InMux I__7564 (
            .O(N__35034),
            .I(N__35031));
    LocalMux I__7563 (
            .O(N__35031),
            .I(N__35027));
    InMux I__7562 (
            .O(N__35030),
            .I(N__35023));
    Span4Mux_h I__7561 (
            .O(N__35027),
            .I(N__35020));
    InMux I__7560 (
            .O(N__35026),
            .I(N__35017));
    LocalMux I__7559 (
            .O(N__35023),
            .I(data_in_0_0));
    Odrv4 I__7558 (
            .O(N__35020),
            .I(data_in_0_0));
    LocalMux I__7557 (
            .O(N__35017),
            .I(data_in_0_0));
    InMux I__7556 (
            .O(N__35010),
            .I(N__35006));
    CascadeMux I__7555 (
            .O(N__35009),
            .I(N__35003));
    LocalMux I__7554 (
            .O(N__35006),
            .I(N__35000));
    InMux I__7553 (
            .O(N__35003),
            .I(N__34996));
    Span4Mux_h I__7552 (
            .O(N__35000),
            .I(N__34993));
    InMux I__7551 (
            .O(N__34999),
            .I(N__34990));
    LocalMux I__7550 (
            .O(N__34996),
            .I(N__34987));
    Odrv4 I__7549 (
            .O(N__34993),
            .I(data_in_3_1));
    LocalMux I__7548 (
            .O(N__34990),
            .I(data_in_3_1));
    Odrv12 I__7547 (
            .O(N__34987),
            .I(data_in_3_1));
    InMux I__7546 (
            .O(N__34980),
            .I(N__34977));
    LocalMux I__7545 (
            .O(N__34977),
            .I(\c0.n2128 ));
    InMux I__7544 (
            .O(N__34974),
            .I(N__34970));
    InMux I__7543 (
            .O(N__34973),
            .I(N__34967));
    LocalMux I__7542 (
            .O(N__34970),
            .I(N__34962));
    LocalMux I__7541 (
            .O(N__34967),
            .I(N__34962));
    Odrv4 I__7540 (
            .O(N__34962),
            .I(data_in_frame_6_7));
    InMux I__7539 (
            .O(N__34959),
            .I(N__34955));
    InMux I__7538 (
            .O(N__34958),
            .I(N__34952));
    LocalMux I__7537 (
            .O(N__34955),
            .I(\c0.data_in_frame_5_0 ));
    LocalMux I__7536 (
            .O(N__34952),
            .I(\c0.data_in_frame_5_0 ));
    CascadeMux I__7535 (
            .O(N__34947),
            .I(\c0.n2128_cascade_ ));
    InMux I__7534 (
            .O(N__34944),
            .I(N__34941));
    LocalMux I__7533 (
            .O(N__34941),
            .I(N__34938));
    Odrv4 I__7532 (
            .O(N__34938),
            .I(\c0.n19_adj_2324 ));
    InMux I__7531 (
            .O(N__34935),
            .I(N__34930));
    InMux I__7530 (
            .O(N__34934),
            .I(N__34927));
    InMux I__7529 (
            .O(N__34933),
            .I(N__34924));
    LocalMux I__7528 (
            .O(N__34930),
            .I(N__34920));
    LocalMux I__7527 (
            .O(N__34927),
            .I(N__34917));
    LocalMux I__7526 (
            .O(N__34924),
            .I(N__34914));
    InMux I__7525 (
            .O(N__34923),
            .I(N__34911));
    Span12Mux_s11_h I__7524 (
            .O(N__34920),
            .I(N__34908));
    Span4Mux_h I__7523 (
            .O(N__34917),
            .I(N__34903));
    Span4Mux_h I__7522 (
            .O(N__34914),
            .I(N__34903));
    LocalMux I__7521 (
            .O(N__34911),
            .I(data_in_3_0));
    Odrv12 I__7520 (
            .O(N__34908),
            .I(data_in_3_0));
    Odrv4 I__7519 (
            .O(N__34903),
            .I(data_in_3_0));
    InMux I__7518 (
            .O(N__34896),
            .I(N__34891));
    InMux I__7517 (
            .O(N__34895),
            .I(N__34887));
    InMux I__7516 (
            .O(N__34894),
            .I(N__34884));
    LocalMux I__7515 (
            .O(N__34891),
            .I(N__34881));
    InMux I__7514 (
            .O(N__34890),
            .I(N__34878));
    LocalMux I__7513 (
            .O(N__34887),
            .I(\c0.data_in_frame_0_3 ));
    LocalMux I__7512 (
            .O(N__34884),
            .I(\c0.data_in_frame_0_3 ));
    Odrv4 I__7511 (
            .O(N__34881),
            .I(\c0.data_in_frame_0_3 ));
    LocalMux I__7510 (
            .O(N__34878),
            .I(\c0.data_in_frame_0_3 ));
    CascadeMux I__7509 (
            .O(N__34869),
            .I(N__34866));
    InMux I__7508 (
            .O(N__34866),
            .I(N__34862));
    CascadeMux I__7507 (
            .O(N__34865),
            .I(N__34859));
    LocalMux I__7506 (
            .O(N__34862),
            .I(N__34856));
    InMux I__7505 (
            .O(N__34859),
            .I(N__34851));
    Span4Mux_v I__7504 (
            .O(N__34856),
            .I(N__34848));
    InMux I__7503 (
            .O(N__34855),
            .I(N__34845));
    InMux I__7502 (
            .O(N__34854),
            .I(N__34842));
    LocalMux I__7501 (
            .O(N__34851),
            .I(\c0.data_in_frame_0_2 ));
    Odrv4 I__7500 (
            .O(N__34848),
            .I(\c0.data_in_frame_0_2 ));
    LocalMux I__7499 (
            .O(N__34845),
            .I(\c0.data_in_frame_0_2 ));
    LocalMux I__7498 (
            .O(N__34842),
            .I(\c0.data_in_frame_0_2 ));
    InMux I__7497 (
            .O(N__34833),
            .I(N__34829));
    InMux I__7496 (
            .O(N__34832),
            .I(N__34826));
    LocalMux I__7495 (
            .O(N__34829),
            .I(N__34821));
    LocalMux I__7494 (
            .O(N__34826),
            .I(N__34821));
    Span4Mux_v I__7493 (
            .O(N__34821),
            .I(N__34817));
    InMux I__7492 (
            .O(N__34820),
            .I(N__34814));
    Odrv4 I__7491 (
            .O(N__34817),
            .I(\c0.n2120 ));
    LocalMux I__7490 (
            .O(N__34814),
            .I(\c0.n2120 ));
    CascadeMux I__7489 (
            .O(N__34809),
            .I(\c0.n22_adj_2201_cascade_ ));
    InMux I__7488 (
            .O(N__34806),
            .I(N__34803));
    LocalMux I__7487 (
            .O(N__34803),
            .I(\c0.n27_adj_2202 ));
    InMux I__7486 (
            .O(N__34800),
            .I(N__34793));
    InMux I__7485 (
            .O(N__34799),
            .I(N__34790));
    InMux I__7484 (
            .O(N__34798),
            .I(N__34785));
    InMux I__7483 (
            .O(N__34797),
            .I(N__34785));
    InMux I__7482 (
            .O(N__34796),
            .I(N__34782));
    LocalMux I__7481 (
            .O(N__34793),
            .I(\c0.data_in_frame_0_5 ));
    LocalMux I__7480 (
            .O(N__34790),
            .I(\c0.data_in_frame_0_5 ));
    LocalMux I__7479 (
            .O(N__34785),
            .I(\c0.data_in_frame_0_5 ));
    LocalMux I__7478 (
            .O(N__34782),
            .I(\c0.data_in_frame_0_5 ));
    InMux I__7477 (
            .O(N__34773),
            .I(N__34768));
    InMux I__7476 (
            .O(N__34772),
            .I(N__34760));
    InMux I__7475 (
            .O(N__34771),
            .I(N__34757));
    LocalMux I__7474 (
            .O(N__34768),
            .I(N__34754));
    InMux I__7473 (
            .O(N__34767),
            .I(N__34751));
    InMux I__7472 (
            .O(N__34766),
            .I(N__34744));
    InMux I__7471 (
            .O(N__34765),
            .I(N__34744));
    InMux I__7470 (
            .O(N__34764),
            .I(N__34744));
    InMux I__7469 (
            .O(N__34763),
            .I(N__34741));
    LocalMux I__7468 (
            .O(N__34760),
            .I(\c0.data_in_frame_0_6 ));
    LocalMux I__7467 (
            .O(N__34757),
            .I(\c0.data_in_frame_0_6 ));
    Odrv12 I__7466 (
            .O(N__34754),
            .I(\c0.data_in_frame_0_6 ));
    LocalMux I__7465 (
            .O(N__34751),
            .I(\c0.data_in_frame_0_6 ));
    LocalMux I__7464 (
            .O(N__34744),
            .I(\c0.data_in_frame_0_6 ));
    LocalMux I__7463 (
            .O(N__34741),
            .I(\c0.data_in_frame_0_6 ));
    CascadeMux I__7462 (
            .O(N__34728),
            .I(\c0.n17469_cascade_ ));
    InMux I__7461 (
            .O(N__34725),
            .I(N__34721));
    InMux I__7460 (
            .O(N__34724),
            .I(N__34718));
    LocalMux I__7459 (
            .O(N__34721),
            .I(N__34715));
    LocalMux I__7458 (
            .O(N__34718),
            .I(N__34711));
    Span4Mux_h I__7457 (
            .O(N__34715),
            .I(N__34707));
    CascadeMux I__7456 (
            .O(N__34714),
            .I(N__34704));
    Span4Mux_v I__7455 (
            .O(N__34711),
            .I(N__34701));
    InMux I__7454 (
            .O(N__34710),
            .I(N__34698));
    Span4Mux_h I__7453 (
            .O(N__34707),
            .I(N__34695));
    InMux I__7452 (
            .O(N__34704),
            .I(N__34692));
    Sp12to4 I__7451 (
            .O(N__34701),
            .I(N__34687));
    LocalMux I__7450 (
            .O(N__34698),
            .I(N__34687));
    Odrv4 I__7449 (
            .O(N__34695),
            .I(\c0.data_out_frame2_0_7 ));
    LocalMux I__7448 (
            .O(N__34692),
            .I(\c0.data_out_frame2_0_7 ));
    Odrv12 I__7447 (
            .O(N__34687),
            .I(\c0.data_out_frame2_0_7 ));
    CascadeMux I__7446 (
            .O(N__34680),
            .I(N__34677));
    InMux I__7445 (
            .O(N__34677),
            .I(N__34674));
    LocalMux I__7444 (
            .O(N__34674),
            .I(N__34670));
    InMux I__7443 (
            .O(N__34673),
            .I(N__34667));
    Span4Mux_h I__7442 (
            .O(N__34670),
            .I(N__34664));
    LocalMux I__7441 (
            .O(N__34667),
            .I(data_in_frame_6_1));
    Odrv4 I__7440 (
            .O(N__34664),
            .I(data_in_frame_6_1));
    InMux I__7439 (
            .O(N__34659),
            .I(N__34656));
    LocalMux I__7438 (
            .O(N__34656),
            .I(N__34652));
    InMux I__7437 (
            .O(N__34655),
            .I(N__34649));
    Span4Mux_h I__7436 (
            .O(N__34652),
            .I(N__34646));
    LocalMux I__7435 (
            .O(N__34649),
            .I(\c0.data_in_frame_5_1 ));
    Odrv4 I__7434 (
            .O(N__34646),
            .I(\c0.data_in_frame_5_1 ));
    CascadeMux I__7433 (
            .O(N__34641),
            .I(\c0.n17114_cascade_ ));
    CascadeMux I__7432 (
            .O(N__34638),
            .I(N__34635));
    InMux I__7431 (
            .O(N__34635),
            .I(N__34632));
    LocalMux I__7430 (
            .O(N__34632),
            .I(N__34629));
    Span4Mux_h I__7429 (
            .O(N__34629),
            .I(N__34625));
    InMux I__7428 (
            .O(N__34628),
            .I(N__34622));
    Span4Mux_h I__7427 (
            .O(N__34625),
            .I(N__34619));
    LocalMux I__7426 (
            .O(N__34622),
            .I(\c0.data_in_frame_5_7 ));
    Odrv4 I__7425 (
            .O(N__34619),
            .I(\c0.data_in_frame_5_7 ));
    CascadeMux I__7424 (
            .O(N__34614),
            .I(N__34610));
    InMux I__7423 (
            .O(N__34613),
            .I(N__34604));
    InMux I__7422 (
            .O(N__34610),
            .I(N__34601));
    InMux I__7421 (
            .O(N__34609),
            .I(N__34596));
    InMux I__7420 (
            .O(N__34608),
            .I(N__34596));
    InMux I__7419 (
            .O(N__34607),
            .I(N__34593));
    LocalMux I__7418 (
            .O(N__34604),
            .I(N__34590));
    LocalMux I__7417 (
            .O(N__34601),
            .I(\c0.data_in_frame_1_4 ));
    LocalMux I__7416 (
            .O(N__34596),
            .I(\c0.data_in_frame_1_4 ));
    LocalMux I__7415 (
            .O(N__34593),
            .I(\c0.data_in_frame_1_4 ));
    Odrv4 I__7414 (
            .O(N__34590),
            .I(\c0.data_in_frame_1_4 ));
    CascadeMux I__7413 (
            .O(N__34581),
            .I(\c0.n17101_cascade_ ));
    CascadeMux I__7412 (
            .O(N__34578),
            .I(\c0.n10_adj_2299_cascade_ ));
    InMux I__7411 (
            .O(N__34575),
            .I(N__34571));
    InMux I__7410 (
            .O(N__34574),
            .I(N__34568));
    LocalMux I__7409 (
            .O(N__34571),
            .I(\c0.n17206 ));
    LocalMux I__7408 (
            .O(N__34568),
            .I(\c0.n17206 ));
    InMux I__7407 (
            .O(N__34563),
            .I(N__34557));
    InMux I__7406 (
            .O(N__34562),
            .I(N__34557));
    LocalMux I__7405 (
            .O(N__34557),
            .I(\c0.n10407 ));
    InMux I__7404 (
            .O(N__34554),
            .I(N__34551));
    LocalMux I__7403 (
            .O(N__34551),
            .I(N__34547));
    InMux I__7402 (
            .O(N__34550),
            .I(N__34544));
    Span4Mux_h I__7401 (
            .O(N__34547),
            .I(N__34541));
    LocalMux I__7400 (
            .O(N__34544),
            .I(N__34536));
    Span4Mux_h I__7399 (
            .O(N__34541),
            .I(N__34536));
    Odrv4 I__7398 (
            .O(N__34536),
            .I(data_in_frame_6_0));
    CascadeMux I__7397 (
            .O(N__34533),
            .I(\c0.n10407_cascade_ ));
    InMux I__7396 (
            .O(N__34530),
            .I(N__34523));
    InMux I__7395 (
            .O(N__34529),
            .I(N__34523));
    InMux I__7394 (
            .O(N__34528),
            .I(N__34518));
    LocalMux I__7393 (
            .O(N__34523),
            .I(N__34515));
    CascadeMux I__7392 (
            .O(N__34522),
            .I(N__34512));
    InMux I__7391 (
            .O(N__34521),
            .I(N__34509));
    LocalMux I__7390 (
            .O(N__34518),
            .I(N__34506));
    Span4Mux_v I__7389 (
            .O(N__34515),
            .I(N__34503));
    InMux I__7388 (
            .O(N__34512),
            .I(N__34500));
    LocalMux I__7387 (
            .O(N__34509),
            .I(\c0.data_in_frame_1_5 ));
    Odrv4 I__7386 (
            .O(N__34506),
            .I(\c0.data_in_frame_1_5 ));
    Odrv4 I__7385 (
            .O(N__34503),
            .I(\c0.data_in_frame_1_5 ));
    LocalMux I__7384 (
            .O(N__34500),
            .I(\c0.data_in_frame_1_5 ));
    InMux I__7383 (
            .O(N__34491),
            .I(N__34488));
    LocalMux I__7382 (
            .O(N__34488),
            .I(\c0.n17215 ));
    InMux I__7381 (
            .O(N__34485),
            .I(N__34481));
    InMux I__7380 (
            .O(N__34484),
            .I(N__34478));
    LocalMux I__7379 (
            .O(N__34481),
            .I(N__34471));
    LocalMux I__7378 (
            .O(N__34478),
            .I(N__34471));
    CascadeMux I__7377 (
            .O(N__34477),
            .I(N__34468));
    InMux I__7376 (
            .O(N__34476),
            .I(N__34465));
    Span4Mux_h I__7375 (
            .O(N__34471),
            .I(N__34462));
    InMux I__7374 (
            .O(N__34468),
            .I(N__34459));
    LocalMux I__7373 (
            .O(N__34465),
            .I(N__34456));
    Span4Mux_h I__7372 (
            .O(N__34462),
            .I(N__34453));
    LocalMux I__7371 (
            .O(N__34459),
            .I(\c0.byte_transmit_counter2_7 ));
    Odrv12 I__7370 (
            .O(N__34456),
            .I(\c0.byte_transmit_counter2_7 ));
    Odrv4 I__7369 (
            .O(N__34453),
            .I(\c0.byte_transmit_counter2_7 ));
    InMux I__7368 (
            .O(N__34446),
            .I(N__34443));
    LocalMux I__7367 (
            .O(N__34443),
            .I(N__34438));
    InMux I__7366 (
            .O(N__34442),
            .I(N__34434));
    InMux I__7365 (
            .O(N__34441),
            .I(N__34431));
    Span4Mux_h I__7364 (
            .O(N__34438),
            .I(N__34428));
    InMux I__7363 (
            .O(N__34437),
            .I(N__34425));
    LocalMux I__7362 (
            .O(N__34434),
            .I(\c0.byte_transmit_counter2_6 ));
    LocalMux I__7361 (
            .O(N__34431),
            .I(\c0.byte_transmit_counter2_6 ));
    Odrv4 I__7360 (
            .O(N__34428),
            .I(\c0.byte_transmit_counter2_6 ));
    LocalMux I__7359 (
            .O(N__34425),
            .I(\c0.byte_transmit_counter2_6 ));
    InMux I__7358 (
            .O(N__34416),
            .I(N__34413));
    LocalMux I__7357 (
            .O(N__34413),
            .I(\c0.n13284 ));
    InMux I__7356 (
            .O(N__34410),
            .I(N__34404));
    InMux I__7355 (
            .O(N__34409),
            .I(N__34404));
    LocalMux I__7354 (
            .O(N__34404),
            .I(\c0.n13628 ));
    CascadeMux I__7353 (
            .O(N__34401),
            .I(\c0.n13628_cascade_ ));
    InMux I__7352 (
            .O(N__34398),
            .I(N__34392));
    InMux I__7351 (
            .O(N__34397),
            .I(N__34387));
    InMux I__7350 (
            .O(N__34396),
            .I(N__34387));
    CascadeMux I__7349 (
            .O(N__34395),
            .I(N__34384));
    LocalMux I__7348 (
            .O(N__34392),
            .I(N__34379));
    LocalMux I__7347 (
            .O(N__34387),
            .I(N__34379));
    InMux I__7346 (
            .O(N__34384),
            .I(N__34376));
    Span4Mux_h I__7345 (
            .O(N__34379),
            .I(N__34373));
    LocalMux I__7344 (
            .O(N__34376),
            .I(tx2_active));
    Odrv4 I__7343 (
            .O(N__34373),
            .I(tx2_active));
    InMux I__7342 (
            .O(N__34368),
            .I(N__34365));
    LocalMux I__7341 (
            .O(N__34365),
            .I(N__34361));
    InMux I__7340 (
            .O(N__34364),
            .I(N__34358));
    Span4Mux_h I__7339 (
            .O(N__34361),
            .I(N__34355));
    LocalMux I__7338 (
            .O(N__34358),
            .I(\c0.data_in_frame_3_2 ));
    Odrv4 I__7337 (
            .O(N__34355),
            .I(\c0.data_in_frame_3_2 ));
    CascadeMux I__7336 (
            .O(N__34350),
            .I(N__34347));
    InMux I__7335 (
            .O(N__34347),
            .I(N__34344));
    LocalMux I__7334 (
            .O(N__34344),
            .I(N__34340));
    InMux I__7333 (
            .O(N__34343),
            .I(N__34337));
    Span4Mux_v I__7332 (
            .O(N__34340),
            .I(N__34334));
    LocalMux I__7331 (
            .O(N__34337),
            .I(data_in_frame_6_2));
    Odrv4 I__7330 (
            .O(N__34334),
            .I(data_in_frame_6_2));
    CascadeMux I__7329 (
            .O(N__34329),
            .I(\c0.n17475_cascade_ ));
    InMux I__7328 (
            .O(N__34326),
            .I(N__34322));
    CascadeMux I__7327 (
            .O(N__34325),
            .I(N__34319));
    LocalMux I__7326 (
            .O(N__34322),
            .I(N__34315));
    InMux I__7325 (
            .O(N__34319),
            .I(N__34309));
    InMux I__7324 (
            .O(N__34318),
            .I(N__34309));
    Span4Mux_h I__7323 (
            .O(N__34315),
            .I(N__34306));
    CascadeMux I__7322 (
            .O(N__34314),
            .I(N__34303));
    LocalMux I__7321 (
            .O(N__34309),
            .I(N__34300));
    Span4Mux_h I__7320 (
            .O(N__34306),
            .I(N__34297));
    InMux I__7319 (
            .O(N__34303),
            .I(N__34294));
    Span12Mux_s4_h I__7318 (
            .O(N__34300),
            .I(N__34291));
    Span4Mux_h I__7317 (
            .O(N__34297),
            .I(N__34288));
    LocalMux I__7316 (
            .O(N__34294),
            .I(\c0.data_out_frame2_0_5 ));
    Odrv12 I__7315 (
            .O(N__34291),
            .I(\c0.data_out_frame2_0_5 ));
    Odrv4 I__7314 (
            .O(N__34288),
            .I(\c0.data_out_frame2_0_5 ));
    InMux I__7313 (
            .O(N__34281),
            .I(N__34278));
    LocalMux I__7312 (
            .O(N__34278),
            .I(N__34275));
    Span4Mux_v I__7311 (
            .O(N__34275),
            .I(N__34272));
    Odrv4 I__7310 (
            .O(N__34272),
            .I(\c0.n16352 ));
    InMux I__7309 (
            .O(N__34269),
            .I(N__34266));
    LocalMux I__7308 (
            .O(N__34266),
            .I(\c0.n24_adj_2340 ));
    CascadeMux I__7307 (
            .O(N__34263),
            .I(N__34260));
    InMux I__7306 (
            .O(N__34260),
            .I(N__34257));
    LocalMux I__7305 (
            .O(N__34257),
            .I(N__34254));
    Span4Mux_h I__7304 (
            .O(N__34254),
            .I(N__34250));
    InMux I__7303 (
            .O(N__34253),
            .I(N__34247));
    Sp12to4 I__7302 (
            .O(N__34250),
            .I(N__34244));
    LocalMux I__7301 (
            .O(N__34247),
            .I(data_in_frame_6_5));
    Odrv12 I__7300 (
            .O(N__34244),
            .I(data_in_frame_6_5));
    InMux I__7299 (
            .O(N__34239),
            .I(N__34233));
    InMux I__7298 (
            .O(N__34238),
            .I(N__34233));
    LocalMux I__7297 (
            .O(N__34233),
            .I(N__34230));
    Odrv4 I__7296 (
            .O(N__34230),
            .I(\c0.n2122 ));
    InMux I__7295 (
            .O(N__34227),
            .I(N__34223));
    InMux I__7294 (
            .O(N__34226),
            .I(N__34220));
    LocalMux I__7293 (
            .O(N__34223),
            .I(data_out_0_5));
    LocalMux I__7292 (
            .O(N__34220),
            .I(data_out_0_5));
    InMux I__7291 (
            .O(N__34215),
            .I(N__34211));
    InMux I__7290 (
            .O(N__34214),
            .I(N__34208));
    LocalMux I__7289 (
            .O(N__34211),
            .I(data_out_2_2));
    LocalMux I__7288 (
            .O(N__34208),
            .I(data_out_2_2));
    CascadeMux I__7287 (
            .O(N__34203),
            .I(n2699_cascade_));
    InMux I__7286 (
            .O(N__34200),
            .I(N__34196));
    InMux I__7285 (
            .O(N__34199),
            .I(N__34193));
    LocalMux I__7284 (
            .O(N__34196),
            .I(N__34190));
    LocalMux I__7283 (
            .O(N__34193),
            .I(data_out_3_4));
    Odrv4 I__7282 (
            .O(N__34190),
            .I(data_out_3_4));
    InMux I__7281 (
            .O(N__34185),
            .I(N__34176));
    InMux I__7280 (
            .O(N__34184),
            .I(N__34176));
    InMux I__7279 (
            .O(N__34183),
            .I(N__34176));
    LocalMux I__7278 (
            .O(N__34176),
            .I(n2699));
    InMux I__7277 (
            .O(N__34173),
            .I(N__34169));
    InMux I__7276 (
            .O(N__34172),
            .I(N__34166));
    LocalMux I__7275 (
            .O(N__34169),
            .I(data_out_3_2));
    LocalMux I__7274 (
            .O(N__34166),
            .I(data_out_3_2));
    InMux I__7273 (
            .O(N__34161),
            .I(N__34157));
    InMux I__7272 (
            .O(N__34160),
            .I(N__34154));
    LocalMux I__7271 (
            .O(N__34157),
            .I(N__34150));
    LocalMux I__7270 (
            .O(N__34154),
            .I(N__34147));
    InMux I__7269 (
            .O(N__34153),
            .I(N__34144));
    Span4Mux_v I__7268 (
            .O(N__34150),
            .I(N__34141));
    Span4Mux_h I__7267 (
            .O(N__34147),
            .I(N__34138));
    LocalMux I__7266 (
            .O(N__34144),
            .I(\c0.data_in_frame_2_6 ));
    Odrv4 I__7265 (
            .O(N__34141),
            .I(\c0.data_in_frame_2_6 ));
    Odrv4 I__7264 (
            .O(N__34138),
            .I(\c0.data_in_frame_2_6 ));
    InMux I__7263 (
            .O(N__34131),
            .I(N__34128));
    LocalMux I__7262 (
            .O(N__34128),
            .I(N__34125));
    Span4Mux_h I__7261 (
            .O(N__34125),
            .I(N__34122));
    Odrv4 I__7260 (
            .O(N__34122),
            .I(\c0.n17713 ));
    SRMux I__7259 (
            .O(N__34119),
            .I(N__34116));
    LocalMux I__7258 (
            .O(N__34116),
            .I(\c0.n4_adj_2325 ));
    InMux I__7257 (
            .O(N__34113),
            .I(N__34099));
    InMux I__7256 (
            .O(N__34112),
            .I(N__34099));
    InMux I__7255 (
            .O(N__34111),
            .I(N__34099));
    InMux I__7254 (
            .O(N__34110),
            .I(N__34088));
    InMux I__7253 (
            .O(N__34109),
            .I(N__34088));
    InMux I__7252 (
            .O(N__34108),
            .I(N__34088));
    InMux I__7251 (
            .O(N__34107),
            .I(N__34088));
    InMux I__7250 (
            .O(N__34106),
            .I(N__34088));
    LocalMux I__7249 (
            .O(N__34099),
            .I(N__34083));
    LocalMux I__7248 (
            .O(N__34088),
            .I(N__34083));
    Odrv12 I__7247 (
            .O(N__34083),
            .I(\c0.tx2_transmit_N_1996 ));
    InMux I__7246 (
            .O(N__34080),
            .I(N__34077));
    LocalMux I__7245 (
            .O(N__34077),
            .I(\c0.n17676 ));
    CascadeMux I__7244 (
            .O(N__34074),
            .I(N__34071));
    InMux I__7243 (
            .O(N__34071),
            .I(N__34068));
    LocalMux I__7242 (
            .O(N__34068),
            .I(N__34064));
    CascadeMux I__7241 (
            .O(N__34067),
            .I(N__34061));
    Span4Mux_v I__7240 (
            .O(N__34064),
            .I(N__34058));
    InMux I__7239 (
            .O(N__34061),
            .I(N__34055));
    Odrv4 I__7238 (
            .O(N__34058),
            .I(rand_setpoint_14));
    LocalMux I__7237 (
            .O(N__34055),
            .I(rand_setpoint_14));
    InMux I__7236 (
            .O(N__34050),
            .I(N__34047));
    LocalMux I__7235 (
            .O(N__34047),
            .I(\c0.n17703 ));
    InMux I__7234 (
            .O(N__34044),
            .I(N__34038));
    InMux I__7233 (
            .O(N__34043),
            .I(N__34038));
    LocalMux I__7232 (
            .O(N__34038),
            .I(\c0.data_out_1_4 ));
    InMux I__7231 (
            .O(N__34035),
            .I(N__34032));
    LocalMux I__7230 (
            .O(N__34032),
            .I(\c0.n17675 ));
    InMux I__7229 (
            .O(N__34029),
            .I(N__34026));
    LocalMux I__7228 (
            .O(N__34026),
            .I(N__34023));
    Odrv4 I__7227 (
            .O(N__34023),
            .I(\c0.n17697 ));
    InMux I__7226 (
            .O(N__34020),
            .I(N__34017));
    LocalMux I__7225 (
            .O(N__34017),
            .I(N__34014));
    Odrv4 I__7224 (
            .O(N__34014),
            .I(n18271));
    CascadeMux I__7223 (
            .O(N__34011),
            .I(n10_adj_2408_cascade_));
    InMux I__7222 (
            .O(N__34008),
            .I(N__34002));
    InMux I__7221 (
            .O(N__34007),
            .I(N__34002));
    LocalMux I__7220 (
            .O(N__34002),
            .I(\c0.data_out_2_3 ));
    CascadeMux I__7219 (
            .O(N__33999),
            .I(\c0.n18268_cascade_ ));
    CascadeMux I__7218 (
            .O(N__33996),
            .I(\c0.tx.n55_cascade_ ));
    CascadeMux I__7217 (
            .O(N__33993),
            .I(N__33990));
    InMux I__7216 (
            .O(N__33990),
            .I(N__33987));
    LocalMux I__7215 (
            .O(N__33987),
            .I(\c0.n5_adj_2136 ));
    InMux I__7214 (
            .O(N__33984),
            .I(N__33980));
    CascadeMux I__7213 (
            .O(N__33983),
            .I(N__33977));
    LocalMux I__7212 (
            .O(N__33980),
            .I(N__33974));
    InMux I__7211 (
            .O(N__33977),
            .I(N__33971));
    Odrv4 I__7210 (
            .O(N__33974),
            .I(rand_setpoint_12));
    LocalMux I__7209 (
            .O(N__33971),
            .I(rand_setpoint_12));
    CascadeMux I__7208 (
            .O(N__33966),
            .I(N__33963));
    InMux I__7207 (
            .O(N__33963),
            .I(N__33960));
    LocalMux I__7206 (
            .O(N__33960),
            .I(\c0.n5 ));
    CascadeMux I__7205 (
            .O(N__33957),
            .I(\c0.n18172_cascade_ ));
    InMux I__7204 (
            .O(N__33954),
            .I(N__33951));
    LocalMux I__7203 (
            .O(N__33951),
            .I(\c0.n17764 ));
    CascadeMux I__7202 (
            .O(N__33948),
            .I(\c0.n17639_cascade_ ));
    CascadeMux I__7201 (
            .O(N__33945),
            .I(N__33941));
    InMux I__7200 (
            .O(N__33944),
            .I(N__33938));
    InMux I__7199 (
            .O(N__33941),
            .I(N__33935));
    LocalMux I__7198 (
            .O(N__33938),
            .I(rand_setpoint_20));
    LocalMux I__7197 (
            .O(N__33935),
            .I(rand_setpoint_20));
    CascadeMux I__7196 (
            .O(N__33930),
            .I(N__33926));
    InMux I__7195 (
            .O(N__33929),
            .I(N__33923));
    InMux I__7194 (
            .O(N__33926),
            .I(N__33920));
    LocalMux I__7193 (
            .O(N__33923),
            .I(rand_setpoint_22));
    LocalMux I__7192 (
            .O(N__33920),
            .I(rand_setpoint_22));
    CascadeMux I__7191 (
            .O(N__33915),
            .I(N__33912));
    InMux I__7190 (
            .O(N__33912),
            .I(N__33909));
    LocalMux I__7189 (
            .O(N__33909),
            .I(N__33906));
    Span4Mux_h I__7188 (
            .O(N__33906),
            .I(N__33903));
    Odrv4 I__7187 (
            .O(N__33903),
            .I(\c0.n17647 ));
    CascadeMux I__7186 (
            .O(N__33900),
            .I(N__33896));
    InMux I__7185 (
            .O(N__33899),
            .I(N__33893));
    InMux I__7184 (
            .O(N__33896),
            .I(N__33890));
    LocalMux I__7183 (
            .O(N__33893),
            .I(rand_setpoint_19));
    LocalMux I__7182 (
            .O(N__33890),
            .I(rand_setpoint_19));
    CascadeMux I__7181 (
            .O(N__33885),
            .I(\c0.n17631_cascade_ ));
    CascadeMux I__7180 (
            .O(N__33882),
            .I(N__33878));
    InMux I__7179 (
            .O(N__33881),
            .I(N__33875));
    InMux I__7178 (
            .O(N__33878),
            .I(N__33872));
    LocalMux I__7177 (
            .O(N__33875),
            .I(rand_setpoint_18));
    LocalMux I__7176 (
            .O(N__33872),
            .I(rand_setpoint_18));
    CascadeMux I__7175 (
            .O(N__33867),
            .I(\c0.n17627_cascade_ ));
    CascadeMux I__7174 (
            .O(N__33864),
            .I(N__33860));
    InMux I__7173 (
            .O(N__33863),
            .I(N__33857));
    InMux I__7172 (
            .O(N__33860),
            .I(N__33854));
    LocalMux I__7171 (
            .O(N__33857),
            .I(rand_setpoint_21));
    LocalMux I__7170 (
            .O(N__33854),
            .I(rand_setpoint_21));
    CascadeMux I__7169 (
            .O(N__33849),
            .I(N__33846));
    InMux I__7168 (
            .O(N__33846),
            .I(N__33843));
    LocalMux I__7167 (
            .O(N__33843),
            .I(N__33840));
    Span4Mux_v I__7166 (
            .O(N__33840),
            .I(N__33837));
    Span4Mux_h I__7165 (
            .O(N__33837),
            .I(N__33834));
    Odrv4 I__7164 (
            .O(N__33834),
            .I(\c0.n17643 ));
    CascadeMux I__7163 (
            .O(N__33831),
            .I(N__33827));
    InMux I__7162 (
            .O(N__33830),
            .I(N__33824));
    InMux I__7161 (
            .O(N__33827),
            .I(N__33821));
    LocalMux I__7160 (
            .O(N__33824),
            .I(rand_setpoint_2));
    LocalMux I__7159 (
            .O(N__33821),
            .I(rand_setpoint_2));
    InMux I__7158 (
            .O(N__33816),
            .I(N__33812));
    CascadeMux I__7157 (
            .O(N__33815),
            .I(N__33809));
    LocalMux I__7156 (
            .O(N__33812),
            .I(N__33806));
    InMux I__7155 (
            .O(N__33809),
            .I(N__33803));
    Odrv4 I__7154 (
            .O(N__33806),
            .I(rand_setpoint_3));
    LocalMux I__7153 (
            .O(N__33803),
            .I(rand_setpoint_3));
    CascadeMux I__7152 (
            .O(N__33798),
            .I(N__33795));
    InMux I__7151 (
            .O(N__33795),
            .I(N__33790));
    InMux I__7150 (
            .O(N__33794),
            .I(N__33787));
    InMux I__7149 (
            .O(N__33793),
            .I(N__33784));
    LocalMux I__7148 (
            .O(N__33790),
            .I(\c0.FRAME_MATCHER_state_7 ));
    LocalMux I__7147 (
            .O(N__33787),
            .I(\c0.FRAME_MATCHER_state_7 ));
    LocalMux I__7146 (
            .O(N__33784),
            .I(\c0.FRAME_MATCHER_state_7 ));
    SRMux I__7145 (
            .O(N__33777),
            .I(N__33774));
    LocalMux I__7144 (
            .O(N__33774),
            .I(N__33771));
    Span4Mux_h I__7143 (
            .O(N__33771),
            .I(N__33768));
    Odrv4 I__7142 (
            .O(N__33768),
            .I(\c0.n16141 ));
    InMux I__7141 (
            .O(N__33765),
            .I(N__33761));
    CascadeMux I__7140 (
            .O(N__33764),
            .I(N__33758));
    LocalMux I__7139 (
            .O(N__33761),
            .I(N__33755));
    InMux I__7138 (
            .O(N__33758),
            .I(N__33752));
    Odrv4 I__7137 (
            .O(N__33755),
            .I(rand_setpoint_23));
    LocalMux I__7136 (
            .O(N__33752),
            .I(rand_setpoint_23));
    CascadeMux I__7135 (
            .O(N__33747),
            .I(n21_adj_2487_cascade_));
    InMux I__7134 (
            .O(N__33744),
            .I(N__33741));
    LocalMux I__7133 (
            .O(N__33741),
            .I(N__33736));
    CascadeMux I__7132 (
            .O(N__33740),
            .I(N__33733));
    CascadeMux I__7131 (
            .O(N__33739),
            .I(N__33729));
    Span4Mux_v I__7130 (
            .O(N__33736),
            .I(N__33725));
    InMux I__7129 (
            .O(N__33733),
            .I(N__33720));
    InMux I__7128 (
            .O(N__33732),
            .I(N__33720));
    InMux I__7127 (
            .O(N__33729),
            .I(N__33715));
    InMux I__7126 (
            .O(N__33728),
            .I(N__33715));
    Odrv4 I__7125 (
            .O(N__33725),
            .I(n63_adj_2418));
    LocalMux I__7124 (
            .O(N__33720),
            .I(n63_adj_2418));
    LocalMux I__7123 (
            .O(N__33715),
            .I(n63_adj_2418));
    InMux I__7122 (
            .O(N__33708),
            .I(N__33705));
    LocalMux I__7121 (
            .O(N__33705),
            .I(n6_adj_2410));
    InMux I__7120 (
            .O(N__33702),
            .I(N__33699));
    LocalMux I__7119 (
            .O(N__33699),
            .I(N__33695));
    InMux I__7118 (
            .O(N__33698),
            .I(N__33692));
    Odrv4 I__7117 (
            .O(N__33695),
            .I(n2061));
    LocalMux I__7116 (
            .O(N__33692),
            .I(n2061));
    CascadeMux I__7115 (
            .O(N__33687),
            .I(N__33684));
    InMux I__7114 (
            .O(N__33684),
            .I(N__33681));
    LocalMux I__7113 (
            .O(N__33681),
            .I(N__33678));
    Span4Mux_h I__7112 (
            .O(N__33678),
            .I(N__33675));
    Span4Mux_h I__7111 (
            .O(N__33675),
            .I(N__33672));
    Odrv4 I__7110 (
            .O(N__33672),
            .I(\c0.n51_adj_2173 ));
    InMux I__7109 (
            .O(N__33669),
            .I(N__33666));
    LocalMux I__7108 (
            .O(N__33666),
            .I(N__33663));
    Span4Mux_h I__7107 (
            .O(N__33663),
            .I(N__33660));
    Odrv4 I__7106 (
            .O(N__33660),
            .I(\c0.n10166 ));
    CascadeMux I__7105 (
            .O(N__33657),
            .I(N__33652));
    InMux I__7104 (
            .O(N__33656),
            .I(N__33648));
    InMux I__7103 (
            .O(N__33655),
            .I(N__33643));
    InMux I__7102 (
            .O(N__33652),
            .I(N__33643));
    InMux I__7101 (
            .O(N__33651),
            .I(N__33640));
    LocalMux I__7100 (
            .O(N__33648),
            .I(N__33637));
    LocalMux I__7099 (
            .O(N__33643),
            .I(N__33634));
    LocalMux I__7098 (
            .O(N__33640),
            .I(N__33631));
    Span12Mux_v I__7097 (
            .O(N__33637),
            .I(N__33628));
    Span4Mux_v I__7096 (
            .O(N__33634),
            .I(N__33625));
    Odrv4 I__7095 (
            .O(N__33631),
            .I(\c0.FRAME_MATCHER_i_30 ));
    Odrv12 I__7094 (
            .O(N__33628),
            .I(\c0.FRAME_MATCHER_i_30 ));
    Odrv4 I__7093 (
            .O(N__33625),
            .I(\c0.FRAME_MATCHER_i_30 ));
    InMux I__7092 (
            .O(N__33618),
            .I(N__33615));
    LocalMux I__7091 (
            .O(N__33615),
            .I(N__33612));
    Span4Mux_v I__7090 (
            .O(N__33612),
            .I(N__33609));
    Span4Mux_h I__7089 (
            .O(N__33609),
            .I(N__33606));
    Span4Mux_h I__7088 (
            .O(N__33606),
            .I(N__33603));
    Odrv4 I__7087 (
            .O(N__33603),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_30 ));
    SRMux I__7086 (
            .O(N__33600),
            .I(N__33597));
    LocalMux I__7085 (
            .O(N__33597),
            .I(N__33594));
    Span4Mux_h I__7084 (
            .O(N__33594),
            .I(N__33591));
    Span4Mux_h I__7083 (
            .O(N__33591),
            .I(N__33588));
    Odrv4 I__7082 (
            .O(N__33588),
            .I(\c0.n16696 ));
    CascadeMux I__7081 (
            .O(N__33585),
            .I(\c0.n8_adj_2385_cascade_ ));
    SRMux I__7080 (
            .O(N__33582),
            .I(N__33579));
    LocalMux I__7079 (
            .O(N__33579),
            .I(N__33576));
    Span4Mux_s2_v I__7078 (
            .O(N__33576),
            .I(N__33573));
    Span4Mux_h I__7077 (
            .O(N__33573),
            .I(N__33570));
    Span4Mux_h I__7076 (
            .O(N__33570),
            .I(N__33567));
    Span4Mux_v I__7075 (
            .O(N__33567),
            .I(N__33564));
    Odrv4 I__7074 (
            .O(N__33564),
            .I(\c0.n16670 ));
    CascadeMux I__7073 (
            .O(N__33561),
            .I(\c0.n17367_cascade_ ));
    CascadeMux I__7072 (
            .O(N__33558),
            .I(n9_cascade_));
    InMux I__7071 (
            .O(N__33555),
            .I(N__33550));
    InMux I__7070 (
            .O(N__33554),
            .I(N__33547));
    InMux I__7069 (
            .O(N__33553),
            .I(N__33544));
    LocalMux I__7068 (
            .O(N__33550),
            .I(\c0.n10139 ));
    LocalMux I__7067 (
            .O(N__33547),
            .I(\c0.n10139 ));
    LocalMux I__7066 (
            .O(N__33544),
            .I(\c0.n10139 ));
    InMux I__7065 (
            .O(N__33537),
            .I(N__33531));
    InMux I__7064 (
            .O(N__33536),
            .I(N__33528));
    InMux I__7063 (
            .O(N__33535),
            .I(N__33523));
    InMux I__7062 (
            .O(N__33534),
            .I(N__33523));
    LocalMux I__7061 (
            .O(N__33531),
            .I(N__33516));
    LocalMux I__7060 (
            .O(N__33528),
            .I(N__33511));
    LocalMux I__7059 (
            .O(N__33523),
            .I(N__33511));
    InMux I__7058 (
            .O(N__33522),
            .I(N__33502));
    InMux I__7057 (
            .O(N__33521),
            .I(N__33502));
    InMux I__7056 (
            .O(N__33520),
            .I(N__33502));
    InMux I__7055 (
            .O(N__33519),
            .I(N__33502));
    Span4Mux_h I__7054 (
            .O(N__33516),
            .I(N__33499));
    Sp12to4 I__7053 (
            .O(N__33511),
            .I(N__33494));
    LocalMux I__7052 (
            .O(N__33502),
            .I(N__33494));
    Odrv4 I__7051 (
            .O(N__33499),
            .I(\c0.n11833 ));
    Odrv12 I__7050 (
            .O(N__33494),
            .I(\c0.n11833 ));
    InMux I__7049 (
            .O(N__33489),
            .I(N__33484));
    InMux I__7048 (
            .O(N__33488),
            .I(N__33479));
    InMux I__7047 (
            .O(N__33487),
            .I(N__33479));
    LocalMux I__7046 (
            .O(N__33484),
            .I(N__33476));
    LocalMux I__7045 (
            .O(N__33479),
            .I(\c0.FRAME_MATCHER_state_3 ));
    Odrv4 I__7044 (
            .O(N__33476),
            .I(\c0.FRAME_MATCHER_state_3 ));
    InMux I__7043 (
            .O(N__33471),
            .I(N__33466));
    InMux I__7042 (
            .O(N__33470),
            .I(N__33463));
    CascadeMux I__7041 (
            .O(N__33469),
            .I(N__33460));
    LocalMux I__7040 (
            .O(N__33466),
            .I(N__33455));
    LocalMux I__7039 (
            .O(N__33463),
            .I(N__33455));
    InMux I__7038 (
            .O(N__33460),
            .I(N__33452));
    Span4Mux_h I__7037 (
            .O(N__33455),
            .I(N__33449));
    LocalMux I__7036 (
            .O(N__33452),
            .I(\c0.FRAME_MATCHER_state_5 ));
    Odrv4 I__7035 (
            .O(N__33449),
            .I(\c0.FRAME_MATCHER_state_5 ));
    InMux I__7034 (
            .O(N__33444),
            .I(N__33441));
    LocalMux I__7033 (
            .O(N__33441),
            .I(N__33438));
    Span4Mux_v I__7032 (
            .O(N__33438),
            .I(N__33433));
    InMux I__7031 (
            .O(N__33437),
            .I(N__33430));
    InMux I__7030 (
            .O(N__33436),
            .I(N__33427));
    Span4Mux_h I__7029 (
            .O(N__33433),
            .I(N__33422));
    LocalMux I__7028 (
            .O(N__33430),
            .I(N__33422));
    LocalMux I__7027 (
            .O(N__33427),
            .I(n9));
    Odrv4 I__7026 (
            .O(N__33422),
            .I(n9));
    CascadeMux I__7025 (
            .O(N__33417),
            .I(N__33413));
    InMux I__7024 (
            .O(N__33416),
            .I(N__33409));
    InMux I__7023 (
            .O(N__33413),
            .I(N__33406));
    InMux I__7022 (
            .O(N__33412),
            .I(N__33403));
    LocalMux I__7021 (
            .O(N__33409),
            .I(N__33400));
    LocalMux I__7020 (
            .O(N__33406),
            .I(N__33397));
    LocalMux I__7019 (
            .O(N__33403),
            .I(\c0.data_in_frame_2_4 ));
    Odrv12 I__7018 (
            .O(N__33400),
            .I(\c0.data_in_frame_2_4 ));
    Odrv4 I__7017 (
            .O(N__33397),
            .I(\c0.data_in_frame_2_4 ));
    CascadeMux I__7016 (
            .O(N__33390),
            .I(FRAME_MATCHER_i_31__N_1273_cascade_));
    CascadeMux I__7015 (
            .O(N__33387),
            .I(n17086_cascade_));
    InMux I__7014 (
            .O(N__33384),
            .I(N__33375));
    InMux I__7013 (
            .O(N__33383),
            .I(N__33375));
    InMux I__7012 (
            .O(N__33382),
            .I(N__33372));
    InMux I__7011 (
            .O(N__33381),
            .I(N__33367));
    InMux I__7010 (
            .O(N__33380),
            .I(N__33367));
    LocalMux I__7009 (
            .O(N__33375),
            .I(n63_adj_2428));
    LocalMux I__7008 (
            .O(N__33372),
            .I(n63_adj_2428));
    LocalMux I__7007 (
            .O(N__33367),
            .I(n63_adj_2428));
    InMux I__7006 (
            .O(N__33360),
            .I(N__33356));
    InMux I__7005 (
            .O(N__33359),
            .I(N__33351));
    LocalMux I__7004 (
            .O(N__33356),
            .I(N__33348));
    InMux I__7003 (
            .O(N__33355),
            .I(N__33343));
    InMux I__7002 (
            .O(N__33354),
            .I(N__33343));
    LocalMux I__7001 (
            .O(N__33351),
            .I(n63));
    Odrv4 I__7000 (
            .O(N__33348),
            .I(n63));
    LocalMux I__6999 (
            .O(N__33343),
            .I(n63));
    InMux I__6998 (
            .O(N__33336),
            .I(N__33333));
    LocalMux I__6997 (
            .O(N__33333),
            .I(N__33329));
    CascadeMux I__6996 (
            .O(N__33332),
            .I(N__33326));
    Span4Mux_v I__6995 (
            .O(N__33329),
            .I(N__33323));
    InMux I__6994 (
            .O(N__33326),
            .I(N__33319));
    Span4Mux_h I__6993 (
            .O(N__33323),
            .I(N__33316));
    InMux I__6992 (
            .O(N__33322),
            .I(N__33313));
    LocalMux I__6991 (
            .O(N__33319),
            .I(\c0.FRAME_MATCHER_state_8 ));
    Odrv4 I__6990 (
            .O(N__33316),
            .I(\c0.FRAME_MATCHER_state_8 ));
    LocalMux I__6989 (
            .O(N__33313),
            .I(\c0.FRAME_MATCHER_state_8 ));
    SRMux I__6988 (
            .O(N__33306),
            .I(N__33303));
    LocalMux I__6987 (
            .O(N__33303),
            .I(N__33300));
    Span4Mux_v I__6986 (
            .O(N__33300),
            .I(N__33297));
    Span4Mux_h I__6985 (
            .O(N__33297),
            .I(N__33294));
    Odrv4 I__6984 (
            .O(N__33294),
            .I(\c0.n16666 ));
    InMux I__6983 (
            .O(N__33291),
            .I(N__33287));
    CascadeMux I__6982 (
            .O(N__33290),
            .I(N__33284));
    LocalMux I__6981 (
            .O(N__33287),
            .I(N__33281));
    InMux I__6980 (
            .O(N__33284),
            .I(N__33277));
    Span4Mux_v I__6979 (
            .O(N__33281),
            .I(N__33274));
    InMux I__6978 (
            .O(N__33280),
            .I(N__33271));
    LocalMux I__6977 (
            .O(N__33277),
            .I(\c0.FRAME_MATCHER_state_9 ));
    Odrv4 I__6976 (
            .O(N__33274),
            .I(\c0.FRAME_MATCHER_state_9 ));
    LocalMux I__6975 (
            .O(N__33271),
            .I(\c0.FRAME_MATCHER_state_9 ));
    SRMux I__6974 (
            .O(N__33264),
            .I(N__33261));
    LocalMux I__6973 (
            .O(N__33261),
            .I(N__33258));
    Span4Mux_h I__6972 (
            .O(N__33258),
            .I(N__33255));
    Odrv4 I__6971 (
            .O(N__33255),
            .I(\c0.n16674 ));
    InMux I__6970 (
            .O(N__33252),
            .I(N__33243));
    InMux I__6969 (
            .O(N__33251),
            .I(N__33240));
    InMux I__6968 (
            .O(N__33250),
            .I(N__33237));
    InMux I__6967 (
            .O(N__33249),
            .I(N__33229));
    InMux I__6966 (
            .O(N__33248),
            .I(N__33226));
    InMux I__6965 (
            .O(N__33247),
            .I(N__33215));
    InMux I__6964 (
            .O(N__33246),
            .I(N__33212));
    LocalMux I__6963 (
            .O(N__33243),
            .I(N__33207));
    LocalMux I__6962 (
            .O(N__33240),
            .I(N__33207));
    LocalMux I__6961 (
            .O(N__33237),
            .I(N__33204));
    InMux I__6960 (
            .O(N__33236),
            .I(N__33201));
    InMux I__6959 (
            .O(N__33235),
            .I(N__33198));
    InMux I__6958 (
            .O(N__33234),
            .I(N__33194));
    InMux I__6957 (
            .O(N__33233),
            .I(N__33191));
    InMux I__6956 (
            .O(N__33232),
            .I(N__33188));
    LocalMux I__6955 (
            .O(N__33229),
            .I(N__33179));
    LocalMux I__6954 (
            .O(N__33226),
            .I(N__33179));
    InMux I__6953 (
            .O(N__33225),
            .I(N__33176));
    InMux I__6952 (
            .O(N__33224),
            .I(N__33173));
    InMux I__6951 (
            .O(N__33223),
            .I(N__33170));
    InMux I__6950 (
            .O(N__33222),
            .I(N__33167));
    InMux I__6949 (
            .O(N__33221),
            .I(N__33164));
    InMux I__6948 (
            .O(N__33220),
            .I(N__33161));
    InMux I__6947 (
            .O(N__33219),
            .I(N__33156));
    InMux I__6946 (
            .O(N__33218),
            .I(N__33153));
    LocalMux I__6945 (
            .O(N__33215),
            .I(N__33143));
    LocalMux I__6944 (
            .O(N__33212),
            .I(N__33143));
    Span4Mux_h I__6943 (
            .O(N__33207),
            .I(N__33134));
    Span4Mux_s2_v I__6942 (
            .O(N__33204),
            .I(N__33134));
    LocalMux I__6941 (
            .O(N__33201),
            .I(N__33134));
    LocalMux I__6940 (
            .O(N__33198),
            .I(N__33134));
    InMux I__6939 (
            .O(N__33197),
            .I(N__33131));
    LocalMux I__6938 (
            .O(N__33194),
            .I(N__33124));
    LocalMux I__6937 (
            .O(N__33191),
            .I(N__33124));
    LocalMux I__6936 (
            .O(N__33188),
            .I(N__33124));
    InMux I__6935 (
            .O(N__33187),
            .I(N__33121));
    InMux I__6934 (
            .O(N__33186),
            .I(N__33118));
    InMux I__6933 (
            .O(N__33185),
            .I(N__33115));
    InMux I__6932 (
            .O(N__33184),
            .I(N__33112));
    Span4Mux_s3_v I__6931 (
            .O(N__33179),
            .I(N__33099));
    LocalMux I__6930 (
            .O(N__33176),
            .I(N__33099));
    LocalMux I__6929 (
            .O(N__33173),
            .I(N__33099));
    LocalMux I__6928 (
            .O(N__33170),
            .I(N__33099));
    LocalMux I__6927 (
            .O(N__33167),
            .I(N__33099));
    LocalMux I__6926 (
            .O(N__33164),
            .I(N__33099));
    LocalMux I__6925 (
            .O(N__33161),
            .I(N__33096));
    InMux I__6924 (
            .O(N__33160),
            .I(N__33093));
    InMux I__6923 (
            .O(N__33159),
            .I(N__33090));
    LocalMux I__6922 (
            .O(N__33156),
            .I(N__33085));
    LocalMux I__6921 (
            .O(N__33153),
            .I(N__33085));
    InMux I__6920 (
            .O(N__33152),
            .I(N__33082));
    InMux I__6919 (
            .O(N__33151),
            .I(N__33079));
    InMux I__6918 (
            .O(N__33150),
            .I(N__33076));
    InMux I__6917 (
            .O(N__33149),
            .I(N__33073));
    InMux I__6916 (
            .O(N__33148),
            .I(N__33070));
    Span4Mux_h I__6915 (
            .O(N__33143),
            .I(N__33063));
    Span4Mux_v I__6914 (
            .O(N__33134),
            .I(N__33063));
    LocalMux I__6913 (
            .O(N__33131),
            .I(N__33063));
    Span4Mux_s3_v I__6912 (
            .O(N__33124),
            .I(N__33052));
    LocalMux I__6911 (
            .O(N__33121),
            .I(N__33052));
    LocalMux I__6910 (
            .O(N__33118),
            .I(N__33052));
    LocalMux I__6909 (
            .O(N__33115),
            .I(N__33052));
    LocalMux I__6908 (
            .O(N__33112),
            .I(N__33052));
    Span4Mux_v I__6907 (
            .O(N__33099),
            .I(N__33045));
    Span4Mux_s2_h I__6906 (
            .O(N__33096),
            .I(N__33045));
    LocalMux I__6905 (
            .O(N__33093),
            .I(N__33045));
    LocalMux I__6904 (
            .O(N__33090),
            .I(N__33040));
    Span4Mux_h I__6903 (
            .O(N__33085),
            .I(N__33040));
    LocalMux I__6902 (
            .O(N__33082),
            .I(N__33028));
    LocalMux I__6901 (
            .O(N__33079),
            .I(N__33028));
    LocalMux I__6900 (
            .O(N__33076),
            .I(N__33028));
    LocalMux I__6899 (
            .O(N__33073),
            .I(N__33028));
    LocalMux I__6898 (
            .O(N__33070),
            .I(N__33028));
    Span4Mux_v I__6897 (
            .O(N__33063),
            .I(N__33025));
    Span4Mux_v I__6896 (
            .O(N__33052),
            .I(N__33020));
    Span4Mux_h I__6895 (
            .O(N__33045),
            .I(N__33020));
    Span4Mux_h I__6894 (
            .O(N__33040),
            .I(N__33017));
    InMux I__6893 (
            .O(N__33039),
            .I(N__33014));
    Span12Mux_s10_v I__6892 (
            .O(N__33028),
            .I(N__33008));
    Span4Mux_h I__6891 (
            .O(N__33025),
            .I(N__33005));
    Span4Mux_h I__6890 (
            .O(N__33020),
            .I(N__33002));
    Span4Mux_v I__6889 (
            .O(N__33017),
            .I(N__32999));
    LocalMux I__6888 (
            .O(N__33014),
            .I(N__32996));
    InMux I__6887 (
            .O(N__33013),
            .I(N__32993));
    InMux I__6886 (
            .O(N__33012),
            .I(N__32990));
    InMux I__6885 (
            .O(N__33011),
            .I(N__32987));
    Odrv12 I__6884 (
            .O(N__33008),
            .I(\c0.n1034 ));
    Odrv4 I__6883 (
            .O(N__33005),
            .I(\c0.n1034 ));
    Odrv4 I__6882 (
            .O(N__33002),
            .I(\c0.n1034 ));
    Odrv4 I__6881 (
            .O(N__32999),
            .I(\c0.n1034 ));
    Odrv12 I__6880 (
            .O(N__32996),
            .I(\c0.n1034 ));
    LocalMux I__6879 (
            .O(N__32993),
            .I(\c0.n1034 ));
    LocalMux I__6878 (
            .O(N__32990),
            .I(\c0.n1034 ));
    LocalMux I__6877 (
            .O(N__32987),
            .I(\c0.n1034 ));
    CascadeMux I__6876 (
            .O(N__32970),
            .I(n10140_cascade_));
    CascadeMux I__6875 (
            .O(N__32967),
            .I(\c0.n23_cascade_ ));
    InMux I__6874 (
            .O(N__32964),
            .I(N__32961));
    LocalMux I__6873 (
            .O(N__32961),
            .I(\c0.n26_adj_2210 ));
    InMux I__6872 (
            .O(N__32958),
            .I(N__32955));
    LocalMux I__6871 (
            .O(N__32955),
            .I(\c0.n18 ));
    CascadeMux I__6870 (
            .O(N__32952),
            .I(\c0.n30_adj_2213_cascade_ ));
    InMux I__6869 (
            .O(N__32949),
            .I(N__32946));
    LocalMux I__6868 (
            .O(N__32946),
            .I(N__32943));
    Odrv4 I__6867 (
            .O(N__32943),
            .I(\c0.n17_adj_2214 ));
    CascadeMux I__6866 (
            .O(N__32940),
            .I(n31_adj_2415_cascade_));
    InMux I__6865 (
            .O(N__32937),
            .I(N__32933));
    InMux I__6864 (
            .O(N__32936),
            .I(N__32930));
    LocalMux I__6863 (
            .O(N__32933),
            .I(N__32927));
    LocalMux I__6862 (
            .O(N__32930),
            .I(data_in_frame_6_3));
    Odrv4 I__6861 (
            .O(N__32927),
            .I(data_in_frame_6_3));
    InMux I__6860 (
            .O(N__32922),
            .I(N__32917));
    InMux I__6859 (
            .O(N__32921),
            .I(N__32911));
    InMux I__6858 (
            .O(N__32920),
            .I(N__32911));
    LocalMux I__6857 (
            .O(N__32917),
            .I(N__32908));
    InMux I__6856 (
            .O(N__32916),
            .I(N__32905));
    LocalMux I__6855 (
            .O(N__32911),
            .I(data_in_3_7));
    Odrv4 I__6854 (
            .O(N__32908),
            .I(data_in_3_7));
    LocalMux I__6853 (
            .O(N__32905),
            .I(data_in_3_7));
    InMux I__6852 (
            .O(N__32898),
            .I(N__32895));
    LocalMux I__6851 (
            .O(N__32895),
            .I(\c0.n6_adj_2358 ));
    InMux I__6850 (
            .O(N__32892),
            .I(N__32889));
    LocalMux I__6849 (
            .O(N__32889),
            .I(N__32885));
    InMux I__6848 (
            .O(N__32888),
            .I(N__32881));
    Span4Mux_v I__6847 (
            .O(N__32885),
            .I(N__32877));
    CascadeMux I__6846 (
            .O(N__32884),
            .I(N__32874));
    LocalMux I__6845 (
            .O(N__32881),
            .I(N__32869));
    InMux I__6844 (
            .O(N__32880),
            .I(N__32866));
    Span4Mux_v I__6843 (
            .O(N__32877),
            .I(N__32862));
    InMux I__6842 (
            .O(N__32874),
            .I(N__32857));
    InMux I__6841 (
            .O(N__32873),
            .I(N__32857));
    CascadeMux I__6840 (
            .O(N__32872),
            .I(N__32854));
    Span4Mux_h I__6839 (
            .O(N__32869),
            .I(N__32849));
    LocalMux I__6838 (
            .O(N__32866),
            .I(N__32849));
    InMux I__6837 (
            .O(N__32865),
            .I(N__32846));
    Span4Mux_h I__6836 (
            .O(N__32862),
            .I(N__32841));
    LocalMux I__6835 (
            .O(N__32857),
            .I(N__32841));
    InMux I__6834 (
            .O(N__32854),
            .I(N__32838));
    Span4Mux_v I__6833 (
            .O(N__32849),
            .I(N__32833));
    LocalMux I__6832 (
            .O(N__32846),
            .I(N__32833));
    Span4Mux_v I__6831 (
            .O(N__32841),
            .I(N__32830));
    LocalMux I__6830 (
            .O(N__32838),
            .I(N__32827));
    Span4Mux_h I__6829 (
            .O(N__32833),
            .I(N__32824));
    Span4Mux_h I__6828 (
            .O(N__32830),
            .I(N__32819));
    Span4Mux_v I__6827 (
            .O(N__32827),
            .I(N__32819));
    Span4Mux_h I__6826 (
            .O(N__32824),
            .I(N__32816));
    Odrv4 I__6825 (
            .O(N__32819),
            .I(\c0.FRAME_MATCHER_i_1 ));
    Odrv4 I__6824 (
            .O(N__32816),
            .I(\c0.FRAME_MATCHER_i_1 ));
    CascadeMux I__6823 (
            .O(N__32811),
            .I(N__32807));
    InMux I__6822 (
            .O(N__32810),
            .I(N__32804));
    InMux I__6821 (
            .O(N__32807),
            .I(N__32801));
    LocalMux I__6820 (
            .O(N__32804),
            .I(N__32798));
    LocalMux I__6819 (
            .O(N__32801),
            .I(N__32795));
    Span4Mux_v I__6818 (
            .O(N__32798),
            .I(N__32792));
    Span4Mux_h I__6817 (
            .O(N__32795),
            .I(N__32788));
    Span4Mux_v I__6816 (
            .O(N__32792),
            .I(N__32785));
    InMux I__6815 (
            .O(N__32791),
            .I(N__32782));
    Span4Mux_h I__6814 (
            .O(N__32788),
            .I(N__32779));
    Span4Mux_h I__6813 (
            .O(N__32785),
            .I(N__32774));
    LocalMux I__6812 (
            .O(N__32782),
            .I(N__32774));
    Odrv4 I__6811 (
            .O(N__32779),
            .I(\c0.n15164 ));
    Odrv4 I__6810 (
            .O(N__32774),
            .I(\c0.n15164 ));
    CascadeMux I__6809 (
            .O(N__32769),
            .I(\c0.n17072_cascade_ ));
    InMux I__6808 (
            .O(N__32766),
            .I(N__32762));
    InMux I__6807 (
            .O(N__32765),
            .I(N__32759));
    LocalMux I__6806 (
            .O(N__32762),
            .I(N__32756));
    LocalMux I__6805 (
            .O(N__32759),
            .I(\c0.n10215 ));
    Odrv4 I__6804 (
            .O(N__32756),
            .I(\c0.n10215 ));
    InMux I__6803 (
            .O(N__32751),
            .I(N__32746));
    InMux I__6802 (
            .O(N__32750),
            .I(N__32742));
    InMux I__6801 (
            .O(N__32749),
            .I(N__32739));
    LocalMux I__6800 (
            .O(N__32746),
            .I(N__32736));
    InMux I__6799 (
            .O(N__32745),
            .I(N__32733));
    LocalMux I__6798 (
            .O(N__32742),
            .I(\c0.data_in_frame_0_4 ));
    LocalMux I__6797 (
            .O(N__32739),
            .I(\c0.data_in_frame_0_4 ));
    Odrv4 I__6796 (
            .O(N__32736),
            .I(\c0.data_in_frame_0_4 ));
    LocalMux I__6795 (
            .O(N__32733),
            .I(\c0.data_in_frame_0_4 ));
    CascadeMux I__6794 (
            .O(N__32724),
            .I(\c0.n10215_cascade_ ));
    CascadeMux I__6793 (
            .O(N__32721),
            .I(\c0.n17206_cascade_ ));
    InMux I__6792 (
            .O(N__32718),
            .I(N__32715));
    LocalMux I__6791 (
            .O(N__32715),
            .I(N__32712));
    Odrv4 I__6790 (
            .O(N__32712),
            .I(\c0.n20_adj_2195 ));
    CascadeMux I__6789 (
            .O(N__32709),
            .I(N__32703));
    InMux I__6788 (
            .O(N__32708),
            .I(N__32697));
    InMux I__6787 (
            .O(N__32707),
            .I(N__32697));
    InMux I__6786 (
            .O(N__32706),
            .I(N__32692));
    InMux I__6785 (
            .O(N__32703),
            .I(N__32687));
    InMux I__6784 (
            .O(N__32702),
            .I(N__32687));
    LocalMux I__6783 (
            .O(N__32697),
            .I(N__32684));
    CascadeMux I__6782 (
            .O(N__32696),
            .I(N__32681));
    CascadeMux I__6781 (
            .O(N__32695),
            .I(N__32677));
    LocalMux I__6780 (
            .O(N__32692),
            .I(N__32674));
    LocalMux I__6779 (
            .O(N__32687),
            .I(N__32671));
    Span4Mux_h I__6778 (
            .O(N__32684),
            .I(N__32668));
    InMux I__6777 (
            .O(N__32681),
            .I(N__32665));
    InMux I__6776 (
            .O(N__32680),
            .I(N__32660));
    InMux I__6775 (
            .O(N__32677),
            .I(N__32660));
    Span4Mux_v I__6774 (
            .O(N__32674),
            .I(N__32655));
    Span4Mux_v I__6773 (
            .O(N__32671),
            .I(N__32655));
    Span4Mux_h I__6772 (
            .O(N__32668),
            .I(N__32652));
    LocalMux I__6771 (
            .O(N__32665),
            .I(N__32647));
    LocalMux I__6770 (
            .O(N__32660),
            .I(N__32647));
    Span4Mux_v I__6769 (
            .O(N__32655),
            .I(N__32644));
    Span4Mux_v I__6768 (
            .O(N__32652),
            .I(N__32641));
    Span12Mux_h I__6767 (
            .O(N__32647),
            .I(N__32637));
    Span4Mux_h I__6766 (
            .O(N__32644),
            .I(N__32634));
    Span4Mux_v I__6765 (
            .O(N__32641),
            .I(N__32631));
    InMux I__6764 (
            .O(N__32640),
            .I(N__32628));
    Odrv12 I__6763 (
            .O(N__32637),
            .I(\c0.n39 ));
    Odrv4 I__6762 (
            .O(N__32634),
            .I(\c0.n39 ));
    Odrv4 I__6761 (
            .O(N__32631),
            .I(\c0.n39 ));
    LocalMux I__6760 (
            .O(N__32628),
            .I(\c0.n39 ));
    InMux I__6759 (
            .O(N__32619),
            .I(N__32615));
    InMux I__6758 (
            .O(N__32618),
            .I(N__32612));
    LocalMux I__6757 (
            .O(N__32615),
            .I(\c0.n2137 ));
    LocalMux I__6756 (
            .O(N__32612),
            .I(\c0.n2137 ));
    InMux I__6755 (
            .O(N__32607),
            .I(N__32604));
    LocalMux I__6754 (
            .O(N__32604),
            .I(\c0.n16475 ));
    InMux I__6753 (
            .O(N__32601),
            .I(N__32597));
    InMux I__6752 (
            .O(N__32600),
            .I(N__32594));
    LocalMux I__6751 (
            .O(N__32597),
            .I(\c0.data_in_frame_5_5 ));
    LocalMux I__6750 (
            .O(N__32594),
            .I(\c0.data_in_frame_5_5 ));
    CascadeMux I__6749 (
            .O(N__32589),
            .I(N__32586));
    InMux I__6748 (
            .O(N__32586),
            .I(N__32583));
    LocalMux I__6747 (
            .O(N__32583),
            .I(N__32580));
    Span4Mux_v I__6746 (
            .O(N__32580),
            .I(N__32577));
    Odrv4 I__6745 (
            .O(N__32577),
            .I(\c0.n17373 ));
    InMux I__6744 (
            .O(N__32574),
            .I(N__32571));
    LocalMux I__6743 (
            .O(N__32571),
            .I(\c0.n19_adj_2303 ));
    CascadeMux I__6742 (
            .O(N__32568),
            .I(\c0.n17076_cascade_ ));
    InMux I__6741 (
            .O(N__32565),
            .I(N__32556));
    InMux I__6740 (
            .O(N__32564),
            .I(N__32553));
    InMux I__6739 (
            .O(N__32563),
            .I(N__32546));
    InMux I__6738 (
            .O(N__32562),
            .I(N__32546));
    InMux I__6737 (
            .O(N__32561),
            .I(N__32546));
    InMux I__6736 (
            .O(N__32560),
            .I(N__32541));
    InMux I__6735 (
            .O(N__32559),
            .I(N__32541));
    LocalMux I__6734 (
            .O(N__32556),
            .I(n17075));
    LocalMux I__6733 (
            .O(N__32553),
            .I(n17075));
    LocalMux I__6732 (
            .O(N__32546),
            .I(n17075));
    LocalMux I__6731 (
            .O(N__32541),
            .I(n17075));
    CascadeMux I__6730 (
            .O(N__32532),
            .I(N__32528));
    InMux I__6729 (
            .O(N__32531),
            .I(N__32525));
    InMux I__6728 (
            .O(N__32528),
            .I(N__32522));
    LocalMux I__6727 (
            .O(N__32525),
            .I(data_in_frame_6_4));
    LocalMux I__6726 (
            .O(N__32522),
            .I(data_in_frame_6_4));
    CascadeMux I__6725 (
            .O(N__32517),
            .I(\c0.n2122_cascade_ ));
    InMux I__6724 (
            .O(N__32514),
            .I(N__32511));
    LocalMux I__6723 (
            .O(N__32511),
            .I(N__32508));
    Span4Mux_h I__6722 (
            .O(N__32508),
            .I(N__32503));
    InMux I__6721 (
            .O(N__32507),
            .I(N__32498));
    InMux I__6720 (
            .O(N__32506),
            .I(N__32498));
    Odrv4 I__6719 (
            .O(N__32503),
            .I(\c0.data_in_frame_2_5 ));
    LocalMux I__6718 (
            .O(N__32498),
            .I(\c0.data_in_frame_2_5 ));
    CascadeMux I__6717 (
            .O(N__32493),
            .I(N__32489));
    InMux I__6716 (
            .O(N__32492),
            .I(N__32486));
    InMux I__6715 (
            .O(N__32489),
            .I(N__32483));
    LocalMux I__6714 (
            .O(N__32486),
            .I(\c0.data_in_frame_5_6 ));
    LocalMux I__6713 (
            .O(N__32483),
            .I(\c0.data_in_frame_5_6 ));
    CascadeMux I__6712 (
            .O(N__32478),
            .I(\c0.n2124_cascade_ ));
    InMux I__6711 (
            .O(N__32475),
            .I(N__32471));
    InMux I__6710 (
            .O(N__32474),
            .I(N__32468));
    LocalMux I__6709 (
            .O(N__32471),
            .I(\c0.data_in_frame_5_3 ));
    LocalMux I__6708 (
            .O(N__32468),
            .I(\c0.data_in_frame_5_3 ));
    InMux I__6707 (
            .O(N__32463),
            .I(N__32455));
    InMux I__6706 (
            .O(N__32462),
            .I(N__32448));
    InMux I__6705 (
            .O(N__32461),
            .I(N__32448));
    InMux I__6704 (
            .O(N__32460),
            .I(N__32448));
    InMux I__6703 (
            .O(N__32459),
            .I(N__32436));
    InMux I__6702 (
            .O(N__32458),
            .I(N__32436));
    LocalMux I__6701 (
            .O(N__32455),
            .I(N__32433));
    LocalMux I__6700 (
            .O(N__32448),
            .I(N__32430));
    InMux I__6699 (
            .O(N__32447),
            .I(N__32425));
    InMux I__6698 (
            .O(N__32446),
            .I(N__32425));
    InMux I__6697 (
            .O(N__32445),
            .I(N__32418));
    InMux I__6696 (
            .O(N__32444),
            .I(N__32418));
    InMux I__6695 (
            .O(N__32443),
            .I(N__32405));
    InMux I__6694 (
            .O(N__32442),
            .I(N__32405));
    InMux I__6693 (
            .O(N__32441),
            .I(N__32405));
    LocalMux I__6692 (
            .O(N__32436),
            .I(N__32402));
    Span4Mux_s1_h I__6691 (
            .O(N__32433),
            .I(N__32395));
    Span4Mux_v I__6690 (
            .O(N__32430),
            .I(N__32395));
    LocalMux I__6689 (
            .O(N__32425),
            .I(N__32395));
    InMux I__6688 (
            .O(N__32424),
            .I(N__32392));
    InMux I__6687 (
            .O(N__32423),
            .I(N__32389));
    LocalMux I__6686 (
            .O(N__32418),
            .I(N__32385));
    InMux I__6685 (
            .O(N__32417),
            .I(N__32378));
    InMux I__6684 (
            .O(N__32416),
            .I(N__32378));
    InMux I__6683 (
            .O(N__32415),
            .I(N__32378));
    InMux I__6682 (
            .O(N__32414),
            .I(N__32371));
    InMux I__6681 (
            .O(N__32413),
            .I(N__32371));
    InMux I__6680 (
            .O(N__32412),
            .I(N__32371));
    LocalMux I__6679 (
            .O(N__32405),
            .I(N__32364));
    Span4Mux_s1_h I__6678 (
            .O(N__32402),
            .I(N__32364));
    Span4Mux_h I__6677 (
            .O(N__32395),
            .I(N__32359));
    LocalMux I__6676 (
            .O(N__32392),
            .I(N__32354));
    LocalMux I__6675 (
            .O(N__32389),
            .I(N__32354));
    InMux I__6674 (
            .O(N__32388),
            .I(N__32351));
    Span4Mux_v I__6673 (
            .O(N__32385),
            .I(N__32348));
    LocalMux I__6672 (
            .O(N__32378),
            .I(N__32343));
    LocalMux I__6671 (
            .O(N__32371),
            .I(N__32343));
    InMux I__6670 (
            .O(N__32370),
            .I(N__32338));
    InMux I__6669 (
            .O(N__32369),
            .I(N__32338));
    Span4Mux_h I__6668 (
            .O(N__32364),
            .I(N__32335));
    InMux I__6667 (
            .O(N__32363),
            .I(N__32330));
    InMux I__6666 (
            .O(N__32362),
            .I(N__32327));
    Span4Mux_h I__6665 (
            .O(N__32359),
            .I(N__32324));
    Span12Mux_s5_h I__6664 (
            .O(N__32354),
            .I(N__32313));
    LocalMux I__6663 (
            .O(N__32351),
            .I(N__32313));
    Sp12to4 I__6662 (
            .O(N__32348),
            .I(N__32313));
    Span12Mux_v I__6661 (
            .O(N__32343),
            .I(N__32313));
    LocalMux I__6660 (
            .O(N__32338),
            .I(N__32313));
    Span4Mux_h I__6659 (
            .O(N__32335),
            .I(N__32310));
    InMux I__6658 (
            .O(N__32334),
            .I(N__32307));
    InMux I__6657 (
            .O(N__32333),
            .I(N__32304));
    LocalMux I__6656 (
            .O(N__32330),
            .I(\c0.byte_transmit_counter2_3 ));
    LocalMux I__6655 (
            .O(N__32327),
            .I(\c0.byte_transmit_counter2_3 ));
    Odrv4 I__6654 (
            .O(N__32324),
            .I(\c0.byte_transmit_counter2_3 ));
    Odrv12 I__6653 (
            .O(N__32313),
            .I(\c0.byte_transmit_counter2_3 ));
    Odrv4 I__6652 (
            .O(N__32310),
            .I(\c0.byte_transmit_counter2_3 ));
    LocalMux I__6651 (
            .O(N__32307),
            .I(\c0.byte_transmit_counter2_3 ));
    LocalMux I__6650 (
            .O(N__32304),
            .I(\c0.byte_transmit_counter2_3 ));
    InMux I__6649 (
            .O(N__32289),
            .I(N__32284));
    InMux I__6648 (
            .O(N__32288),
            .I(N__32281));
    InMux I__6647 (
            .O(N__32287),
            .I(N__32278));
    LocalMux I__6646 (
            .O(N__32284),
            .I(N__32268));
    LocalMux I__6645 (
            .O(N__32281),
            .I(N__32268));
    LocalMux I__6644 (
            .O(N__32278),
            .I(N__32268));
    InMux I__6643 (
            .O(N__32277),
            .I(N__32265));
    CascadeMux I__6642 (
            .O(N__32276),
            .I(N__32262));
    InMux I__6641 (
            .O(N__32275),
            .I(N__32257));
    Span4Mux_v I__6640 (
            .O(N__32268),
            .I(N__32254));
    LocalMux I__6639 (
            .O(N__32265),
            .I(N__32251));
    InMux I__6638 (
            .O(N__32262),
            .I(N__32248));
    InMux I__6637 (
            .O(N__32261),
            .I(N__32244));
    InMux I__6636 (
            .O(N__32260),
            .I(N__32241));
    LocalMux I__6635 (
            .O(N__32257),
            .I(N__32236));
    IoSpan4Mux I__6634 (
            .O(N__32254),
            .I(N__32236));
    Span4Mux_v I__6633 (
            .O(N__32251),
            .I(N__32229));
    LocalMux I__6632 (
            .O(N__32248),
            .I(N__32229));
    InMux I__6631 (
            .O(N__32247),
            .I(N__32226));
    LocalMux I__6630 (
            .O(N__32244),
            .I(N__32218));
    LocalMux I__6629 (
            .O(N__32241),
            .I(N__32218));
    Span4Mux_s3_h I__6628 (
            .O(N__32236),
            .I(N__32218));
    InMux I__6627 (
            .O(N__32235),
            .I(N__32215));
    InMux I__6626 (
            .O(N__32234),
            .I(N__32212));
    Span4Mux_h I__6625 (
            .O(N__32229),
            .I(N__32209));
    LocalMux I__6624 (
            .O(N__32226),
            .I(N__32206));
    InMux I__6623 (
            .O(N__32225),
            .I(N__32203));
    Span4Mux_h I__6622 (
            .O(N__32218),
            .I(N__32198));
    LocalMux I__6621 (
            .O(N__32215),
            .I(N__32198));
    LocalMux I__6620 (
            .O(N__32212),
            .I(\c0.byte_transmit_counter2_4 ));
    Odrv4 I__6619 (
            .O(N__32209),
            .I(\c0.byte_transmit_counter2_4 ));
    Odrv12 I__6618 (
            .O(N__32206),
            .I(\c0.byte_transmit_counter2_4 ));
    LocalMux I__6617 (
            .O(N__32203),
            .I(\c0.byte_transmit_counter2_4 ));
    Odrv4 I__6616 (
            .O(N__32198),
            .I(\c0.byte_transmit_counter2_4 ));
    InMux I__6615 (
            .O(N__32187),
            .I(N__32184));
    LocalMux I__6614 (
            .O(N__32184),
            .I(N__32181));
    Span4Mux_h I__6613 (
            .O(N__32181),
            .I(N__32178));
    Odrv4 I__6612 (
            .O(N__32178),
            .I(\c0.n17710 ));
    InMux I__6611 (
            .O(N__32175),
            .I(N__32162));
    InMux I__6610 (
            .O(N__32174),
            .I(N__32162));
    InMux I__6609 (
            .O(N__32173),
            .I(N__32157));
    InMux I__6608 (
            .O(N__32172),
            .I(N__32157));
    InMux I__6607 (
            .O(N__32171),
            .I(N__32154));
    CascadeMux I__6606 (
            .O(N__32170),
            .I(N__32150));
    InMux I__6605 (
            .O(N__32169),
            .I(N__32143));
    InMux I__6604 (
            .O(N__32168),
            .I(N__32136));
    InMux I__6603 (
            .O(N__32167),
            .I(N__32136));
    LocalMux I__6602 (
            .O(N__32162),
            .I(N__32133));
    LocalMux I__6601 (
            .O(N__32157),
            .I(N__32128));
    LocalMux I__6600 (
            .O(N__32154),
            .I(N__32128));
    InMux I__6599 (
            .O(N__32153),
            .I(N__32123));
    InMux I__6598 (
            .O(N__32150),
            .I(N__32123));
    InMux I__6597 (
            .O(N__32149),
            .I(N__32120));
    InMux I__6596 (
            .O(N__32148),
            .I(N__32113));
    InMux I__6595 (
            .O(N__32147),
            .I(N__32113));
    InMux I__6594 (
            .O(N__32146),
            .I(N__32113));
    LocalMux I__6593 (
            .O(N__32143),
            .I(N__32110));
    InMux I__6592 (
            .O(N__32142),
            .I(N__32104));
    InMux I__6591 (
            .O(N__32141),
            .I(N__32104));
    LocalMux I__6590 (
            .O(N__32136),
            .I(N__32101));
    Span4Mux_v I__6589 (
            .O(N__32133),
            .I(N__32096));
    Span4Mux_v I__6588 (
            .O(N__32128),
            .I(N__32096));
    LocalMux I__6587 (
            .O(N__32123),
            .I(N__32087));
    LocalMux I__6586 (
            .O(N__32120),
            .I(N__32087));
    LocalMux I__6585 (
            .O(N__32113),
            .I(N__32087));
    Span4Mux_v I__6584 (
            .O(N__32110),
            .I(N__32087));
    InMux I__6583 (
            .O(N__32109),
            .I(N__32084));
    LocalMux I__6582 (
            .O(N__32104),
            .I(N__32077));
    Span4Mux_v I__6581 (
            .O(N__32101),
            .I(N__32077));
    Span4Mux_h I__6580 (
            .O(N__32096),
            .I(N__32077));
    Span4Mux_h I__6579 (
            .O(N__32087),
            .I(N__32072));
    LocalMux I__6578 (
            .O(N__32084),
            .I(N__32072));
    Span4Mux_h I__6577 (
            .O(N__32077),
            .I(N__32066));
    Span4Mux_h I__6576 (
            .O(N__32072),
            .I(N__32063));
    InMux I__6575 (
            .O(N__32071),
            .I(N__32056));
    InMux I__6574 (
            .O(N__32070),
            .I(N__32056));
    InMux I__6573 (
            .O(N__32069),
            .I(N__32056));
    Odrv4 I__6572 (
            .O(N__32066),
            .I(\c0.byte_transmit_counter2_2 ));
    Odrv4 I__6571 (
            .O(N__32063),
            .I(\c0.byte_transmit_counter2_2 ));
    LocalMux I__6570 (
            .O(N__32056),
            .I(\c0.byte_transmit_counter2_2 ));
    SRMux I__6569 (
            .O(N__32049),
            .I(N__32046));
    LocalMux I__6568 (
            .O(N__32046),
            .I(\c0.n4_adj_2154 ));
    SRMux I__6567 (
            .O(N__32043),
            .I(N__32040));
    LocalMux I__6566 (
            .O(N__32040),
            .I(N__32037));
    Span4Mux_h I__6565 (
            .O(N__32037),
            .I(N__32034));
    Odrv4 I__6564 (
            .O(N__32034),
            .I(\c0.n4_adj_2345 ));
    CascadeMux I__6563 (
            .O(N__32031),
            .I(N__32027));
    InMux I__6562 (
            .O(N__32030),
            .I(N__32024));
    InMux I__6561 (
            .O(N__32027),
            .I(N__32021));
    LocalMux I__6560 (
            .O(N__32024),
            .I(rand_setpoint_28));
    LocalMux I__6559 (
            .O(N__32021),
            .I(rand_setpoint_28));
    InMux I__6558 (
            .O(N__32016),
            .I(N__32013));
    LocalMux I__6557 (
            .O(N__32013),
            .I(N__32009));
    CascadeMux I__6556 (
            .O(N__32012),
            .I(N__32006));
    Span12Mux_s3_v I__6555 (
            .O(N__32009),
            .I(N__32003));
    InMux I__6554 (
            .O(N__32006),
            .I(N__32000));
    Odrv12 I__6553 (
            .O(N__32003),
            .I(rand_setpoint_11));
    LocalMux I__6552 (
            .O(N__32000),
            .I(rand_setpoint_11));
    CascadeMux I__6551 (
            .O(N__31995),
            .I(N__31992));
    InMux I__6550 (
            .O(N__31992),
            .I(N__31989));
    LocalMux I__6549 (
            .O(N__31989),
            .I(N__31986));
    Span4Mux_s2_v I__6548 (
            .O(N__31986),
            .I(N__31983));
    Span4Mux_h I__6547 (
            .O(N__31983),
            .I(N__31980));
    Odrv4 I__6546 (
            .O(N__31980),
            .I(\c0.n17585 ));
    InMux I__6545 (
            .O(N__31977),
            .I(N__31974));
    LocalMux I__6544 (
            .O(N__31974),
            .I(N__31970));
    CascadeMux I__6543 (
            .O(N__31973),
            .I(N__31967));
    Span4Mux_s3_v I__6542 (
            .O(N__31970),
            .I(N__31964));
    InMux I__6541 (
            .O(N__31967),
            .I(N__31961));
    Odrv4 I__6540 (
            .O(N__31964),
            .I(rand_setpoint_10));
    LocalMux I__6539 (
            .O(N__31961),
            .I(rand_setpoint_10));
    CascadeMux I__6538 (
            .O(N__31956),
            .I(\c0.n17583_cascade_ ));
    InMux I__6537 (
            .O(N__31953),
            .I(N__31949));
    CascadeMux I__6536 (
            .O(N__31952),
            .I(N__31946));
    LocalMux I__6535 (
            .O(N__31949),
            .I(N__31943));
    InMux I__6534 (
            .O(N__31946),
            .I(N__31940));
    Span4Mux_h I__6533 (
            .O(N__31943),
            .I(N__31934));
    LocalMux I__6532 (
            .O(N__31940),
            .I(N__31930));
    InMux I__6531 (
            .O(N__31939),
            .I(N__31927));
    InMux I__6530 (
            .O(N__31938),
            .I(N__31922));
    InMux I__6529 (
            .O(N__31937),
            .I(N__31922));
    Span4Mux_h I__6528 (
            .O(N__31934),
            .I(N__31919));
    InMux I__6527 (
            .O(N__31933),
            .I(N__31916));
    Span4Mux_h I__6526 (
            .O(N__31930),
            .I(N__31913));
    LocalMux I__6525 (
            .O(N__31927),
            .I(N__31908));
    LocalMux I__6524 (
            .O(N__31922),
            .I(N__31908));
    Odrv4 I__6523 (
            .O(N__31919),
            .I(\c0.rx.r_Clock_Count_5 ));
    LocalMux I__6522 (
            .O(N__31916),
            .I(\c0.rx.r_Clock_Count_5 ));
    Odrv4 I__6521 (
            .O(N__31913),
            .I(\c0.rx.r_Clock_Count_5 ));
    Odrv12 I__6520 (
            .O(N__31908),
            .I(\c0.rx.r_Clock_Count_5 ));
    InMux I__6519 (
            .O(N__31899),
            .I(N__31896));
    LocalMux I__6518 (
            .O(N__31896),
            .I(N__31892));
    InMux I__6517 (
            .O(N__31895),
            .I(N__31887));
    Span4Mux_h I__6516 (
            .O(N__31892),
            .I(N__31884));
    InMux I__6515 (
            .O(N__31891),
            .I(N__31879));
    InMux I__6514 (
            .O(N__31890),
            .I(N__31879));
    LocalMux I__6513 (
            .O(N__31887),
            .I(N__31876));
    Odrv4 I__6512 (
            .O(N__31884),
            .I(\c0.rx.n17022 ));
    LocalMux I__6511 (
            .O(N__31879),
            .I(\c0.rx.n17022 ));
    Odrv4 I__6510 (
            .O(N__31876),
            .I(\c0.rx.n17022 ));
    CascadeMux I__6509 (
            .O(N__31869),
            .I(N__31863));
    InMux I__6508 (
            .O(N__31868),
            .I(N__31854));
    InMux I__6507 (
            .O(N__31867),
            .I(N__31854));
    InMux I__6506 (
            .O(N__31866),
            .I(N__31854));
    InMux I__6505 (
            .O(N__31863),
            .I(N__31854));
    LocalMux I__6504 (
            .O(N__31854),
            .I(N__31845));
    InMux I__6503 (
            .O(N__31853),
            .I(N__31842));
    InMux I__6502 (
            .O(N__31852),
            .I(N__31839));
    InMux I__6501 (
            .O(N__31851),
            .I(N__31836));
    InMux I__6500 (
            .O(N__31850),
            .I(N__31829));
    InMux I__6499 (
            .O(N__31849),
            .I(N__31829));
    InMux I__6498 (
            .O(N__31848),
            .I(N__31829));
    Span4Mux_s1_v I__6497 (
            .O(N__31845),
            .I(N__31826));
    LocalMux I__6496 (
            .O(N__31842),
            .I(N__31823));
    LocalMux I__6495 (
            .O(N__31839),
            .I(N__31818));
    LocalMux I__6494 (
            .O(N__31836),
            .I(N__31818));
    LocalMux I__6493 (
            .O(N__31829),
            .I(N__31815));
    Sp12to4 I__6492 (
            .O(N__31826),
            .I(N__31810));
    Span12Mux_s1_v I__6491 (
            .O(N__31823),
            .I(N__31810));
    Span4Mux_h I__6490 (
            .O(N__31818),
            .I(N__31805));
    Span4Mux_v I__6489 (
            .O(N__31815),
            .I(N__31805));
    Odrv12 I__6488 (
            .O(N__31810),
            .I(r_SM_Main_2));
    Odrv4 I__6487 (
            .O(N__31805),
            .I(r_SM_Main_2));
    SRMux I__6486 (
            .O(N__31800),
            .I(N__31797));
    LocalMux I__6485 (
            .O(N__31797),
            .I(N__31794));
    Span4Mux_h I__6484 (
            .O(N__31794),
            .I(N__31791));
    Span4Mux_h I__6483 (
            .O(N__31791),
            .I(N__31788));
    Odrv4 I__6482 (
            .O(N__31788),
            .I(\c0.rx.n17058 ));
    CascadeMux I__6481 (
            .O(N__31785),
            .I(N__31782));
    InMux I__6480 (
            .O(N__31782),
            .I(N__31776));
    InMux I__6479 (
            .O(N__31781),
            .I(N__31776));
    LocalMux I__6478 (
            .O(N__31776),
            .I(N__31771));
    InMux I__6477 (
            .O(N__31775),
            .I(N__31768));
    InMux I__6476 (
            .O(N__31774),
            .I(N__31764));
    Span4Mux_h I__6475 (
            .O(N__31771),
            .I(N__31761));
    LocalMux I__6474 (
            .O(N__31768),
            .I(N__31758));
    InMux I__6473 (
            .O(N__31767),
            .I(N__31755));
    LocalMux I__6472 (
            .O(N__31764),
            .I(N__31752));
    Span4Mux_h I__6471 (
            .O(N__31761),
            .I(N__31749));
    Span4Mux_h I__6470 (
            .O(N__31758),
            .I(N__31746));
    LocalMux I__6469 (
            .O(N__31755),
            .I(\c0.rx.r_Clock_Count_7 ));
    Odrv12 I__6468 (
            .O(N__31752),
            .I(\c0.rx.r_Clock_Count_7 ));
    Odrv4 I__6467 (
            .O(N__31749),
            .I(\c0.rx.r_Clock_Count_7 ));
    Odrv4 I__6466 (
            .O(N__31746),
            .I(\c0.rx.r_Clock_Count_7 ));
    InMux I__6465 (
            .O(N__31737),
            .I(N__31730));
    InMux I__6464 (
            .O(N__31736),
            .I(N__31730));
    InMux I__6463 (
            .O(N__31735),
            .I(N__31727));
    LocalMux I__6462 (
            .O(N__31730),
            .I(N__31723));
    LocalMux I__6461 (
            .O(N__31727),
            .I(N__31720));
    InMux I__6460 (
            .O(N__31726),
            .I(N__31716));
    Span4Mux_v I__6459 (
            .O(N__31723),
            .I(N__31713));
    Span4Mux_v I__6458 (
            .O(N__31720),
            .I(N__31710));
    InMux I__6457 (
            .O(N__31719),
            .I(N__31707));
    LocalMux I__6456 (
            .O(N__31716),
            .I(N__31698));
    Span4Mux_h I__6455 (
            .O(N__31713),
            .I(N__31698));
    Span4Mux_s0_v I__6454 (
            .O(N__31710),
            .I(N__31698));
    LocalMux I__6453 (
            .O(N__31707),
            .I(N__31698));
    Odrv4 I__6452 (
            .O(N__31698),
            .I(\c0.rx.r_Clock_Count_6 ));
    CascadeMux I__6451 (
            .O(N__31695),
            .I(N__31692));
    InMux I__6450 (
            .O(N__31692),
            .I(N__31686));
    InMux I__6449 (
            .O(N__31691),
            .I(N__31686));
    LocalMux I__6448 (
            .O(N__31686),
            .I(N__31683));
    Span4Mux_h I__6447 (
            .O(N__31683),
            .I(N__31680));
    Odrv4 I__6446 (
            .O(N__31680),
            .I(\c0.rx.n17080 ));
    InMux I__6445 (
            .O(N__31677),
            .I(N__31671));
    InMux I__6444 (
            .O(N__31676),
            .I(N__31668));
    InMux I__6443 (
            .O(N__31675),
            .I(N__31665));
    InMux I__6442 (
            .O(N__31674),
            .I(N__31662));
    LocalMux I__6441 (
            .O(N__31671),
            .I(N__31659));
    LocalMux I__6440 (
            .O(N__31668),
            .I(N__31656));
    LocalMux I__6439 (
            .O(N__31665),
            .I(N__31652));
    LocalMux I__6438 (
            .O(N__31662),
            .I(N__31649));
    Span4Mux_v I__6437 (
            .O(N__31659),
            .I(N__31646));
    Span4Mux_v I__6436 (
            .O(N__31656),
            .I(N__31643));
    InMux I__6435 (
            .O(N__31655),
            .I(N__31640));
    Span4Mux_h I__6434 (
            .O(N__31652),
            .I(N__31633));
    Span4Mux_v I__6433 (
            .O(N__31649),
            .I(N__31633));
    Span4Mux_h I__6432 (
            .O(N__31646),
            .I(N__31633));
    Odrv4 I__6431 (
            .O(N__31643),
            .I(rand_data_26));
    LocalMux I__6430 (
            .O(N__31640),
            .I(rand_data_26));
    Odrv4 I__6429 (
            .O(N__31633),
            .I(rand_data_26));
    InMux I__6428 (
            .O(N__31626),
            .I(n16035));
    InMux I__6427 (
            .O(N__31623),
            .I(N__31619));
    InMux I__6426 (
            .O(N__31622),
            .I(N__31615));
    LocalMux I__6425 (
            .O(N__31619),
            .I(N__31611));
    InMux I__6424 (
            .O(N__31618),
            .I(N__31608));
    LocalMux I__6423 (
            .O(N__31615),
            .I(N__31605));
    InMux I__6422 (
            .O(N__31614),
            .I(N__31602));
    Span4Mux_v I__6421 (
            .O(N__31611),
            .I(N__31597));
    LocalMux I__6420 (
            .O(N__31608),
            .I(N__31597));
    Span4Mux_v I__6419 (
            .O(N__31605),
            .I(N__31593));
    LocalMux I__6418 (
            .O(N__31602),
            .I(N__31590));
    Span4Mux_h I__6417 (
            .O(N__31597),
            .I(N__31587));
    InMux I__6416 (
            .O(N__31596),
            .I(N__31584));
    Span4Mux_v I__6415 (
            .O(N__31593),
            .I(N__31581));
    Span12Mux_s6_v I__6414 (
            .O(N__31590),
            .I(N__31578));
    Odrv4 I__6413 (
            .O(N__31587),
            .I(rand_data_27));
    LocalMux I__6412 (
            .O(N__31584),
            .I(rand_data_27));
    Odrv4 I__6411 (
            .O(N__31581),
            .I(rand_data_27));
    Odrv12 I__6410 (
            .O(N__31578),
            .I(rand_data_27));
    InMux I__6409 (
            .O(N__31569),
            .I(n16036));
    InMux I__6408 (
            .O(N__31566),
            .I(N__31560));
    InMux I__6407 (
            .O(N__31565),
            .I(N__31557));
    InMux I__6406 (
            .O(N__31564),
            .I(N__31554));
    InMux I__6405 (
            .O(N__31563),
            .I(N__31551));
    LocalMux I__6404 (
            .O(N__31560),
            .I(N__31548));
    LocalMux I__6403 (
            .O(N__31557),
            .I(N__31545));
    LocalMux I__6402 (
            .O(N__31554),
            .I(N__31539));
    LocalMux I__6401 (
            .O(N__31551),
            .I(N__31539));
    Span4Mux_h I__6400 (
            .O(N__31548),
            .I(N__31536));
    Span4Mux_v I__6399 (
            .O(N__31545),
            .I(N__31533));
    InMux I__6398 (
            .O(N__31544),
            .I(N__31530));
    Span4Mux_v I__6397 (
            .O(N__31539),
            .I(N__31525));
    Span4Mux_h I__6396 (
            .O(N__31536),
            .I(N__31525));
    Odrv4 I__6395 (
            .O(N__31533),
            .I(rand_data_28));
    LocalMux I__6394 (
            .O(N__31530),
            .I(rand_data_28));
    Odrv4 I__6393 (
            .O(N__31525),
            .I(rand_data_28));
    InMux I__6392 (
            .O(N__31518),
            .I(n16037));
    InMux I__6391 (
            .O(N__31515),
            .I(N__31510));
    InMux I__6390 (
            .O(N__31514),
            .I(N__31507));
    InMux I__6389 (
            .O(N__31513),
            .I(N__31503));
    LocalMux I__6388 (
            .O(N__31510),
            .I(N__31500));
    LocalMux I__6387 (
            .O(N__31507),
            .I(N__31497));
    InMux I__6386 (
            .O(N__31506),
            .I(N__31494));
    LocalMux I__6385 (
            .O(N__31503),
            .I(N__31491));
    Span4Mux_h I__6384 (
            .O(N__31500),
            .I(N__31488));
    Span4Mux_v I__6383 (
            .O(N__31497),
            .I(N__31483));
    LocalMux I__6382 (
            .O(N__31494),
            .I(N__31483));
    Span4Mux_h I__6381 (
            .O(N__31491),
            .I(N__31479));
    Span4Mux_v I__6380 (
            .O(N__31488),
            .I(N__31474));
    Span4Mux_h I__6379 (
            .O(N__31483),
            .I(N__31474));
    InMux I__6378 (
            .O(N__31482),
            .I(N__31471));
    Span4Mux_h I__6377 (
            .O(N__31479),
            .I(N__31468));
    Odrv4 I__6376 (
            .O(N__31474),
            .I(rand_data_29));
    LocalMux I__6375 (
            .O(N__31471),
            .I(rand_data_29));
    Odrv4 I__6374 (
            .O(N__31468),
            .I(rand_data_29));
    InMux I__6373 (
            .O(N__31461),
            .I(n16038));
    InMux I__6372 (
            .O(N__31458),
            .I(N__31455));
    LocalMux I__6371 (
            .O(N__31455),
            .I(N__31450));
    InMux I__6370 (
            .O(N__31454),
            .I(N__31446));
    InMux I__6369 (
            .O(N__31453),
            .I(N__31443));
    Span4Mux_s1_h I__6368 (
            .O(N__31450),
            .I(N__31440));
    InMux I__6367 (
            .O(N__31449),
            .I(N__31437));
    LocalMux I__6366 (
            .O(N__31446),
            .I(N__31434));
    LocalMux I__6365 (
            .O(N__31443),
            .I(N__31431));
    Span4Mux_v I__6364 (
            .O(N__31440),
            .I(N__31425));
    LocalMux I__6363 (
            .O(N__31437),
            .I(N__31425));
    Span4Mux_v I__6362 (
            .O(N__31434),
            .I(N__31422));
    Span4Mux_v I__6361 (
            .O(N__31431),
            .I(N__31419));
    InMux I__6360 (
            .O(N__31430),
            .I(N__31416));
    Span4Mux_h I__6359 (
            .O(N__31425),
            .I(N__31411));
    Span4Mux_h I__6358 (
            .O(N__31422),
            .I(N__31411));
    Odrv4 I__6357 (
            .O(N__31419),
            .I(rand_data_30));
    LocalMux I__6356 (
            .O(N__31416),
            .I(rand_data_30));
    Odrv4 I__6355 (
            .O(N__31411),
            .I(rand_data_30));
    InMux I__6354 (
            .O(N__31404),
            .I(n16039));
    InMux I__6353 (
            .O(N__31401),
            .I(N__31396));
    InMux I__6352 (
            .O(N__31400),
            .I(N__31393));
    InMux I__6351 (
            .O(N__31399),
            .I(N__31389));
    LocalMux I__6350 (
            .O(N__31396),
            .I(N__31386));
    LocalMux I__6349 (
            .O(N__31393),
            .I(N__31383));
    InMux I__6348 (
            .O(N__31392),
            .I(N__31380));
    LocalMux I__6347 (
            .O(N__31389),
            .I(N__31377));
    Span4Mux_h I__6346 (
            .O(N__31386),
            .I(N__31373));
    Span4Mux_v I__6345 (
            .O(N__31383),
            .I(N__31368));
    LocalMux I__6344 (
            .O(N__31380),
            .I(N__31368));
    Span4Mux_v I__6343 (
            .O(N__31377),
            .I(N__31365));
    InMux I__6342 (
            .O(N__31376),
            .I(N__31362));
    Span4Mux_h I__6341 (
            .O(N__31373),
            .I(N__31357));
    Span4Mux_h I__6340 (
            .O(N__31368),
            .I(N__31357));
    Sp12to4 I__6339 (
            .O(N__31365),
            .I(N__31354));
    LocalMux I__6338 (
            .O(N__31362),
            .I(rand_data_31));
    Odrv4 I__6337 (
            .O(N__31357),
            .I(rand_data_31));
    Odrv12 I__6336 (
            .O(N__31354),
            .I(rand_data_31));
    InMux I__6335 (
            .O(N__31347),
            .I(n16040));
    InMux I__6334 (
            .O(N__31344),
            .I(N__31341));
    LocalMux I__6333 (
            .O(N__31341),
            .I(N__31338));
    Span4Mux_s2_v I__6332 (
            .O(N__31338),
            .I(N__31335));
    Span4Mux_h I__6331 (
            .O(N__31335),
            .I(N__31331));
    InMux I__6330 (
            .O(N__31334),
            .I(N__31328));
    Span4Mux_h I__6329 (
            .O(N__31331),
            .I(N__31325));
    LocalMux I__6328 (
            .O(N__31328),
            .I(rand_setpoint_31));
    Odrv4 I__6327 (
            .O(N__31325),
            .I(rand_setpoint_31));
    InMux I__6326 (
            .O(N__31320),
            .I(N__31316));
    CascadeMux I__6325 (
            .O(N__31319),
            .I(N__31313));
    LocalMux I__6324 (
            .O(N__31316),
            .I(N__31310));
    InMux I__6323 (
            .O(N__31313),
            .I(N__31307));
    Odrv4 I__6322 (
            .O(N__31310),
            .I(rand_setpoint_26));
    LocalMux I__6321 (
            .O(N__31307),
            .I(rand_setpoint_26));
    CascadeMux I__6320 (
            .O(N__31302),
            .I(N__31298));
    InMux I__6319 (
            .O(N__31301),
            .I(N__31295));
    InMux I__6318 (
            .O(N__31298),
            .I(N__31292));
    LocalMux I__6317 (
            .O(N__31295),
            .I(rand_setpoint_29));
    LocalMux I__6316 (
            .O(N__31292),
            .I(rand_setpoint_29));
    CascadeMux I__6315 (
            .O(N__31287),
            .I(N__31283));
    InMux I__6314 (
            .O(N__31286),
            .I(N__31280));
    InMux I__6313 (
            .O(N__31283),
            .I(N__31277));
    LocalMux I__6312 (
            .O(N__31280),
            .I(rand_setpoint_27));
    LocalMux I__6311 (
            .O(N__31277),
            .I(rand_setpoint_27));
    InMux I__6310 (
            .O(N__31272),
            .I(N__31269));
    LocalMux I__6309 (
            .O(N__31269),
            .I(N__31265));
    InMux I__6308 (
            .O(N__31268),
            .I(N__31260));
    Span4Mux_v I__6307 (
            .O(N__31265),
            .I(N__31257));
    InMux I__6306 (
            .O(N__31264),
            .I(N__31254));
    InMux I__6305 (
            .O(N__31263),
            .I(N__31251));
    LocalMux I__6304 (
            .O(N__31260),
            .I(N__31248));
    Span4Mux_v I__6303 (
            .O(N__31257),
            .I(N__31245));
    LocalMux I__6302 (
            .O(N__31254),
            .I(N__31242));
    LocalMux I__6301 (
            .O(N__31251),
            .I(N__31239));
    Span4Mux_v I__6300 (
            .O(N__31248),
            .I(N__31235));
    Span4Mux_s3_h I__6299 (
            .O(N__31245),
            .I(N__31232));
    Span4Mux_v I__6298 (
            .O(N__31242),
            .I(N__31227));
    Span4Mux_h I__6297 (
            .O(N__31239),
            .I(N__31227));
    InMux I__6296 (
            .O(N__31238),
            .I(N__31224));
    Span4Mux_h I__6295 (
            .O(N__31235),
            .I(N__31221));
    Odrv4 I__6294 (
            .O(N__31232),
            .I(rand_data_18));
    Odrv4 I__6293 (
            .O(N__31227),
            .I(rand_data_18));
    LocalMux I__6292 (
            .O(N__31224),
            .I(rand_data_18));
    Odrv4 I__6291 (
            .O(N__31221),
            .I(rand_data_18));
    InMux I__6290 (
            .O(N__31212),
            .I(n16027));
    InMux I__6289 (
            .O(N__31209),
            .I(N__31205));
    InMux I__6288 (
            .O(N__31208),
            .I(N__31202));
    LocalMux I__6287 (
            .O(N__31205),
            .I(N__31198));
    LocalMux I__6286 (
            .O(N__31202),
            .I(N__31195));
    InMux I__6285 (
            .O(N__31201),
            .I(N__31191));
    Span4Mux_h I__6284 (
            .O(N__31198),
            .I(N__31188));
    Span4Mux_h I__6283 (
            .O(N__31195),
            .I(N__31185));
    InMux I__6282 (
            .O(N__31194),
            .I(N__31182));
    LocalMux I__6281 (
            .O(N__31191),
            .I(N__31178));
    Sp12to4 I__6280 (
            .O(N__31188),
            .I(N__31171));
    Sp12to4 I__6279 (
            .O(N__31185),
            .I(N__31171));
    LocalMux I__6278 (
            .O(N__31182),
            .I(N__31171));
    InMux I__6277 (
            .O(N__31181),
            .I(N__31168));
    Span12Mux_s7_v I__6276 (
            .O(N__31178),
            .I(N__31165));
    Odrv12 I__6275 (
            .O(N__31171),
            .I(rand_data_19));
    LocalMux I__6274 (
            .O(N__31168),
            .I(rand_data_19));
    Odrv12 I__6273 (
            .O(N__31165),
            .I(rand_data_19));
    InMux I__6272 (
            .O(N__31158),
            .I(n16028));
    CascadeMux I__6271 (
            .O(N__31155),
            .I(N__31151));
    InMux I__6270 (
            .O(N__31154),
            .I(N__31146));
    InMux I__6269 (
            .O(N__31151),
            .I(N__31143));
    InMux I__6268 (
            .O(N__31150),
            .I(N__31140));
    InMux I__6267 (
            .O(N__31149),
            .I(N__31137));
    LocalMux I__6266 (
            .O(N__31146),
            .I(N__31134));
    LocalMux I__6265 (
            .O(N__31143),
            .I(N__31131));
    LocalMux I__6264 (
            .O(N__31140),
            .I(N__31128));
    LocalMux I__6263 (
            .O(N__31137),
            .I(N__31124));
    Span4Mux_v I__6262 (
            .O(N__31134),
            .I(N__31121));
    Span4Mux_h I__6261 (
            .O(N__31131),
            .I(N__31118));
    Span4Mux_v I__6260 (
            .O(N__31128),
            .I(N__31115));
    InMux I__6259 (
            .O(N__31127),
            .I(N__31112));
    Span4Mux_v I__6258 (
            .O(N__31124),
            .I(N__31107));
    Span4Mux_h I__6257 (
            .O(N__31121),
            .I(N__31107));
    Odrv4 I__6256 (
            .O(N__31118),
            .I(rand_data_20));
    Odrv4 I__6255 (
            .O(N__31115),
            .I(rand_data_20));
    LocalMux I__6254 (
            .O(N__31112),
            .I(rand_data_20));
    Odrv4 I__6253 (
            .O(N__31107),
            .I(rand_data_20));
    InMux I__6252 (
            .O(N__31098),
            .I(n16029));
    InMux I__6251 (
            .O(N__31095),
            .I(N__31091));
    InMux I__6250 (
            .O(N__31094),
            .I(N__31086));
    LocalMux I__6249 (
            .O(N__31091),
            .I(N__31083));
    InMux I__6248 (
            .O(N__31090),
            .I(N__31080));
    InMux I__6247 (
            .O(N__31089),
            .I(N__31077));
    LocalMux I__6246 (
            .O(N__31086),
            .I(N__31074));
    Span4Mux_h I__6245 (
            .O(N__31083),
            .I(N__31071));
    LocalMux I__6244 (
            .O(N__31080),
            .I(N__31068));
    LocalMux I__6243 (
            .O(N__31077),
            .I(N__31065));
    Span4Mux_h I__6242 (
            .O(N__31074),
            .I(N__31061));
    Span4Mux_v I__6241 (
            .O(N__31071),
            .I(N__31058));
    Span4Mux_v I__6240 (
            .O(N__31068),
            .I(N__31055));
    Span4Mux_h I__6239 (
            .O(N__31065),
            .I(N__31052));
    InMux I__6238 (
            .O(N__31064),
            .I(N__31049));
    Span4Mux_h I__6237 (
            .O(N__31061),
            .I(N__31046));
    Odrv4 I__6236 (
            .O(N__31058),
            .I(rand_data_21));
    Odrv4 I__6235 (
            .O(N__31055),
            .I(rand_data_21));
    Odrv4 I__6234 (
            .O(N__31052),
            .I(rand_data_21));
    LocalMux I__6233 (
            .O(N__31049),
            .I(rand_data_21));
    Odrv4 I__6232 (
            .O(N__31046),
            .I(rand_data_21));
    InMux I__6231 (
            .O(N__31035),
            .I(n16030));
    CascadeMux I__6230 (
            .O(N__31032),
            .I(N__31027));
    InMux I__6229 (
            .O(N__31031),
            .I(N__31023));
    InMux I__6228 (
            .O(N__31030),
            .I(N__31020));
    InMux I__6227 (
            .O(N__31027),
            .I(N__31017));
    InMux I__6226 (
            .O(N__31026),
            .I(N__31014));
    LocalMux I__6225 (
            .O(N__31023),
            .I(N__31011));
    LocalMux I__6224 (
            .O(N__31020),
            .I(N__31008));
    LocalMux I__6223 (
            .O(N__31017),
            .I(N__31003));
    LocalMux I__6222 (
            .O(N__31014),
            .I(N__31003));
    Span4Mux_h I__6221 (
            .O(N__31011),
            .I(N__30999));
    Span4Mux_v I__6220 (
            .O(N__31008),
            .I(N__30996));
    Span4Mux_v I__6219 (
            .O(N__31003),
            .I(N__30993));
    InMux I__6218 (
            .O(N__31002),
            .I(N__30990));
    Span4Mux_h I__6217 (
            .O(N__30999),
            .I(N__30987));
    Odrv4 I__6216 (
            .O(N__30996),
            .I(rand_data_22));
    Odrv4 I__6215 (
            .O(N__30993),
            .I(rand_data_22));
    LocalMux I__6214 (
            .O(N__30990),
            .I(rand_data_22));
    Odrv4 I__6213 (
            .O(N__30987),
            .I(rand_data_22));
    InMux I__6212 (
            .O(N__30978),
            .I(n16031));
    InMux I__6211 (
            .O(N__30975),
            .I(N__30971));
    InMux I__6210 (
            .O(N__30974),
            .I(N__30967));
    LocalMux I__6209 (
            .O(N__30971),
            .I(N__30964));
    InMux I__6208 (
            .O(N__30970),
            .I(N__30961));
    LocalMux I__6207 (
            .O(N__30967),
            .I(N__30957));
    Span4Mux_h I__6206 (
            .O(N__30964),
            .I(N__30952));
    LocalMux I__6205 (
            .O(N__30961),
            .I(N__30952));
    InMux I__6204 (
            .O(N__30960),
            .I(N__30949));
    Span4Mux_h I__6203 (
            .O(N__30957),
            .I(N__30945));
    Span4Mux_v I__6202 (
            .O(N__30952),
            .I(N__30942));
    LocalMux I__6201 (
            .O(N__30949),
            .I(N__30939));
    InMux I__6200 (
            .O(N__30948),
            .I(N__30936));
    Span4Mux_h I__6199 (
            .O(N__30945),
            .I(N__30933));
    Odrv4 I__6198 (
            .O(N__30942),
            .I(rand_data_23));
    Odrv12 I__6197 (
            .O(N__30939),
            .I(rand_data_23));
    LocalMux I__6196 (
            .O(N__30936),
            .I(rand_data_23));
    Odrv4 I__6195 (
            .O(N__30933),
            .I(rand_data_23));
    InMux I__6194 (
            .O(N__30924),
            .I(n16032));
    InMux I__6193 (
            .O(N__30921),
            .I(N__30916));
    InMux I__6192 (
            .O(N__30920),
            .I(N__30912));
    InMux I__6191 (
            .O(N__30919),
            .I(N__30909));
    LocalMux I__6190 (
            .O(N__30916),
            .I(N__30906));
    InMux I__6189 (
            .O(N__30915),
            .I(N__30903));
    LocalMux I__6188 (
            .O(N__30912),
            .I(N__30900));
    LocalMux I__6187 (
            .O(N__30909),
            .I(N__30896));
    Span4Mux_v I__6186 (
            .O(N__30906),
            .I(N__30891));
    LocalMux I__6185 (
            .O(N__30903),
            .I(N__30891));
    Span4Mux_h I__6184 (
            .O(N__30900),
            .I(N__30888));
    InMux I__6183 (
            .O(N__30899),
            .I(N__30885));
    Span4Mux_v I__6182 (
            .O(N__30896),
            .I(N__30878));
    Span4Mux_h I__6181 (
            .O(N__30891),
            .I(N__30878));
    Span4Mux_h I__6180 (
            .O(N__30888),
            .I(N__30878));
    LocalMux I__6179 (
            .O(N__30885),
            .I(rand_data_24));
    Odrv4 I__6178 (
            .O(N__30878),
            .I(rand_data_24));
    InMux I__6177 (
            .O(N__30873),
            .I(N__30870));
    LocalMux I__6176 (
            .O(N__30870),
            .I(N__30867));
    Span4Mux_s2_v I__6175 (
            .O(N__30867),
            .I(N__30864));
    Span4Mux_h I__6174 (
            .O(N__30864),
            .I(N__30860));
    CascadeMux I__6173 (
            .O(N__30863),
            .I(N__30857));
    Span4Mux_h I__6172 (
            .O(N__30860),
            .I(N__30854));
    InMux I__6171 (
            .O(N__30857),
            .I(N__30851));
    Odrv4 I__6170 (
            .O(N__30854),
            .I(rand_setpoint_24));
    LocalMux I__6169 (
            .O(N__30851),
            .I(rand_setpoint_24));
    InMux I__6168 (
            .O(N__30846),
            .I(bfn_10_28_0_));
    InMux I__6167 (
            .O(N__30843),
            .I(N__30839));
    InMux I__6166 (
            .O(N__30842),
            .I(N__30835));
    LocalMux I__6165 (
            .O(N__30839),
            .I(N__30831));
    InMux I__6164 (
            .O(N__30838),
            .I(N__30828));
    LocalMux I__6163 (
            .O(N__30835),
            .I(N__30825));
    InMux I__6162 (
            .O(N__30834),
            .I(N__30822));
    Span4Mux_v I__6161 (
            .O(N__30831),
            .I(N__30819));
    LocalMux I__6160 (
            .O(N__30828),
            .I(N__30816));
    Span4Mux_v I__6159 (
            .O(N__30825),
            .I(N__30811));
    LocalMux I__6158 (
            .O(N__30822),
            .I(N__30811));
    Span4Mux_s0_h I__6157 (
            .O(N__30819),
            .I(N__30807));
    Span4Mux_h I__6156 (
            .O(N__30816),
            .I(N__30804));
    Span4Mux_v I__6155 (
            .O(N__30811),
            .I(N__30801));
    InMux I__6154 (
            .O(N__30810),
            .I(N__30798));
    Span4Mux_h I__6153 (
            .O(N__30807),
            .I(N__30793));
    Span4Mux_h I__6152 (
            .O(N__30804),
            .I(N__30793));
    Odrv4 I__6151 (
            .O(N__30801),
            .I(rand_data_25));
    LocalMux I__6150 (
            .O(N__30798),
            .I(rand_data_25));
    Odrv4 I__6149 (
            .O(N__30793),
            .I(rand_data_25));
    InMux I__6148 (
            .O(N__30786),
            .I(n16034));
    InMux I__6147 (
            .O(N__30783),
            .I(N__30776));
    InMux I__6146 (
            .O(N__30782),
            .I(N__30773));
    InMux I__6145 (
            .O(N__30781),
            .I(N__30770));
    InMux I__6144 (
            .O(N__30780),
            .I(N__30767));
    InMux I__6143 (
            .O(N__30779),
            .I(N__30764));
    LocalMux I__6142 (
            .O(N__30776),
            .I(N__30761));
    LocalMux I__6141 (
            .O(N__30773),
            .I(N__30758));
    LocalMux I__6140 (
            .O(N__30770),
            .I(N__30755));
    LocalMux I__6139 (
            .O(N__30767),
            .I(N__30752));
    LocalMux I__6138 (
            .O(N__30764),
            .I(N__30748));
    Span4Mux_h I__6137 (
            .O(N__30761),
            .I(N__30743));
    Span4Mux_h I__6136 (
            .O(N__30758),
            .I(N__30743));
    Span12Mux_h I__6135 (
            .O(N__30755),
            .I(N__30740));
    Span4Mux_h I__6134 (
            .O(N__30752),
            .I(N__30737));
    InMux I__6133 (
            .O(N__30751),
            .I(N__30734));
    Span12Mux_h I__6132 (
            .O(N__30748),
            .I(N__30731));
    Odrv4 I__6131 (
            .O(N__30743),
            .I(rand_data_10));
    Odrv12 I__6130 (
            .O(N__30740),
            .I(rand_data_10));
    Odrv4 I__6129 (
            .O(N__30737),
            .I(rand_data_10));
    LocalMux I__6128 (
            .O(N__30734),
            .I(rand_data_10));
    Odrv12 I__6127 (
            .O(N__30731),
            .I(rand_data_10));
    InMux I__6126 (
            .O(N__30720),
            .I(n16019));
    InMux I__6125 (
            .O(N__30717),
            .I(N__30713));
    InMux I__6124 (
            .O(N__30716),
            .I(N__30710));
    LocalMux I__6123 (
            .O(N__30713),
            .I(N__30704));
    LocalMux I__6122 (
            .O(N__30710),
            .I(N__30701));
    InMux I__6121 (
            .O(N__30709),
            .I(N__30698));
    InMux I__6120 (
            .O(N__30708),
            .I(N__30695));
    InMux I__6119 (
            .O(N__30707),
            .I(N__30692));
    Span4Mux_v I__6118 (
            .O(N__30704),
            .I(N__30689));
    Span4Mux_h I__6117 (
            .O(N__30701),
            .I(N__30682));
    LocalMux I__6116 (
            .O(N__30698),
            .I(N__30682));
    LocalMux I__6115 (
            .O(N__30695),
            .I(N__30682));
    LocalMux I__6114 (
            .O(N__30692),
            .I(N__30678));
    Span4Mux_h I__6113 (
            .O(N__30689),
            .I(N__30673));
    Span4Mux_h I__6112 (
            .O(N__30682),
            .I(N__30673));
    InMux I__6111 (
            .O(N__30681),
            .I(N__30670));
    Span12Mux_s8_v I__6110 (
            .O(N__30678),
            .I(N__30667));
    Odrv4 I__6109 (
            .O(N__30673),
            .I(rand_data_11));
    LocalMux I__6108 (
            .O(N__30670),
            .I(rand_data_11));
    Odrv12 I__6107 (
            .O(N__30667),
            .I(rand_data_11));
    InMux I__6106 (
            .O(N__30660),
            .I(n16020));
    InMux I__6105 (
            .O(N__30657),
            .I(N__30650));
    InMux I__6104 (
            .O(N__30656),
            .I(N__30650));
    InMux I__6103 (
            .O(N__30655),
            .I(N__30647));
    LocalMux I__6102 (
            .O(N__30650),
            .I(N__30642));
    LocalMux I__6101 (
            .O(N__30647),
            .I(N__30639));
    InMux I__6100 (
            .O(N__30646),
            .I(N__30636));
    InMux I__6099 (
            .O(N__30645),
            .I(N__30633));
    Span4Mux_v I__6098 (
            .O(N__30642),
            .I(N__30630));
    Span4Mux_h I__6097 (
            .O(N__30639),
            .I(N__30626));
    LocalMux I__6096 (
            .O(N__30636),
            .I(N__30621));
    LocalMux I__6095 (
            .O(N__30633),
            .I(N__30621));
    Sp12to4 I__6094 (
            .O(N__30630),
            .I(N__30618));
    InMux I__6093 (
            .O(N__30629),
            .I(N__30615));
    Span4Mux_h I__6092 (
            .O(N__30626),
            .I(N__30612));
    Odrv12 I__6091 (
            .O(N__30621),
            .I(rand_data_12));
    Odrv12 I__6090 (
            .O(N__30618),
            .I(rand_data_12));
    LocalMux I__6089 (
            .O(N__30615),
            .I(rand_data_12));
    Odrv4 I__6088 (
            .O(N__30612),
            .I(rand_data_12));
    InMux I__6087 (
            .O(N__30603),
            .I(n16021));
    InMux I__6086 (
            .O(N__30600),
            .I(N__30595));
    InMux I__6085 (
            .O(N__30599),
            .I(N__30591));
    InMux I__6084 (
            .O(N__30598),
            .I(N__30588));
    LocalMux I__6083 (
            .O(N__30595),
            .I(N__30585));
    InMux I__6082 (
            .O(N__30594),
            .I(N__30581));
    LocalMux I__6081 (
            .O(N__30591),
            .I(N__30578));
    LocalMux I__6080 (
            .O(N__30588),
            .I(N__30575));
    Span4Mux_h I__6079 (
            .O(N__30585),
            .I(N__30571));
    InMux I__6078 (
            .O(N__30584),
            .I(N__30568));
    LocalMux I__6077 (
            .O(N__30581),
            .I(N__30565));
    Span4Mux_h I__6076 (
            .O(N__30578),
            .I(N__30562));
    Span4Mux_v I__6075 (
            .O(N__30575),
            .I(N__30559));
    InMux I__6074 (
            .O(N__30574),
            .I(N__30556));
    Span4Mux_h I__6073 (
            .O(N__30571),
            .I(N__30553));
    LocalMux I__6072 (
            .O(N__30568),
            .I(rand_data_13));
    Odrv12 I__6071 (
            .O(N__30565),
            .I(rand_data_13));
    Odrv4 I__6070 (
            .O(N__30562),
            .I(rand_data_13));
    Odrv4 I__6069 (
            .O(N__30559),
            .I(rand_data_13));
    LocalMux I__6068 (
            .O(N__30556),
            .I(rand_data_13));
    Odrv4 I__6067 (
            .O(N__30553),
            .I(rand_data_13));
    InMux I__6066 (
            .O(N__30540),
            .I(n16022));
    CascadeMux I__6065 (
            .O(N__30537),
            .I(N__30530));
    InMux I__6064 (
            .O(N__30536),
            .I(N__30527));
    InMux I__6063 (
            .O(N__30535),
            .I(N__30524));
    InMux I__6062 (
            .O(N__30534),
            .I(N__30521));
    InMux I__6061 (
            .O(N__30533),
            .I(N__30518));
    InMux I__6060 (
            .O(N__30530),
            .I(N__30515));
    LocalMux I__6059 (
            .O(N__30527),
            .I(N__30512));
    LocalMux I__6058 (
            .O(N__30524),
            .I(N__30509));
    LocalMux I__6057 (
            .O(N__30521),
            .I(N__30506));
    LocalMux I__6056 (
            .O(N__30518),
            .I(N__30503));
    LocalMux I__6055 (
            .O(N__30515),
            .I(N__30497));
    Span4Mux_h I__6054 (
            .O(N__30512),
            .I(N__30497));
    Span4Mux_v I__6053 (
            .O(N__30509),
            .I(N__30494));
    Span4Mux_h I__6052 (
            .O(N__30506),
            .I(N__30491));
    Sp12to4 I__6051 (
            .O(N__30503),
            .I(N__30488));
    InMux I__6050 (
            .O(N__30502),
            .I(N__30485));
    Span4Mux_v I__6049 (
            .O(N__30497),
            .I(N__30480));
    Span4Mux_h I__6048 (
            .O(N__30494),
            .I(N__30480));
    Odrv4 I__6047 (
            .O(N__30491),
            .I(rand_data_14));
    Odrv12 I__6046 (
            .O(N__30488),
            .I(rand_data_14));
    LocalMux I__6045 (
            .O(N__30485),
            .I(rand_data_14));
    Odrv4 I__6044 (
            .O(N__30480),
            .I(rand_data_14));
    InMux I__6043 (
            .O(N__30471),
            .I(n16023));
    InMux I__6042 (
            .O(N__30468),
            .I(N__30462));
    InMux I__6041 (
            .O(N__30467),
            .I(N__30459));
    InMux I__6040 (
            .O(N__30466),
            .I(N__30454));
    InMux I__6039 (
            .O(N__30465),
            .I(N__30454));
    LocalMux I__6038 (
            .O(N__30462),
            .I(N__30451));
    LocalMux I__6037 (
            .O(N__30459),
            .I(N__30448));
    LocalMux I__6036 (
            .O(N__30454),
            .I(N__30443));
    Span4Mux_v I__6035 (
            .O(N__30451),
            .I(N__30440));
    Span4Mux_v I__6034 (
            .O(N__30448),
            .I(N__30437));
    InMux I__6033 (
            .O(N__30447),
            .I(N__30434));
    InMux I__6032 (
            .O(N__30446),
            .I(N__30431));
    Span4Mux_s2_h I__6031 (
            .O(N__30443),
            .I(N__30426));
    Span4Mux_h I__6030 (
            .O(N__30440),
            .I(N__30426));
    Odrv4 I__6029 (
            .O(N__30437),
            .I(rand_data_15));
    LocalMux I__6028 (
            .O(N__30434),
            .I(rand_data_15));
    LocalMux I__6027 (
            .O(N__30431),
            .I(rand_data_15));
    Odrv4 I__6026 (
            .O(N__30426),
            .I(rand_data_15));
    InMux I__6025 (
            .O(N__30417),
            .I(n16024));
    InMux I__6024 (
            .O(N__30414),
            .I(N__30410));
    InMux I__6023 (
            .O(N__30413),
            .I(N__30407));
    LocalMux I__6022 (
            .O(N__30410),
            .I(N__30402));
    LocalMux I__6021 (
            .O(N__30407),
            .I(N__30399));
    InMux I__6020 (
            .O(N__30406),
            .I(N__30396));
    InMux I__6019 (
            .O(N__30405),
            .I(N__30393));
    Span4Mux_h I__6018 (
            .O(N__30402),
            .I(N__30389));
    Span12Mux_s4_h I__6017 (
            .O(N__30399),
            .I(N__30384));
    LocalMux I__6016 (
            .O(N__30396),
            .I(N__30384));
    LocalMux I__6015 (
            .O(N__30393),
            .I(N__30381));
    InMux I__6014 (
            .O(N__30392),
            .I(N__30378));
    Span4Mux_h I__6013 (
            .O(N__30389),
            .I(N__30375));
    Odrv12 I__6012 (
            .O(N__30384),
            .I(rand_data_16));
    Odrv12 I__6011 (
            .O(N__30381),
            .I(rand_data_16));
    LocalMux I__6010 (
            .O(N__30378),
            .I(rand_data_16));
    Odrv4 I__6009 (
            .O(N__30375),
            .I(rand_data_16));
    InMux I__6008 (
            .O(N__30366),
            .I(bfn_10_27_0_));
    InMux I__6007 (
            .O(N__30363),
            .I(N__30360));
    LocalMux I__6006 (
            .O(N__30360),
            .I(N__30356));
    InMux I__6005 (
            .O(N__30359),
            .I(N__30352));
    Span4Mux_h I__6004 (
            .O(N__30356),
            .I(N__30348));
    InMux I__6003 (
            .O(N__30355),
            .I(N__30345));
    LocalMux I__6002 (
            .O(N__30352),
            .I(N__30342));
    CascadeMux I__6001 (
            .O(N__30351),
            .I(N__30339));
    Span4Mux_v I__6000 (
            .O(N__30348),
            .I(N__30336));
    LocalMux I__5999 (
            .O(N__30345),
            .I(N__30333));
    Span4Mux_h I__5998 (
            .O(N__30342),
            .I(N__30330));
    InMux I__5997 (
            .O(N__30339),
            .I(N__30326));
    Span4Mux_v I__5996 (
            .O(N__30336),
            .I(N__30321));
    Span4Mux_h I__5995 (
            .O(N__30333),
            .I(N__30321));
    Span4Mux_v I__5994 (
            .O(N__30330),
            .I(N__30318));
    InMux I__5993 (
            .O(N__30329),
            .I(N__30315));
    LocalMux I__5992 (
            .O(N__30326),
            .I(N__30310));
    Span4Mux_h I__5991 (
            .O(N__30321),
            .I(N__30310));
    Odrv4 I__5990 (
            .O(N__30318),
            .I(rand_data_17));
    LocalMux I__5989 (
            .O(N__30315),
            .I(rand_data_17));
    Odrv4 I__5988 (
            .O(N__30310),
            .I(rand_data_17));
    InMux I__5987 (
            .O(N__30303),
            .I(N__30300));
    LocalMux I__5986 (
            .O(N__30300),
            .I(N__30296));
    CascadeMux I__5985 (
            .O(N__30299),
            .I(N__30293));
    Span4Mux_v I__5984 (
            .O(N__30296),
            .I(N__30290));
    InMux I__5983 (
            .O(N__30293),
            .I(N__30287));
    Odrv4 I__5982 (
            .O(N__30290),
            .I(rand_setpoint_17));
    LocalMux I__5981 (
            .O(N__30287),
            .I(rand_setpoint_17));
    InMux I__5980 (
            .O(N__30282),
            .I(n16026));
    InMux I__5979 (
            .O(N__30279),
            .I(N__30275));
    InMux I__5978 (
            .O(N__30278),
            .I(N__30271));
    LocalMux I__5977 (
            .O(N__30275),
            .I(N__30268));
    CascadeMux I__5976 (
            .O(N__30274),
            .I(N__30265));
    LocalMux I__5975 (
            .O(N__30271),
            .I(N__30261));
    Span4Mux_v I__5974 (
            .O(N__30268),
            .I(N__30258));
    InMux I__5973 (
            .O(N__30265),
            .I(N__30254));
    InMux I__5972 (
            .O(N__30264),
            .I(N__30251));
    Span4Mux_v I__5971 (
            .O(N__30261),
            .I(N__30247));
    Span4Mux_h I__5970 (
            .O(N__30258),
            .I(N__30244));
    InMux I__5969 (
            .O(N__30257),
            .I(N__30241));
    LocalMux I__5968 (
            .O(N__30254),
            .I(N__30236));
    LocalMux I__5967 (
            .O(N__30251),
            .I(N__30236));
    InMux I__5966 (
            .O(N__30250),
            .I(N__30233));
    Span4Mux_s2_h I__5965 (
            .O(N__30247),
            .I(N__30228));
    Span4Mux_h I__5964 (
            .O(N__30244),
            .I(N__30228));
    LocalMux I__5963 (
            .O(N__30241),
            .I(rand_data_1));
    Odrv12 I__5962 (
            .O(N__30236),
            .I(rand_data_1));
    LocalMux I__5961 (
            .O(N__30233),
            .I(rand_data_1));
    Odrv4 I__5960 (
            .O(N__30228),
            .I(rand_data_1));
    InMux I__5959 (
            .O(N__30219),
            .I(n16010));
    InMux I__5958 (
            .O(N__30216),
            .I(N__30212));
    InMux I__5957 (
            .O(N__30215),
            .I(N__30206));
    LocalMux I__5956 (
            .O(N__30212),
            .I(N__30202));
    InMux I__5955 (
            .O(N__30211),
            .I(N__30197));
    InMux I__5954 (
            .O(N__30210),
            .I(N__30197));
    InMux I__5953 (
            .O(N__30209),
            .I(N__30194));
    LocalMux I__5952 (
            .O(N__30206),
            .I(N__30191));
    InMux I__5951 (
            .O(N__30205),
            .I(N__30188));
    Span12Mux_h I__5950 (
            .O(N__30202),
            .I(N__30185));
    LocalMux I__5949 (
            .O(N__30197),
            .I(rand_data_2));
    LocalMux I__5948 (
            .O(N__30194),
            .I(rand_data_2));
    Odrv4 I__5947 (
            .O(N__30191),
            .I(rand_data_2));
    LocalMux I__5946 (
            .O(N__30188),
            .I(rand_data_2));
    Odrv12 I__5945 (
            .O(N__30185),
            .I(rand_data_2));
    InMux I__5944 (
            .O(N__30174),
            .I(n16011));
    InMux I__5943 (
            .O(N__30171),
            .I(N__30166));
    InMux I__5942 (
            .O(N__30170),
            .I(N__30163));
    InMux I__5941 (
            .O(N__30169),
            .I(N__30159));
    LocalMux I__5940 (
            .O(N__30166),
            .I(N__30153));
    LocalMux I__5939 (
            .O(N__30163),
            .I(N__30153));
    InMux I__5938 (
            .O(N__30162),
            .I(N__30150));
    LocalMux I__5937 (
            .O(N__30159),
            .I(N__30147));
    InMux I__5936 (
            .O(N__30158),
            .I(N__30144));
    Span4Mux_v I__5935 (
            .O(N__30153),
            .I(N__30140));
    LocalMux I__5934 (
            .O(N__30150),
            .I(N__30137));
    Span4Mux_h I__5933 (
            .O(N__30147),
            .I(N__30134));
    LocalMux I__5932 (
            .O(N__30144),
            .I(N__30131));
    InMux I__5931 (
            .O(N__30143),
            .I(N__30128));
    Sp12to4 I__5930 (
            .O(N__30140),
            .I(N__30123));
    Span12Mux_s9_v I__5929 (
            .O(N__30137),
            .I(N__30123));
    Odrv4 I__5928 (
            .O(N__30134),
            .I(rand_data_3));
    Odrv12 I__5927 (
            .O(N__30131),
            .I(rand_data_3));
    LocalMux I__5926 (
            .O(N__30128),
            .I(rand_data_3));
    Odrv12 I__5925 (
            .O(N__30123),
            .I(rand_data_3));
    InMux I__5924 (
            .O(N__30114),
            .I(n16012));
    InMux I__5923 (
            .O(N__30111),
            .I(N__30106));
    InMux I__5922 (
            .O(N__30110),
            .I(N__30101));
    InMux I__5921 (
            .O(N__30109),
            .I(N__30098));
    LocalMux I__5920 (
            .O(N__30106),
            .I(N__30095));
    InMux I__5919 (
            .O(N__30105),
            .I(N__30092));
    InMux I__5918 (
            .O(N__30104),
            .I(N__30089));
    LocalMux I__5917 (
            .O(N__30101),
            .I(N__30083));
    LocalMux I__5916 (
            .O(N__30098),
            .I(N__30083));
    Span4Mux_h I__5915 (
            .O(N__30095),
            .I(N__30080));
    LocalMux I__5914 (
            .O(N__30092),
            .I(N__30077));
    LocalMux I__5913 (
            .O(N__30089),
            .I(N__30074));
    InMux I__5912 (
            .O(N__30088),
            .I(N__30071));
    Span4Mux_h I__5911 (
            .O(N__30083),
            .I(N__30066));
    Span4Mux_h I__5910 (
            .O(N__30080),
            .I(N__30066));
    Odrv12 I__5909 (
            .O(N__30077),
            .I(rand_data_4));
    Odrv4 I__5908 (
            .O(N__30074),
            .I(rand_data_4));
    LocalMux I__5907 (
            .O(N__30071),
            .I(rand_data_4));
    Odrv4 I__5906 (
            .O(N__30066),
            .I(rand_data_4));
    InMux I__5905 (
            .O(N__30057),
            .I(n16013));
    InMux I__5904 (
            .O(N__30054),
            .I(N__30050));
    InMux I__5903 (
            .O(N__30053),
            .I(N__30046));
    LocalMux I__5902 (
            .O(N__30050),
            .I(N__30043));
    InMux I__5901 (
            .O(N__30049),
            .I(N__30040));
    LocalMux I__5900 (
            .O(N__30046),
            .I(N__30036));
    Span4Mux_h I__5899 (
            .O(N__30043),
            .I(N__30033));
    LocalMux I__5898 (
            .O(N__30040),
            .I(N__30028));
    InMux I__5897 (
            .O(N__30039),
            .I(N__30025));
    Span4Mux_h I__5896 (
            .O(N__30036),
            .I(N__30022));
    Span4Mux_h I__5895 (
            .O(N__30033),
            .I(N__30019));
    InMux I__5894 (
            .O(N__30032),
            .I(N__30016));
    InMux I__5893 (
            .O(N__30031),
            .I(N__30013));
    Span4Mux_h I__5892 (
            .O(N__30028),
            .I(N__30006));
    LocalMux I__5891 (
            .O(N__30025),
            .I(N__30006));
    Span4Mux_h I__5890 (
            .O(N__30022),
            .I(N__30006));
    Odrv4 I__5889 (
            .O(N__30019),
            .I(rand_data_5));
    LocalMux I__5888 (
            .O(N__30016),
            .I(rand_data_5));
    LocalMux I__5887 (
            .O(N__30013),
            .I(rand_data_5));
    Odrv4 I__5886 (
            .O(N__30006),
            .I(rand_data_5));
    InMux I__5885 (
            .O(N__29997),
            .I(n16014));
    InMux I__5884 (
            .O(N__29994),
            .I(N__29988));
    InMux I__5883 (
            .O(N__29993),
            .I(N__29985));
    InMux I__5882 (
            .O(N__29992),
            .I(N__29982));
    InMux I__5881 (
            .O(N__29991),
            .I(N__29979));
    LocalMux I__5880 (
            .O(N__29988),
            .I(N__29976));
    LocalMux I__5879 (
            .O(N__29985),
            .I(N__29973));
    LocalMux I__5878 (
            .O(N__29982),
            .I(N__29970));
    LocalMux I__5877 (
            .O(N__29979),
            .I(N__29967));
    Span4Mux_h I__5876 (
            .O(N__29976),
            .I(N__29962));
    Span4Mux_h I__5875 (
            .O(N__29973),
            .I(N__29959));
    Span4Mux_v I__5874 (
            .O(N__29970),
            .I(N__29954));
    Span4Mux_h I__5873 (
            .O(N__29967),
            .I(N__29954));
    InMux I__5872 (
            .O(N__29966),
            .I(N__29951));
    InMux I__5871 (
            .O(N__29965),
            .I(N__29948));
    Span4Mux_h I__5870 (
            .O(N__29962),
            .I(N__29945));
    Odrv4 I__5869 (
            .O(N__29959),
            .I(rand_data_6));
    Odrv4 I__5868 (
            .O(N__29954),
            .I(rand_data_6));
    LocalMux I__5867 (
            .O(N__29951),
            .I(rand_data_6));
    LocalMux I__5866 (
            .O(N__29948),
            .I(rand_data_6));
    Odrv4 I__5865 (
            .O(N__29945),
            .I(rand_data_6));
    InMux I__5864 (
            .O(N__29934),
            .I(n16015));
    InMux I__5863 (
            .O(N__29931),
            .I(N__29926));
    InMux I__5862 (
            .O(N__29930),
            .I(N__29923));
    InMux I__5861 (
            .O(N__29929),
            .I(N__29920));
    LocalMux I__5860 (
            .O(N__29926),
            .I(N__29917));
    LocalMux I__5859 (
            .O(N__29923),
            .I(N__29913));
    LocalMux I__5858 (
            .O(N__29920),
            .I(N__29907));
    Span4Mux_v I__5857 (
            .O(N__29917),
            .I(N__29907));
    InMux I__5856 (
            .O(N__29916),
            .I(N__29904));
    Span4Mux_h I__5855 (
            .O(N__29913),
            .I(N__29900));
    InMux I__5854 (
            .O(N__29912),
            .I(N__29897));
    Span4Mux_h I__5853 (
            .O(N__29907),
            .I(N__29892));
    LocalMux I__5852 (
            .O(N__29904),
            .I(N__29892));
    InMux I__5851 (
            .O(N__29903),
            .I(N__29889));
    Span4Mux_h I__5850 (
            .O(N__29900),
            .I(N__29886));
    LocalMux I__5849 (
            .O(N__29897),
            .I(rand_data_7));
    Odrv4 I__5848 (
            .O(N__29892),
            .I(rand_data_7));
    LocalMux I__5847 (
            .O(N__29889),
            .I(rand_data_7));
    Odrv4 I__5846 (
            .O(N__29886),
            .I(rand_data_7));
    InMux I__5845 (
            .O(N__29877),
            .I(n16016));
    InMux I__5844 (
            .O(N__29874),
            .I(N__29869));
    InMux I__5843 (
            .O(N__29873),
            .I(N__29866));
    InMux I__5842 (
            .O(N__29872),
            .I(N__29863));
    LocalMux I__5841 (
            .O(N__29869),
            .I(N__29858));
    LocalMux I__5840 (
            .O(N__29866),
            .I(N__29855));
    LocalMux I__5839 (
            .O(N__29863),
            .I(N__29852));
    InMux I__5838 (
            .O(N__29862),
            .I(N__29847));
    InMux I__5837 (
            .O(N__29861),
            .I(N__29847));
    Span4Mux_h I__5836 (
            .O(N__29858),
            .I(N__29843));
    Span4Mux_h I__5835 (
            .O(N__29855),
            .I(N__29840));
    Span4Mux_h I__5834 (
            .O(N__29852),
            .I(N__29835));
    LocalMux I__5833 (
            .O(N__29847),
            .I(N__29835));
    InMux I__5832 (
            .O(N__29846),
            .I(N__29832));
    Span4Mux_h I__5831 (
            .O(N__29843),
            .I(N__29827));
    Span4Mux_h I__5830 (
            .O(N__29840),
            .I(N__29827));
    Odrv4 I__5829 (
            .O(N__29835),
            .I(rand_data_8));
    LocalMux I__5828 (
            .O(N__29832),
            .I(rand_data_8));
    Odrv4 I__5827 (
            .O(N__29827),
            .I(rand_data_8));
    InMux I__5826 (
            .O(N__29820),
            .I(bfn_10_26_0_));
    InMux I__5825 (
            .O(N__29817),
            .I(N__29813));
    InMux I__5824 (
            .O(N__29816),
            .I(N__29807));
    LocalMux I__5823 (
            .O(N__29813),
            .I(N__29804));
    InMux I__5822 (
            .O(N__29812),
            .I(N__29799));
    InMux I__5821 (
            .O(N__29811),
            .I(N__29799));
    InMux I__5820 (
            .O(N__29810),
            .I(N__29796));
    LocalMux I__5819 (
            .O(N__29807),
            .I(N__29793));
    Span4Mux_v I__5818 (
            .O(N__29804),
            .I(N__29790));
    LocalMux I__5817 (
            .O(N__29799),
            .I(N__29787));
    LocalMux I__5816 (
            .O(N__29796),
            .I(N__29784));
    Span4Mux_v I__5815 (
            .O(N__29793),
            .I(N__29780));
    Span4Mux_h I__5814 (
            .O(N__29790),
            .I(N__29775));
    Span4Mux_v I__5813 (
            .O(N__29787),
            .I(N__29775));
    Sp12to4 I__5812 (
            .O(N__29784),
            .I(N__29772));
    InMux I__5811 (
            .O(N__29783),
            .I(N__29769));
    Span4Mux_h I__5810 (
            .O(N__29780),
            .I(N__29766));
    Odrv4 I__5809 (
            .O(N__29775),
            .I(rand_data_9));
    Odrv12 I__5808 (
            .O(N__29772),
            .I(rand_data_9));
    LocalMux I__5807 (
            .O(N__29769),
            .I(rand_data_9));
    Odrv4 I__5806 (
            .O(N__29766),
            .I(rand_data_9));
    InMux I__5805 (
            .O(N__29757),
            .I(N__29754));
    LocalMux I__5804 (
            .O(N__29754),
            .I(N__29750));
    CascadeMux I__5803 (
            .O(N__29753),
            .I(N__29747));
    Span4Mux_v I__5802 (
            .O(N__29750),
            .I(N__29744));
    InMux I__5801 (
            .O(N__29747),
            .I(N__29741));
    Odrv4 I__5800 (
            .O(N__29744),
            .I(rand_setpoint_9));
    LocalMux I__5799 (
            .O(N__29741),
            .I(rand_setpoint_9));
    InMux I__5798 (
            .O(N__29736),
            .I(n16018));
    InMux I__5797 (
            .O(N__29733),
            .I(N__29727));
    InMux I__5796 (
            .O(N__29732),
            .I(N__29724));
    InMux I__5795 (
            .O(N__29731),
            .I(N__29719));
    InMux I__5794 (
            .O(N__29730),
            .I(N__29719));
    LocalMux I__5793 (
            .O(N__29727),
            .I(data_in_3_4));
    LocalMux I__5792 (
            .O(N__29724),
            .I(data_in_3_4));
    LocalMux I__5791 (
            .O(N__29719),
            .I(data_in_3_4));
    InMux I__5790 (
            .O(N__29712),
            .I(N__29707));
    InMux I__5789 (
            .O(N__29711),
            .I(N__29704));
    InMux I__5788 (
            .O(N__29710),
            .I(N__29701));
    LocalMux I__5787 (
            .O(N__29707),
            .I(N__29698));
    LocalMux I__5786 (
            .O(N__29704),
            .I(N__29695));
    LocalMux I__5785 (
            .O(N__29701),
            .I(N__29692));
    Span4Mux_h I__5784 (
            .O(N__29698),
            .I(N__29689));
    Span4Mux_v I__5783 (
            .O(N__29695),
            .I(N__29686));
    Span4Mux_h I__5782 (
            .O(N__29692),
            .I(N__29683));
    Span4Mux_v I__5781 (
            .O(N__29689),
            .I(N__29680));
    Span4Mux_v I__5780 (
            .O(N__29686),
            .I(N__29676));
    Span4Mux_v I__5779 (
            .O(N__29683),
            .I(N__29673));
    Span4Mux_v I__5778 (
            .O(N__29680),
            .I(N__29670));
    InMux I__5777 (
            .O(N__29679),
            .I(N__29667));
    Span4Mux_h I__5776 (
            .O(N__29676),
            .I(N__29662));
    Span4Mux_v I__5775 (
            .O(N__29673),
            .I(N__29662));
    Odrv4 I__5774 (
            .O(N__29670),
            .I(data_in_1_6));
    LocalMux I__5773 (
            .O(N__29667),
            .I(data_in_1_6));
    Odrv4 I__5772 (
            .O(N__29662),
            .I(data_in_1_6));
    CascadeMux I__5771 (
            .O(N__29655),
            .I(N__29652));
    InMux I__5770 (
            .O(N__29652),
            .I(N__29648));
    InMux I__5769 (
            .O(N__29651),
            .I(N__29643));
    LocalMux I__5768 (
            .O(N__29648),
            .I(N__29640));
    InMux I__5767 (
            .O(N__29647),
            .I(N__29637));
    InMux I__5766 (
            .O(N__29646),
            .I(N__29634));
    LocalMux I__5765 (
            .O(N__29643),
            .I(N__29627));
    Span4Mux_v I__5764 (
            .O(N__29640),
            .I(N__29627));
    LocalMux I__5763 (
            .O(N__29637),
            .I(N__29627));
    LocalMux I__5762 (
            .O(N__29634),
            .I(data_in_3_5));
    Odrv4 I__5761 (
            .O(N__29627),
            .I(data_in_3_5));
    InMux I__5760 (
            .O(N__29622),
            .I(N__29619));
    LocalMux I__5759 (
            .O(N__29619),
            .I(\c0.n17402 ));
    InMux I__5758 (
            .O(N__29616),
            .I(N__29613));
    LocalMux I__5757 (
            .O(N__29613),
            .I(N__29610));
    Span4Mux_h I__5756 (
            .O(N__29610),
            .I(N__29605));
    InMux I__5755 (
            .O(N__29609),
            .I(N__29602));
    InMux I__5754 (
            .O(N__29608),
            .I(N__29599));
    Span4Mux_v I__5753 (
            .O(N__29605),
            .I(N__29596));
    LocalMux I__5752 (
            .O(N__29602),
            .I(N__29593));
    LocalMux I__5751 (
            .O(N__29599),
            .I(\c0.FRAME_MATCHER_state_20 ));
    Odrv4 I__5750 (
            .O(N__29596),
            .I(\c0.FRAME_MATCHER_state_20 ));
    Odrv12 I__5749 (
            .O(N__29593),
            .I(\c0.FRAME_MATCHER_state_20 ));
    SRMux I__5748 (
            .O(N__29586),
            .I(N__29583));
    LocalMux I__5747 (
            .O(N__29583),
            .I(N__29580));
    Span4Mux_v I__5746 (
            .O(N__29580),
            .I(N__29577));
    Span4Mux_v I__5745 (
            .O(N__29577),
            .I(N__29574));
    Odrv4 I__5744 (
            .O(N__29574),
            .I(\c0.n8_adj_2327 ));
    CascadeMux I__5743 (
            .O(N__29571),
            .I(N__29568));
    InMux I__5742 (
            .O(N__29568),
            .I(N__29565));
    LocalMux I__5741 (
            .O(N__29565),
            .I(N__29561));
    InMux I__5740 (
            .O(N__29564),
            .I(N__29555));
    Span4Mux_v I__5739 (
            .O(N__29561),
            .I(N__29552));
    InMux I__5738 (
            .O(N__29560),
            .I(N__29549));
    InMux I__5737 (
            .O(N__29559),
            .I(N__29546));
    InMux I__5736 (
            .O(N__29558),
            .I(N__29543));
    LocalMux I__5735 (
            .O(N__29555),
            .I(N__29539));
    Span4Mux_h I__5734 (
            .O(N__29552),
            .I(N__29534));
    LocalMux I__5733 (
            .O(N__29549),
            .I(N__29534));
    LocalMux I__5732 (
            .O(N__29546),
            .I(N__29529));
    LocalMux I__5731 (
            .O(N__29543),
            .I(N__29529));
    InMux I__5730 (
            .O(N__29542),
            .I(N__29526));
    Span4Mux_v I__5729 (
            .O(N__29539),
            .I(N__29523));
    Span4Mux_h I__5728 (
            .O(N__29534),
            .I(N__29520));
    Span4Mux_h I__5727 (
            .O(N__29529),
            .I(N__29517));
    LocalMux I__5726 (
            .O(N__29526),
            .I(\c0.FRAME_MATCHER_i_31 ));
    Odrv4 I__5725 (
            .O(N__29523),
            .I(\c0.FRAME_MATCHER_i_31 ));
    Odrv4 I__5724 (
            .O(N__29520),
            .I(\c0.FRAME_MATCHER_i_31 ));
    Odrv4 I__5723 (
            .O(N__29517),
            .I(\c0.FRAME_MATCHER_i_31 ));
    InMux I__5722 (
            .O(N__29508),
            .I(N__29505));
    LocalMux I__5721 (
            .O(N__29505),
            .I(N__29502));
    Span4Mux_v I__5720 (
            .O(N__29502),
            .I(N__29499));
    Odrv4 I__5719 (
            .O(N__29499),
            .I(\c0.n10161 ));
    CascadeMux I__5718 (
            .O(N__29496),
            .I(n2061_cascade_));
    InMux I__5717 (
            .O(N__29493),
            .I(N__29490));
    LocalMux I__5716 (
            .O(N__29490),
            .I(\c0.n47_adj_2347 ));
    CascadeMux I__5715 (
            .O(N__29487),
            .I(\c0.n9334_cascade_ ));
    InMux I__5714 (
            .O(N__29484),
            .I(N__29481));
    LocalMux I__5713 (
            .O(N__29481),
            .I(\c0.n4 ));
    CascadeMux I__5712 (
            .O(N__29478),
            .I(\c0.n15821_cascade_ ));
    SRMux I__5711 (
            .O(N__29475),
            .I(N__29472));
    LocalMux I__5710 (
            .O(N__29472),
            .I(N__29469));
    Span4Mux_h I__5709 (
            .O(N__29469),
            .I(N__29466));
    Span4Mux_h I__5708 (
            .O(N__29466),
            .I(N__29463));
    Odrv4 I__5707 (
            .O(N__29463),
            .I(\c0.n8_adj_2335 ));
    InMux I__5706 (
            .O(N__29460),
            .I(N__29455));
    InMux I__5705 (
            .O(N__29459),
            .I(N__29450));
    InMux I__5704 (
            .O(N__29458),
            .I(N__29447));
    LocalMux I__5703 (
            .O(N__29455),
            .I(N__29444));
    InMux I__5702 (
            .O(N__29454),
            .I(N__29441));
    InMux I__5701 (
            .O(N__29453),
            .I(N__29438));
    LocalMux I__5700 (
            .O(N__29450),
            .I(N__29435));
    LocalMux I__5699 (
            .O(N__29447),
            .I(N__29432));
    Span4Mux_h I__5698 (
            .O(N__29444),
            .I(N__29428));
    LocalMux I__5697 (
            .O(N__29441),
            .I(N__29425));
    LocalMux I__5696 (
            .O(N__29438),
            .I(N__29420));
    Span4Mux_v I__5695 (
            .O(N__29435),
            .I(N__29420));
    Span12Mux_h I__5694 (
            .O(N__29432),
            .I(N__29417));
    InMux I__5693 (
            .O(N__29431),
            .I(N__29414));
    Span4Mux_h I__5692 (
            .O(N__29428),
            .I(N__29411));
    Odrv4 I__5691 (
            .O(N__29425),
            .I(rand_data_0));
    Odrv4 I__5690 (
            .O(N__29420),
            .I(rand_data_0));
    Odrv12 I__5689 (
            .O(N__29417),
            .I(rand_data_0));
    LocalMux I__5688 (
            .O(N__29414),
            .I(rand_data_0));
    Odrv4 I__5687 (
            .O(N__29411),
            .I(rand_data_0));
    CascadeMux I__5686 (
            .O(N__29400),
            .I(n63_cascade_));
    InMux I__5685 (
            .O(N__29397),
            .I(N__29394));
    LocalMux I__5684 (
            .O(N__29394),
            .I(N__29388));
    InMux I__5683 (
            .O(N__29393),
            .I(N__29381));
    InMux I__5682 (
            .O(N__29392),
            .I(N__29381));
    InMux I__5681 (
            .O(N__29391),
            .I(N__29381));
    Odrv4 I__5680 (
            .O(N__29388),
            .I(data_in_2_7));
    LocalMux I__5679 (
            .O(N__29381),
            .I(data_in_2_7));
    CascadeMux I__5678 (
            .O(N__29376),
            .I(N__29372));
    InMux I__5677 (
            .O(N__29375),
            .I(N__29369));
    InMux I__5676 (
            .O(N__29372),
            .I(N__29366));
    LocalMux I__5675 (
            .O(N__29369),
            .I(N__29361));
    LocalMux I__5674 (
            .O(N__29366),
            .I(N__29361));
    Span4Mux_v I__5673 (
            .O(N__29361),
            .I(N__29358));
    Odrv4 I__5672 (
            .O(N__29358),
            .I(\c0.n10141 ));
    InMux I__5671 (
            .O(N__29355),
            .I(N__29352));
    LocalMux I__5670 (
            .O(N__29352),
            .I(\c0.n10027 ));
    InMux I__5669 (
            .O(N__29349),
            .I(N__29346));
    LocalMux I__5668 (
            .O(N__29346),
            .I(N__29343));
    Span4Mux_v I__5667 (
            .O(N__29343),
            .I(N__29340));
    Odrv4 I__5666 (
            .O(N__29340),
            .I(\c0.n17_adj_2370 ));
    CascadeMux I__5665 (
            .O(N__29337),
            .I(\c0.n16_adj_2366_cascade_ ));
    InMux I__5664 (
            .O(N__29334),
            .I(N__29330));
    InMux I__5663 (
            .O(N__29333),
            .I(N__29325));
    LocalMux I__5662 (
            .O(N__29330),
            .I(N__29322));
    InMux I__5661 (
            .O(N__29329),
            .I(N__29317));
    InMux I__5660 (
            .O(N__29328),
            .I(N__29317));
    LocalMux I__5659 (
            .O(N__29325),
            .I(data_in_1_7));
    Odrv12 I__5658 (
            .O(N__29322),
            .I(data_in_1_7));
    LocalMux I__5657 (
            .O(N__29317),
            .I(data_in_1_7));
    CascadeMux I__5656 (
            .O(N__29310),
            .I(n9378_cascade_));
    CascadeMux I__5655 (
            .O(N__29307),
            .I(\c0.n47_adj_2347_cascade_ ));
    CascadeMux I__5654 (
            .O(N__29304),
            .I(\c0.n13146_cascade_ ));
    CascadeMux I__5653 (
            .O(N__29301),
            .I(N__29297));
    CascadeMux I__5652 (
            .O(N__29300),
            .I(N__29294));
    InMux I__5651 (
            .O(N__29297),
            .I(N__29291));
    InMux I__5650 (
            .O(N__29294),
            .I(N__29288));
    LocalMux I__5649 (
            .O(N__29291),
            .I(N__29285));
    LocalMux I__5648 (
            .O(N__29288),
            .I(\c0.data_in_frame_3_4 ));
    Odrv4 I__5647 (
            .O(N__29285),
            .I(\c0.data_in_frame_3_4 ));
    InMux I__5646 (
            .O(N__29280),
            .I(N__29275));
    InMux I__5645 (
            .O(N__29279),
            .I(N__29270));
    InMux I__5644 (
            .O(N__29278),
            .I(N__29270));
    LocalMux I__5643 (
            .O(N__29275),
            .I(data_in_0_1));
    LocalMux I__5642 (
            .O(N__29270),
            .I(data_in_0_1));
    CascadeMux I__5641 (
            .O(N__29265),
            .I(\c0.n7_adj_2384_cascade_ ));
    SRMux I__5640 (
            .O(N__29262),
            .I(N__29259));
    LocalMux I__5639 (
            .O(N__29259),
            .I(N__29256));
    Odrv4 I__5638 (
            .O(N__29256),
            .I(\c0.n6_adj_2336 ));
    InMux I__5637 (
            .O(N__29253),
            .I(N__29249));
    InMux I__5636 (
            .O(N__29252),
            .I(N__29246));
    LocalMux I__5635 (
            .O(N__29249),
            .I(\c0.n10136 ));
    LocalMux I__5634 (
            .O(N__29246),
            .I(\c0.n10136 ));
    InMux I__5633 (
            .O(N__29241),
            .I(N__29237));
    CascadeMux I__5632 (
            .O(N__29240),
            .I(N__29234));
    LocalMux I__5631 (
            .O(N__29237),
            .I(N__29229));
    InMux I__5630 (
            .O(N__29234),
            .I(N__29226));
    InMux I__5629 (
            .O(N__29233),
            .I(N__29221));
    InMux I__5628 (
            .O(N__29232),
            .I(N__29221));
    Odrv12 I__5627 (
            .O(N__29229),
            .I(data_in_1_4));
    LocalMux I__5626 (
            .O(N__29226),
            .I(data_in_1_4));
    LocalMux I__5625 (
            .O(N__29221),
            .I(data_in_1_4));
    InMux I__5624 (
            .O(N__29214),
            .I(N__29206));
    InMux I__5623 (
            .O(N__29213),
            .I(N__29206));
    InMux I__5622 (
            .O(N__29212),
            .I(N__29203));
    InMux I__5621 (
            .O(N__29211),
            .I(N__29200));
    LocalMux I__5620 (
            .O(N__29206),
            .I(data_in_2_3));
    LocalMux I__5619 (
            .O(N__29203),
            .I(data_in_2_3));
    LocalMux I__5618 (
            .O(N__29200),
            .I(data_in_2_3));
    CascadeMux I__5617 (
            .O(N__29193),
            .I(\c0.n16_adj_2361_cascade_ ));
    InMux I__5616 (
            .O(N__29190),
            .I(N__29187));
    LocalMux I__5615 (
            .O(N__29187),
            .I(\c0.n17_adj_2362 ));
    CascadeMux I__5614 (
            .O(N__29184),
            .I(n17075_cascade_));
    InMux I__5613 (
            .O(N__29181),
            .I(N__29177));
    InMux I__5612 (
            .O(N__29180),
            .I(N__29172));
    LocalMux I__5611 (
            .O(N__29177),
            .I(N__29169));
    InMux I__5610 (
            .O(N__29176),
            .I(N__29166));
    InMux I__5609 (
            .O(N__29175),
            .I(N__29163));
    LocalMux I__5608 (
            .O(N__29172),
            .I(data_in_2_5));
    Odrv12 I__5607 (
            .O(N__29169),
            .I(data_in_2_5));
    LocalMux I__5606 (
            .O(N__29166),
            .I(data_in_2_5));
    LocalMux I__5605 (
            .O(N__29163),
            .I(data_in_2_5));
    CascadeMux I__5604 (
            .O(N__29154),
            .I(N__29150));
    InMux I__5603 (
            .O(N__29153),
            .I(N__29144));
    InMux I__5602 (
            .O(N__29150),
            .I(N__29144));
    InMux I__5601 (
            .O(N__29149),
            .I(N__29141));
    LocalMux I__5600 (
            .O(N__29144),
            .I(N__29135));
    LocalMux I__5599 (
            .O(N__29141),
            .I(N__29135));
    InMux I__5598 (
            .O(N__29140),
            .I(N__29132));
    Span4Mux_v I__5597 (
            .O(N__29135),
            .I(N__29129));
    LocalMux I__5596 (
            .O(N__29132),
            .I(data_in_2_0));
    Odrv4 I__5595 (
            .O(N__29129),
            .I(data_in_2_0));
    CascadeMux I__5594 (
            .O(N__29124),
            .I(\c0.n17400_cascade_ ));
    CascadeMux I__5593 (
            .O(N__29121),
            .I(\c0.n8_adj_2359_cascade_ ));
    InMux I__5592 (
            .O(N__29118),
            .I(N__29115));
    LocalMux I__5591 (
            .O(N__29115),
            .I(\c0.n13450 ));
    CascadeMux I__5590 (
            .O(N__29112),
            .I(\c0.n15_adj_2310_cascade_ ));
    InMux I__5589 (
            .O(N__29109),
            .I(N__29105));
    InMux I__5588 (
            .O(N__29108),
            .I(N__29102));
    LocalMux I__5587 (
            .O(N__29105),
            .I(\c0.data_in_frame_3_3 ));
    LocalMux I__5586 (
            .O(N__29102),
            .I(\c0.data_in_frame_3_3 ));
    InMux I__5585 (
            .O(N__29097),
            .I(N__29094));
    LocalMux I__5584 (
            .O(N__29094),
            .I(\c0.n17659 ));
    CascadeMux I__5583 (
            .O(N__29091),
            .I(\c0.n11867_cascade_ ));
    SRMux I__5582 (
            .O(N__29088),
            .I(N__29085));
    LocalMux I__5581 (
            .O(N__29085),
            .I(N__29082));
    Odrv4 I__5580 (
            .O(N__29082),
            .I(\c0.n4_adj_2187 ));
    SRMux I__5579 (
            .O(N__29079),
            .I(N__29076));
    LocalMux I__5578 (
            .O(N__29076),
            .I(\c0.n4_adj_2152 ));
    CascadeMux I__5577 (
            .O(N__29073),
            .I(N__29070));
    InMux I__5576 (
            .O(N__29070),
            .I(N__29067));
    LocalMux I__5575 (
            .O(N__29067),
            .I(N__29063));
    CascadeMux I__5574 (
            .O(N__29066),
            .I(N__29060));
    Span4Mux_v I__5573 (
            .O(N__29063),
            .I(N__29044));
    InMux I__5572 (
            .O(N__29060),
            .I(N__29041));
    InMux I__5571 (
            .O(N__29059),
            .I(N__29036));
    InMux I__5570 (
            .O(N__29058),
            .I(N__29036));
    InMux I__5569 (
            .O(N__29057),
            .I(N__29033));
    InMux I__5568 (
            .O(N__29056),
            .I(N__29028));
    InMux I__5567 (
            .O(N__29055),
            .I(N__29028));
    InMux I__5566 (
            .O(N__29054),
            .I(N__29025));
    InMux I__5565 (
            .O(N__29053),
            .I(N__29019));
    InMux I__5564 (
            .O(N__29052),
            .I(N__29014));
    InMux I__5563 (
            .O(N__29051),
            .I(N__29014));
    InMux I__5562 (
            .O(N__29050),
            .I(N__29009));
    InMux I__5561 (
            .O(N__29049),
            .I(N__29009));
    InMux I__5560 (
            .O(N__29048),
            .I(N__29000));
    InMux I__5559 (
            .O(N__29047),
            .I(N__28994));
    Span4Mux_h I__5558 (
            .O(N__29044),
            .I(N__28989));
    LocalMux I__5557 (
            .O(N__29041),
            .I(N__28989));
    LocalMux I__5556 (
            .O(N__29036),
            .I(N__28986));
    LocalMux I__5555 (
            .O(N__29033),
            .I(N__28981));
    LocalMux I__5554 (
            .O(N__29028),
            .I(N__28981));
    LocalMux I__5553 (
            .O(N__29025),
            .I(N__28978));
    InMux I__5552 (
            .O(N__29024),
            .I(N__28973));
    InMux I__5551 (
            .O(N__29023),
            .I(N__28973));
    CascadeMux I__5550 (
            .O(N__29022),
            .I(N__28963));
    LocalMux I__5549 (
            .O(N__29019),
            .I(N__28954));
    LocalMux I__5548 (
            .O(N__29014),
            .I(N__28954));
    LocalMux I__5547 (
            .O(N__29009),
            .I(N__28951));
    InMux I__5546 (
            .O(N__29008),
            .I(N__28944));
    InMux I__5545 (
            .O(N__29007),
            .I(N__28944));
    InMux I__5544 (
            .O(N__29006),
            .I(N__28944));
    InMux I__5543 (
            .O(N__29005),
            .I(N__28939));
    InMux I__5542 (
            .O(N__29004),
            .I(N__28939));
    InMux I__5541 (
            .O(N__29003),
            .I(N__28935));
    LocalMux I__5540 (
            .O(N__29000),
            .I(N__28929));
    InMux I__5539 (
            .O(N__28999),
            .I(N__28926));
    InMux I__5538 (
            .O(N__28998),
            .I(N__28920));
    InMux I__5537 (
            .O(N__28997),
            .I(N__28917));
    LocalMux I__5536 (
            .O(N__28994),
            .I(N__28914));
    Span4Mux_v I__5535 (
            .O(N__28989),
            .I(N__28911));
    Span4Mux_s2_h I__5534 (
            .O(N__28986),
            .I(N__28902));
    Span4Mux_v I__5533 (
            .O(N__28981),
            .I(N__28902));
    Span4Mux_v I__5532 (
            .O(N__28978),
            .I(N__28902));
    LocalMux I__5531 (
            .O(N__28973),
            .I(N__28902));
    InMux I__5530 (
            .O(N__28972),
            .I(N__28896));
    InMux I__5529 (
            .O(N__28971),
            .I(N__28896));
    InMux I__5528 (
            .O(N__28970),
            .I(N__28893));
    InMux I__5527 (
            .O(N__28969),
            .I(N__28888));
    InMux I__5526 (
            .O(N__28968),
            .I(N__28881));
    InMux I__5525 (
            .O(N__28967),
            .I(N__28881));
    InMux I__5524 (
            .O(N__28966),
            .I(N__28881));
    InMux I__5523 (
            .O(N__28963),
            .I(N__28878));
    InMux I__5522 (
            .O(N__28962),
            .I(N__28873));
    InMux I__5521 (
            .O(N__28961),
            .I(N__28873));
    InMux I__5520 (
            .O(N__28960),
            .I(N__28870));
    InMux I__5519 (
            .O(N__28959),
            .I(N__28867));
    Span4Mux_v I__5518 (
            .O(N__28954),
            .I(N__28862));
    Span4Mux_h I__5517 (
            .O(N__28951),
            .I(N__28862));
    LocalMux I__5516 (
            .O(N__28944),
            .I(N__28857));
    LocalMux I__5515 (
            .O(N__28939),
            .I(N__28857));
    InMux I__5514 (
            .O(N__28938),
            .I(N__28854));
    LocalMux I__5513 (
            .O(N__28935),
            .I(N__28851));
    InMux I__5512 (
            .O(N__28934),
            .I(N__28846));
    InMux I__5511 (
            .O(N__28933),
            .I(N__28846));
    InMux I__5510 (
            .O(N__28932),
            .I(N__28843));
    Span4Mux_s2_h I__5509 (
            .O(N__28929),
            .I(N__28838));
    LocalMux I__5508 (
            .O(N__28926),
            .I(N__28838));
    InMux I__5507 (
            .O(N__28925),
            .I(N__28831));
    InMux I__5506 (
            .O(N__28924),
            .I(N__28831));
    InMux I__5505 (
            .O(N__28923),
            .I(N__28831));
    LocalMux I__5504 (
            .O(N__28920),
            .I(N__28826));
    LocalMux I__5503 (
            .O(N__28917),
            .I(N__28826));
    Span4Mux_v I__5502 (
            .O(N__28914),
            .I(N__28819));
    Span4Mux_h I__5501 (
            .O(N__28911),
            .I(N__28819));
    Span4Mux_v I__5500 (
            .O(N__28902),
            .I(N__28819));
    InMux I__5499 (
            .O(N__28901),
            .I(N__28813));
    LocalMux I__5498 (
            .O(N__28896),
            .I(N__28808));
    LocalMux I__5497 (
            .O(N__28893),
            .I(N__28808));
    InMux I__5496 (
            .O(N__28892),
            .I(N__28803));
    InMux I__5495 (
            .O(N__28891),
            .I(N__28803));
    LocalMux I__5494 (
            .O(N__28888),
            .I(N__28794));
    LocalMux I__5493 (
            .O(N__28881),
            .I(N__28794));
    LocalMux I__5492 (
            .O(N__28878),
            .I(N__28794));
    LocalMux I__5491 (
            .O(N__28873),
            .I(N__28794));
    LocalMux I__5490 (
            .O(N__28870),
            .I(N__28791));
    LocalMux I__5489 (
            .O(N__28867),
            .I(N__28784));
    Span4Mux_v I__5488 (
            .O(N__28862),
            .I(N__28784));
    Span4Mux_h I__5487 (
            .O(N__28857),
            .I(N__28784));
    LocalMux I__5486 (
            .O(N__28854),
            .I(N__28776));
    Span4Mux_v I__5485 (
            .O(N__28851),
            .I(N__28776));
    LocalMux I__5484 (
            .O(N__28846),
            .I(N__28776));
    LocalMux I__5483 (
            .O(N__28843),
            .I(N__28773));
    Span4Mux_h I__5482 (
            .O(N__28838),
            .I(N__28764));
    LocalMux I__5481 (
            .O(N__28831),
            .I(N__28764));
    Span4Mux_v I__5480 (
            .O(N__28826),
            .I(N__28764));
    Span4Mux_h I__5479 (
            .O(N__28819),
            .I(N__28764));
    InMux I__5478 (
            .O(N__28818),
            .I(N__28757));
    InMux I__5477 (
            .O(N__28817),
            .I(N__28757));
    InMux I__5476 (
            .O(N__28816),
            .I(N__28757));
    LocalMux I__5475 (
            .O(N__28813),
            .I(N__28748));
    Span4Mux_v I__5474 (
            .O(N__28808),
            .I(N__28748));
    LocalMux I__5473 (
            .O(N__28803),
            .I(N__28748));
    Span4Mux_h I__5472 (
            .O(N__28794),
            .I(N__28748));
    Span4Mux_h I__5471 (
            .O(N__28791),
            .I(N__28743));
    Span4Mux_h I__5470 (
            .O(N__28784),
            .I(N__28743));
    InMux I__5469 (
            .O(N__28783),
            .I(N__28740));
    Span4Mux_h I__5468 (
            .O(N__28776),
            .I(N__28735));
    Span4Mux_h I__5467 (
            .O(N__28773),
            .I(N__28735));
    Span4Mux_h I__5466 (
            .O(N__28764),
            .I(N__28732));
    LocalMux I__5465 (
            .O(N__28757),
            .I(N__28725));
    Span4Mux_h I__5464 (
            .O(N__28748),
            .I(N__28725));
    Span4Mux_v I__5463 (
            .O(N__28743),
            .I(N__28725));
    LocalMux I__5462 (
            .O(N__28740),
            .I(\c0.byte_transmit_counter2_0 ));
    Odrv4 I__5461 (
            .O(N__28735),
            .I(\c0.byte_transmit_counter2_0 ));
    Odrv4 I__5460 (
            .O(N__28732),
            .I(\c0.byte_transmit_counter2_0 ));
    Odrv4 I__5459 (
            .O(N__28725),
            .I(\c0.byte_transmit_counter2_0 ));
    InMux I__5458 (
            .O(N__28716),
            .I(N__28713));
    LocalMux I__5457 (
            .O(N__28713),
            .I(N__28710));
    Span4Mux_h I__5456 (
            .O(N__28710),
            .I(N__28707));
    Span4Mux_h I__5455 (
            .O(N__28707),
            .I(N__28704));
    Odrv4 I__5454 (
            .O(N__28704),
            .I(\c0.n17761 ));
    InMux I__5453 (
            .O(N__28701),
            .I(N__28696));
    InMux I__5452 (
            .O(N__28700),
            .I(N__28689));
    InMux I__5451 (
            .O(N__28699),
            .I(N__28689));
    LocalMux I__5450 (
            .O(N__28696),
            .I(N__28686));
    InMux I__5449 (
            .O(N__28695),
            .I(N__28680));
    InMux I__5448 (
            .O(N__28694),
            .I(N__28677));
    LocalMux I__5447 (
            .O(N__28689),
            .I(N__28672));
    Span4Mux_v I__5446 (
            .O(N__28686),
            .I(N__28669));
    InMux I__5445 (
            .O(N__28685),
            .I(N__28664));
    InMux I__5444 (
            .O(N__28684),
            .I(N__28664));
    CascadeMux I__5443 (
            .O(N__28683),
            .I(N__28656));
    LocalMux I__5442 (
            .O(N__28680),
            .I(N__28642));
    LocalMux I__5441 (
            .O(N__28677),
            .I(N__28642));
    CascadeMux I__5440 (
            .O(N__28676),
            .I(N__28633));
    CascadeMux I__5439 (
            .O(N__28675),
            .I(N__28628));
    Span4Mux_v I__5438 (
            .O(N__28672),
            .I(N__28621));
    Span4Mux_h I__5437 (
            .O(N__28669),
            .I(N__28621));
    LocalMux I__5436 (
            .O(N__28664),
            .I(N__28621));
    InMux I__5435 (
            .O(N__28663),
            .I(N__28616));
    InMux I__5434 (
            .O(N__28662),
            .I(N__28616));
    CascadeMux I__5433 (
            .O(N__28661),
            .I(N__28607));
    InMux I__5432 (
            .O(N__28660),
            .I(N__28602));
    InMux I__5431 (
            .O(N__28659),
            .I(N__28602));
    InMux I__5430 (
            .O(N__28656),
            .I(N__28591));
    InMux I__5429 (
            .O(N__28655),
            .I(N__28591));
    CascadeMux I__5428 (
            .O(N__28654),
            .I(N__28586));
    InMux I__5427 (
            .O(N__28653),
            .I(N__28580));
    InMux I__5426 (
            .O(N__28652),
            .I(N__28580));
    InMux I__5425 (
            .O(N__28651),
            .I(N__28577));
    InMux I__5424 (
            .O(N__28650),
            .I(N__28572));
    InMux I__5423 (
            .O(N__28649),
            .I(N__28572));
    InMux I__5422 (
            .O(N__28648),
            .I(N__28567));
    InMux I__5421 (
            .O(N__28647),
            .I(N__28567));
    Span4Mux_h I__5420 (
            .O(N__28642),
            .I(N__28564));
    InMux I__5419 (
            .O(N__28641),
            .I(N__28561));
    InMux I__5418 (
            .O(N__28640),
            .I(N__28556));
    InMux I__5417 (
            .O(N__28639),
            .I(N__28556));
    InMux I__5416 (
            .O(N__28638),
            .I(N__28551));
    InMux I__5415 (
            .O(N__28637),
            .I(N__28551));
    InMux I__5414 (
            .O(N__28636),
            .I(N__28539));
    InMux I__5413 (
            .O(N__28633),
            .I(N__28539));
    InMux I__5412 (
            .O(N__28632),
            .I(N__28539));
    InMux I__5411 (
            .O(N__28631),
            .I(N__28534));
    InMux I__5410 (
            .O(N__28628),
            .I(N__28534));
    Span4Mux_v I__5409 (
            .O(N__28621),
            .I(N__28531));
    LocalMux I__5408 (
            .O(N__28616),
            .I(N__28528));
    InMux I__5407 (
            .O(N__28615),
            .I(N__28523));
    InMux I__5406 (
            .O(N__28614),
            .I(N__28523));
    InMux I__5405 (
            .O(N__28613),
            .I(N__28520));
    InMux I__5404 (
            .O(N__28612),
            .I(N__28517));
    InMux I__5403 (
            .O(N__28611),
            .I(N__28510));
    InMux I__5402 (
            .O(N__28610),
            .I(N__28510));
    InMux I__5401 (
            .O(N__28607),
            .I(N__28510));
    LocalMux I__5400 (
            .O(N__28602),
            .I(N__28507));
    CascadeMux I__5399 (
            .O(N__28601),
            .I(N__28500));
    CascadeMux I__5398 (
            .O(N__28600),
            .I(N__28494));
    CascadeMux I__5397 (
            .O(N__28599),
            .I(N__28490));
    InMux I__5396 (
            .O(N__28598),
            .I(N__28487));
    CascadeMux I__5395 (
            .O(N__28597),
            .I(N__28484));
    InMux I__5394 (
            .O(N__28596),
            .I(N__28480));
    LocalMux I__5393 (
            .O(N__28591),
            .I(N__28477));
    InMux I__5392 (
            .O(N__28590),
            .I(N__28474));
    InMux I__5391 (
            .O(N__28589),
            .I(N__28469));
    InMux I__5390 (
            .O(N__28586),
            .I(N__28469));
    InMux I__5389 (
            .O(N__28585),
            .I(N__28466));
    LocalMux I__5388 (
            .O(N__28580),
            .I(N__28462));
    LocalMux I__5387 (
            .O(N__28577),
            .I(N__28455));
    LocalMux I__5386 (
            .O(N__28572),
            .I(N__28455));
    LocalMux I__5385 (
            .O(N__28567),
            .I(N__28455));
    Span4Mux_h I__5384 (
            .O(N__28564),
            .I(N__28450));
    LocalMux I__5383 (
            .O(N__28561),
            .I(N__28450));
    LocalMux I__5382 (
            .O(N__28556),
            .I(N__28442));
    LocalMux I__5381 (
            .O(N__28551),
            .I(N__28442));
    InMux I__5380 (
            .O(N__28550),
            .I(N__28431));
    InMux I__5379 (
            .O(N__28549),
            .I(N__28431));
    InMux I__5378 (
            .O(N__28548),
            .I(N__28431));
    InMux I__5377 (
            .O(N__28547),
            .I(N__28431));
    InMux I__5376 (
            .O(N__28546),
            .I(N__28431));
    LocalMux I__5375 (
            .O(N__28539),
            .I(N__28426));
    LocalMux I__5374 (
            .O(N__28534),
            .I(N__28426));
    IoSpan4Mux I__5373 (
            .O(N__28531),
            .I(N__28423));
    Span4Mux_v I__5372 (
            .O(N__28528),
            .I(N__28420));
    LocalMux I__5371 (
            .O(N__28523),
            .I(N__28411));
    LocalMux I__5370 (
            .O(N__28520),
            .I(N__28411));
    LocalMux I__5369 (
            .O(N__28517),
            .I(N__28411));
    LocalMux I__5368 (
            .O(N__28510),
            .I(N__28411));
    Span4Mux_v I__5367 (
            .O(N__28507),
            .I(N__28408));
    InMux I__5366 (
            .O(N__28506),
            .I(N__28401));
    InMux I__5365 (
            .O(N__28505),
            .I(N__28401));
    InMux I__5364 (
            .O(N__28504),
            .I(N__28401));
    InMux I__5363 (
            .O(N__28503),
            .I(N__28394));
    InMux I__5362 (
            .O(N__28500),
            .I(N__28394));
    InMux I__5361 (
            .O(N__28499),
            .I(N__28394));
    InMux I__5360 (
            .O(N__28498),
            .I(N__28387));
    InMux I__5359 (
            .O(N__28497),
            .I(N__28387));
    InMux I__5358 (
            .O(N__28494),
            .I(N__28387));
    InMux I__5357 (
            .O(N__28493),
            .I(N__28384));
    InMux I__5356 (
            .O(N__28490),
            .I(N__28381));
    LocalMux I__5355 (
            .O(N__28487),
            .I(N__28378));
    InMux I__5354 (
            .O(N__28484),
            .I(N__28373));
    InMux I__5353 (
            .O(N__28483),
            .I(N__28373));
    LocalMux I__5352 (
            .O(N__28480),
            .I(N__28368));
    Span4Mux_s3_h I__5351 (
            .O(N__28477),
            .I(N__28368));
    LocalMux I__5350 (
            .O(N__28474),
            .I(N__28363));
    LocalMux I__5349 (
            .O(N__28469),
            .I(N__28363));
    LocalMux I__5348 (
            .O(N__28466),
            .I(N__28357));
    InMux I__5347 (
            .O(N__28465),
            .I(N__28354));
    Span4Mux_h I__5346 (
            .O(N__28462),
            .I(N__28347));
    Span4Mux_v I__5345 (
            .O(N__28455),
            .I(N__28347));
    Span4Mux_v I__5344 (
            .O(N__28450),
            .I(N__28347));
    InMux I__5343 (
            .O(N__28449),
            .I(N__28340));
    InMux I__5342 (
            .O(N__28448),
            .I(N__28340));
    InMux I__5341 (
            .O(N__28447),
            .I(N__28340));
    Span4Mux_v I__5340 (
            .O(N__28442),
            .I(N__28329));
    LocalMux I__5339 (
            .O(N__28431),
            .I(N__28329));
    Span4Mux_v I__5338 (
            .O(N__28426),
            .I(N__28329));
    Span4Mux_s2_h I__5337 (
            .O(N__28423),
            .I(N__28329));
    Span4Mux_v I__5336 (
            .O(N__28420),
            .I(N__28329));
    Span4Mux_v I__5335 (
            .O(N__28411),
            .I(N__28314));
    Span4Mux_h I__5334 (
            .O(N__28408),
            .I(N__28314));
    LocalMux I__5333 (
            .O(N__28401),
            .I(N__28314));
    LocalMux I__5332 (
            .O(N__28394),
            .I(N__28314));
    LocalMux I__5331 (
            .O(N__28387),
            .I(N__28314));
    LocalMux I__5330 (
            .O(N__28384),
            .I(N__28314));
    LocalMux I__5329 (
            .O(N__28381),
            .I(N__28314));
    Span4Mux_v I__5328 (
            .O(N__28378),
            .I(N__28305));
    LocalMux I__5327 (
            .O(N__28373),
            .I(N__28305));
    Span4Mux_v I__5326 (
            .O(N__28368),
            .I(N__28305));
    Span4Mux_v I__5325 (
            .O(N__28363),
            .I(N__28305));
    InMux I__5324 (
            .O(N__28362),
            .I(N__28302));
    InMux I__5323 (
            .O(N__28361),
            .I(N__28299));
    InMux I__5322 (
            .O(N__28360),
            .I(N__28296));
    Span4Mux_h I__5321 (
            .O(N__28357),
            .I(N__28293));
    LocalMux I__5320 (
            .O(N__28354),
            .I(N__28288));
    Span4Mux_h I__5319 (
            .O(N__28347),
            .I(N__28288));
    LocalMux I__5318 (
            .O(N__28340),
            .I(N__28281));
    Span4Mux_h I__5317 (
            .O(N__28329),
            .I(N__28281));
    Span4Mux_v I__5316 (
            .O(N__28314),
            .I(N__28281));
    Span4Mux_h I__5315 (
            .O(N__28305),
            .I(N__28278));
    LocalMux I__5314 (
            .O(N__28302),
            .I(\c0.byte_transmit_counter2_1 ));
    LocalMux I__5313 (
            .O(N__28299),
            .I(\c0.byte_transmit_counter2_1 ));
    LocalMux I__5312 (
            .O(N__28296),
            .I(\c0.byte_transmit_counter2_1 ));
    Odrv4 I__5311 (
            .O(N__28293),
            .I(\c0.byte_transmit_counter2_1 ));
    Odrv4 I__5310 (
            .O(N__28288),
            .I(\c0.byte_transmit_counter2_1 ));
    Odrv4 I__5309 (
            .O(N__28281),
            .I(\c0.byte_transmit_counter2_1 ));
    Odrv4 I__5308 (
            .O(N__28278),
            .I(\c0.byte_transmit_counter2_1 ));
    SRMux I__5307 (
            .O(N__28263),
            .I(N__28260));
    LocalMux I__5306 (
            .O(N__28260),
            .I(\c0.n4_adj_2155 ));
    InMux I__5305 (
            .O(N__28257),
            .I(N__28251));
    InMux I__5304 (
            .O(N__28256),
            .I(N__28251));
    LocalMux I__5303 (
            .O(N__28251),
            .I(\c0.data_in_frame_3_6 ));
    InMux I__5302 (
            .O(N__28248),
            .I(N__28245));
    LocalMux I__5301 (
            .O(N__28245),
            .I(n7));
    InMux I__5300 (
            .O(N__28242),
            .I(n16059));
    InMux I__5299 (
            .O(N__28239),
            .I(N__28236));
    LocalMux I__5298 (
            .O(N__28236),
            .I(n6_adj_2429));
    InMux I__5297 (
            .O(N__28233),
            .I(n16060));
    InMux I__5296 (
            .O(N__28230),
            .I(n16061));
    InMux I__5295 (
            .O(N__28227),
            .I(n16062));
    InMux I__5294 (
            .O(N__28224),
            .I(n16063));
    InMux I__5293 (
            .O(N__28221),
            .I(bfn_9_32_0_));
    InMux I__5292 (
            .O(N__28218),
            .I(n16065));
    InMux I__5291 (
            .O(N__28215),
            .I(N__28212));
    LocalMux I__5290 (
            .O(N__28212),
            .I(\c0.n17711 ));
    InMux I__5289 (
            .O(N__28209),
            .I(N__28206));
    LocalMux I__5288 (
            .O(N__28206),
            .I(n15));
    InMux I__5287 (
            .O(N__28203),
            .I(n16051));
    InMux I__5286 (
            .O(N__28200),
            .I(N__28197));
    LocalMux I__5285 (
            .O(N__28197),
            .I(n14));
    InMux I__5284 (
            .O(N__28194),
            .I(n16052));
    InMux I__5283 (
            .O(N__28191),
            .I(N__28188));
    LocalMux I__5282 (
            .O(N__28188),
            .I(n13));
    InMux I__5281 (
            .O(N__28185),
            .I(n16053));
    InMux I__5280 (
            .O(N__28182),
            .I(N__28179));
    LocalMux I__5279 (
            .O(N__28179),
            .I(n12));
    InMux I__5278 (
            .O(N__28176),
            .I(n16054));
    InMux I__5277 (
            .O(N__28173),
            .I(N__28170));
    LocalMux I__5276 (
            .O(N__28170),
            .I(n11));
    InMux I__5275 (
            .O(N__28167),
            .I(n16055));
    InMux I__5274 (
            .O(N__28164),
            .I(N__28161));
    LocalMux I__5273 (
            .O(N__28161),
            .I(n10_adj_2420));
    InMux I__5272 (
            .O(N__28158),
            .I(bfn_9_31_0_));
    InMux I__5271 (
            .O(N__28155),
            .I(N__28152));
    LocalMux I__5270 (
            .O(N__28152),
            .I(n9_adj_2421));
    InMux I__5269 (
            .O(N__28149),
            .I(n16057));
    InMux I__5268 (
            .O(N__28146),
            .I(N__28143));
    LocalMux I__5267 (
            .O(N__28143),
            .I(n8_adj_2412));
    InMux I__5266 (
            .O(N__28140),
            .I(n16058));
    InMux I__5265 (
            .O(N__28137),
            .I(N__28134));
    LocalMux I__5264 (
            .O(N__28134),
            .I(n24));
    InMux I__5263 (
            .O(N__28131),
            .I(n16042));
    InMux I__5262 (
            .O(N__28128),
            .I(N__28125));
    LocalMux I__5261 (
            .O(N__28125),
            .I(n23_adj_2425));
    InMux I__5260 (
            .O(N__28122),
            .I(n16043));
    InMux I__5259 (
            .O(N__28119),
            .I(N__28116));
    LocalMux I__5258 (
            .O(N__28116),
            .I(n22_adj_2426));
    InMux I__5257 (
            .O(N__28113),
            .I(n16044));
    InMux I__5256 (
            .O(N__28110),
            .I(N__28107));
    LocalMux I__5255 (
            .O(N__28107),
            .I(n21));
    InMux I__5254 (
            .O(N__28104),
            .I(n16045));
    InMux I__5253 (
            .O(N__28101),
            .I(N__28098));
    LocalMux I__5252 (
            .O(N__28098),
            .I(n20));
    InMux I__5251 (
            .O(N__28095),
            .I(n16046));
    InMux I__5250 (
            .O(N__28092),
            .I(N__28089));
    LocalMux I__5249 (
            .O(N__28089),
            .I(n19));
    InMux I__5248 (
            .O(N__28086),
            .I(n16047));
    InMux I__5247 (
            .O(N__28083),
            .I(N__28080));
    LocalMux I__5246 (
            .O(N__28080),
            .I(n18));
    InMux I__5245 (
            .O(N__28077),
            .I(bfn_9_30_0_));
    InMux I__5244 (
            .O(N__28074),
            .I(N__28071));
    LocalMux I__5243 (
            .O(N__28071),
            .I(n17));
    InMux I__5242 (
            .O(N__28068),
            .I(n16049));
    InMux I__5241 (
            .O(N__28065),
            .I(N__28062));
    LocalMux I__5240 (
            .O(N__28062),
            .I(n16));
    InMux I__5239 (
            .O(N__28059),
            .I(n16050));
    InMux I__5238 (
            .O(N__28056),
            .I(N__28049));
    InMux I__5237 (
            .O(N__28055),
            .I(N__28049));
    InMux I__5236 (
            .O(N__28054),
            .I(N__28045));
    LocalMux I__5235 (
            .O(N__28049),
            .I(N__28042));
    InMux I__5234 (
            .O(N__28048),
            .I(N__28039));
    LocalMux I__5233 (
            .O(N__28045),
            .I(N__28034));
    Span12Mux_s5_v I__5232 (
            .O(N__28042),
            .I(N__28034));
    LocalMux I__5231 (
            .O(N__28039),
            .I(data_in_1_2));
    Odrv12 I__5230 (
            .O(N__28034),
            .I(data_in_1_2));
    InMux I__5229 (
            .O(N__28029),
            .I(N__28026));
    LocalMux I__5228 (
            .O(N__28026),
            .I(N__28023));
    Span4Mux_v I__5227 (
            .O(N__28023),
            .I(N__28020));
    Odrv4 I__5226 (
            .O(N__28020),
            .I(\c0.n17388 ));
    SRMux I__5225 (
            .O(N__28017),
            .I(N__28014));
    LocalMux I__5224 (
            .O(N__28014),
            .I(N__28011));
    Span4Mux_h I__5223 (
            .O(N__28011),
            .I(N__28008));
    Odrv4 I__5222 (
            .O(N__28008),
            .I(\c0.n3_adj_2272 ));
    CascadeMux I__5221 (
            .O(N__28005),
            .I(N__28002));
    InMux I__5220 (
            .O(N__28002),
            .I(N__27997));
    InMux I__5219 (
            .O(N__28001),
            .I(N__27993));
    InMux I__5218 (
            .O(N__28000),
            .I(N__27990));
    LocalMux I__5217 (
            .O(N__27997),
            .I(N__27987));
    InMux I__5216 (
            .O(N__27996),
            .I(N__27984));
    LocalMux I__5215 (
            .O(N__27993),
            .I(N__27979));
    LocalMux I__5214 (
            .O(N__27990),
            .I(N__27979));
    Span4Mux_h I__5213 (
            .O(N__27987),
            .I(N__27974));
    LocalMux I__5212 (
            .O(N__27984),
            .I(N__27974));
    Odrv4 I__5211 (
            .O(N__27979),
            .I(\c0.FRAME_MATCHER_i_10 ));
    Odrv4 I__5210 (
            .O(N__27974),
            .I(\c0.FRAME_MATCHER_i_10 ));
    InMux I__5209 (
            .O(N__27969),
            .I(N__27966));
    LocalMux I__5208 (
            .O(N__27966),
            .I(N__27963));
    Span4Mux_h I__5207 (
            .O(N__27963),
            .I(N__27960));
    Odrv4 I__5206 (
            .O(N__27960),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_10 ));
    SRMux I__5205 (
            .O(N__27957),
            .I(N__27954));
    LocalMux I__5204 (
            .O(N__27954),
            .I(N__27951));
    Span4Mux_s1_h I__5203 (
            .O(N__27951),
            .I(N__27948));
    Span4Mux_h I__5202 (
            .O(N__27948),
            .I(N__27945));
    Odrv4 I__5201 (
            .O(N__27945),
            .I(\c0.n3_adj_2264 ));
    CascadeMux I__5200 (
            .O(N__27942),
            .I(N__27938));
    CascadeMux I__5199 (
            .O(N__27941),
            .I(N__27934));
    InMux I__5198 (
            .O(N__27938),
            .I(N__27929));
    InMux I__5197 (
            .O(N__27937),
            .I(N__27929));
    InMux I__5196 (
            .O(N__27934),
            .I(N__27925));
    LocalMux I__5195 (
            .O(N__27929),
            .I(N__27922));
    InMux I__5194 (
            .O(N__27928),
            .I(N__27919));
    LocalMux I__5193 (
            .O(N__27925),
            .I(N__27916));
    Span4Mux_v I__5192 (
            .O(N__27922),
            .I(N__27911));
    LocalMux I__5191 (
            .O(N__27919),
            .I(N__27911));
    Span4Mux_v I__5190 (
            .O(N__27916),
            .I(N__27906));
    Span4Mux_h I__5189 (
            .O(N__27911),
            .I(N__27906));
    Span4Mux_h I__5188 (
            .O(N__27906),
            .I(N__27903));
    Odrv4 I__5187 (
            .O(N__27903),
            .I(\c0.FRAME_MATCHER_i_14 ));
    InMux I__5186 (
            .O(N__27900),
            .I(N__27897));
    LocalMux I__5185 (
            .O(N__27897),
            .I(N__27894));
    Odrv12 I__5184 (
            .O(N__27894),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_14 ));
    InMux I__5183 (
            .O(N__27891),
            .I(N__27886));
    CascadeMux I__5182 (
            .O(N__27890),
            .I(N__27883));
    InMux I__5181 (
            .O(N__27889),
            .I(N__27880));
    LocalMux I__5180 (
            .O(N__27886),
            .I(N__27877));
    InMux I__5179 (
            .O(N__27883),
            .I(N__27874));
    LocalMux I__5178 (
            .O(N__27880),
            .I(N__27870));
    Span4Mux_h I__5177 (
            .O(N__27877),
            .I(N__27867));
    LocalMux I__5176 (
            .O(N__27874),
            .I(N__27864));
    InMux I__5175 (
            .O(N__27873),
            .I(N__27861));
    Span4Mux_v I__5174 (
            .O(N__27870),
            .I(N__27858));
    Span4Mux_h I__5173 (
            .O(N__27867),
            .I(N__27855));
    Span4Mux_v I__5172 (
            .O(N__27864),
            .I(N__27852));
    LocalMux I__5171 (
            .O(N__27861),
            .I(\c0.FRAME_MATCHER_i_16 ));
    Odrv4 I__5170 (
            .O(N__27858),
            .I(\c0.FRAME_MATCHER_i_16 ));
    Odrv4 I__5169 (
            .O(N__27855),
            .I(\c0.FRAME_MATCHER_i_16 ));
    Odrv4 I__5168 (
            .O(N__27852),
            .I(\c0.FRAME_MATCHER_i_16 ));
    CascadeMux I__5167 (
            .O(N__27843),
            .I(N__27836));
    InMux I__5166 (
            .O(N__27842),
            .I(N__27823));
    InMux I__5165 (
            .O(N__27841),
            .I(N__27823));
    InMux I__5164 (
            .O(N__27840),
            .I(N__27823));
    InMux I__5163 (
            .O(N__27839),
            .I(N__27813));
    InMux I__5162 (
            .O(N__27836),
            .I(N__27808));
    InMux I__5161 (
            .O(N__27835),
            .I(N__27808));
    InMux I__5160 (
            .O(N__27834),
            .I(N__27805));
    CascadeMux I__5159 (
            .O(N__27833),
            .I(N__27802));
    CascadeMux I__5158 (
            .O(N__27832),
            .I(N__27790));
    CascadeMux I__5157 (
            .O(N__27831),
            .I(N__27787));
    CascadeMux I__5156 (
            .O(N__27830),
            .I(N__27783));
    LocalMux I__5155 (
            .O(N__27823),
            .I(N__27777));
    InMux I__5154 (
            .O(N__27822),
            .I(N__27770));
    InMux I__5153 (
            .O(N__27821),
            .I(N__27770));
    InMux I__5152 (
            .O(N__27820),
            .I(N__27770));
    InMux I__5151 (
            .O(N__27819),
            .I(N__27761));
    InMux I__5150 (
            .O(N__27818),
            .I(N__27761));
    InMux I__5149 (
            .O(N__27817),
            .I(N__27761));
    InMux I__5148 (
            .O(N__27816),
            .I(N__27761));
    LocalMux I__5147 (
            .O(N__27813),
            .I(N__27756));
    LocalMux I__5146 (
            .O(N__27808),
            .I(N__27756));
    LocalMux I__5145 (
            .O(N__27805),
            .I(N__27753));
    InMux I__5144 (
            .O(N__27802),
            .I(N__27748));
    InMux I__5143 (
            .O(N__27801),
            .I(N__27748));
    InMux I__5142 (
            .O(N__27800),
            .I(N__27739));
    InMux I__5141 (
            .O(N__27799),
            .I(N__27739));
    InMux I__5140 (
            .O(N__27798),
            .I(N__27739));
    InMux I__5139 (
            .O(N__27797),
            .I(N__27739));
    InMux I__5138 (
            .O(N__27796),
            .I(N__27730));
    InMux I__5137 (
            .O(N__27795),
            .I(N__27730));
    InMux I__5136 (
            .O(N__27794),
            .I(N__27730));
    InMux I__5135 (
            .O(N__27793),
            .I(N__27730));
    InMux I__5134 (
            .O(N__27790),
            .I(N__27721));
    InMux I__5133 (
            .O(N__27787),
            .I(N__27721));
    InMux I__5132 (
            .O(N__27786),
            .I(N__27721));
    InMux I__5131 (
            .O(N__27783),
            .I(N__27721));
    InMux I__5130 (
            .O(N__27782),
            .I(N__27714));
    InMux I__5129 (
            .O(N__27781),
            .I(N__27714));
    InMux I__5128 (
            .O(N__27780),
            .I(N__27714));
    Span12Mux_s3_h I__5127 (
            .O(N__27777),
            .I(N__27709));
    LocalMux I__5126 (
            .O(N__27770),
            .I(N__27709));
    LocalMux I__5125 (
            .O(N__27761),
            .I(N__27702));
    Span4Mux_h I__5124 (
            .O(N__27756),
            .I(N__27702));
    Span4Mux_v I__5123 (
            .O(N__27753),
            .I(N__27702));
    LocalMux I__5122 (
            .O(N__27748),
            .I(\c0.n10009 ));
    LocalMux I__5121 (
            .O(N__27739),
            .I(\c0.n10009 ));
    LocalMux I__5120 (
            .O(N__27730),
            .I(\c0.n10009 ));
    LocalMux I__5119 (
            .O(N__27721),
            .I(\c0.n10009 ));
    LocalMux I__5118 (
            .O(N__27714),
            .I(\c0.n10009 ));
    Odrv12 I__5117 (
            .O(N__27709),
            .I(\c0.n10009 ));
    Odrv4 I__5116 (
            .O(N__27702),
            .I(\c0.n10009 ));
    SRMux I__5115 (
            .O(N__27687),
            .I(N__27684));
    LocalMux I__5114 (
            .O(N__27684),
            .I(N__27681));
    Span4Mux_h I__5113 (
            .O(N__27681),
            .I(N__27678));
    Odrv4 I__5112 (
            .O(N__27678),
            .I(\c0.n3_adj_2259 ));
    InMux I__5111 (
            .O(N__27675),
            .I(N__27672));
    LocalMux I__5110 (
            .O(N__27672),
            .I(n26_adj_2423));
    InMux I__5109 (
            .O(N__27669),
            .I(bfn_9_29_0_));
    InMux I__5108 (
            .O(N__27666),
            .I(N__27663));
    LocalMux I__5107 (
            .O(N__27663),
            .I(n25_adj_2424));
    InMux I__5106 (
            .O(N__27660),
            .I(n16041));
    CascadeMux I__5105 (
            .O(N__27657),
            .I(N__27652));
    InMux I__5104 (
            .O(N__27656),
            .I(N__27649));
    InMux I__5103 (
            .O(N__27655),
            .I(N__27645));
    InMux I__5102 (
            .O(N__27652),
            .I(N__27642));
    LocalMux I__5101 (
            .O(N__27649),
            .I(N__27639));
    InMux I__5100 (
            .O(N__27648),
            .I(N__27636));
    LocalMux I__5099 (
            .O(N__27645),
            .I(N__27632));
    LocalMux I__5098 (
            .O(N__27642),
            .I(N__27627));
    Span4Mux_v I__5097 (
            .O(N__27639),
            .I(N__27627));
    LocalMux I__5096 (
            .O(N__27636),
            .I(N__27624));
    InMux I__5095 (
            .O(N__27635),
            .I(N__27621));
    Span4Mux_h I__5094 (
            .O(N__27632),
            .I(N__27616));
    Span4Mux_h I__5093 (
            .O(N__27627),
            .I(N__27616));
    Span12Mux_s5_h I__5092 (
            .O(N__27624),
            .I(N__27613));
    LocalMux I__5091 (
            .O(N__27621),
            .I(data_out_frame2_16_7));
    Odrv4 I__5090 (
            .O(N__27616),
            .I(data_out_frame2_16_7));
    Odrv12 I__5089 (
            .O(N__27613),
            .I(data_out_frame2_16_7));
    InMux I__5088 (
            .O(N__27606),
            .I(N__27603));
    LocalMux I__5087 (
            .O(N__27603),
            .I(N__27600));
    Span4Mux_v I__5086 (
            .O(N__27600),
            .I(N__27597));
    Span4Mux_h I__5085 (
            .O(N__27597),
            .I(N__27592));
    InMux I__5084 (
            .O(N__27596),
            .I(N__27589));
    InMux I__5083 (
            .O(N__27595),
            .I(N__27586));
    Odrv4 I__5082 (
            .O(N__27592),
            .I(\c0.n17194 ));
    LocalMux I__5081 (
            .O(N__27589),
            .I(\c0.n17194 ));
    LocalMux I__5080 (
            .O(N__27586),
            .I(\c0.n17194 ));
    InMux I__5079 (
            .O(N__27579),
            .I(N__27576));
    LocalMux I__5078 (
            .O(N__27576),
            .I(N__27573));
    Span4Mux_h I__5077 (
            .O(N__27573),
            .I(N__27570));
    Odrv4 I__5076 (
            .O(N__27570),
            .I(\c0.n10459 ));
    CascadeMux I__5075 (
            .O(N__27567),
            .I(N__27563));
    InMux I__5074 (
            .O(N__27566),
            .I(N__27557));
    InMux I__5073 (
            .O(N__27563),
            .I(N__27557));
    InMux I__5072 (
            .O(N__27562),
            .I(N__27554));
    LocalMux I__5071 (
            .O(N__27557),
            .I(N__27551));
    LocalMux I__5070 (
            .O(N__27554),
            .I(data_in_0_5));
    Odrv4 I__5069 (
            .O(N__27551),
            .I(data_in_0_5));
    InMux I__5068 (
            .O(N__27546),
            .I(N__27542));
    InMux I__5067 (
            .O(N__27545),
            .I(N__27539));
    LocalMux I__5066 (
            .O(N__27542),
            .I(N__27536));
    LocalMux I__5065 (
            .O(N__27539),
            .I(data_in_0_4));
    Odrv12 I__5064 (
            .O(N__27536),
            .I(data_in_0_4));
    InMux I__5063 (
            .O(N__27531),
            .I(N__27527));
    InMux I__5062 (
            .O(N__27530),
            .I(N__27524));
    LocalMux I__5061 (
            .O(N__27527),
            .I(N__27521));
    LocalMux I__5060 (
            .O(N__27524),
            .I(data_in_0_2));
    Odrv12 I__5059 (
            .O(N__27521),
            .I(data_in_0_2));
    InMux I__5058 (
            .O(N__27516),
            .I(N__27511));
    InMux I__5057 (
            .O(N__27515),
            .I(N__27506));
    InMux I__5056 (
            .O(N__27514),
            .I(N__27506));
    LocalMux I__5055 (
            .O(N__27511),
            .I(N__27503));
    LocalMux I__5054 (
            .O(N__27506),
            .I(data_in_1_5));
    Odrv12 I__5053 (
            .O(N__27503),
            .I(data_in_1_5));
    InMux I__5052 (
            .O(N__27498),
            .I(N__27495));
    LocalMux I__5051 (
            .O(N__27495),
            .I(N__27492));
    Span4Mux_h I__5050 (
            .O(N__27492),
            .I(N__27489));
    Span4Mux_h I__5049 (
            .O(N__27489),
            .I(N__27486));
    Odrv4 I__5048 (
            .O(N__27486),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_16 ));
    InMux I__5047 (
            .O(N__27483),
            .I(N__27478));
    InMux I__5046 (
            .O(N__27482),
            .I(N__27475));
    InMux I__5045 (
            .O(N__27481),
            .I(N__27472));
    LocalMux I__5044 (
            .O(N__27478),
            .I(N__27467));
    LocalMux I__5043 (
            .O(N__27475),
            .I(N__27467));
    LocalMux I__5042 (
            .O(N__27472),
            .I(\c0.FRAME_MATCHER_state_4 ));
    Odrv4 I__5041 (
            .O(N__27467),
            .I(\c0.FRAME_MATCHER_state_4 ));
    SRMux I__5040 (
            .O(N__27462),
            .I(N__27459));
    LocalMux I__5039 (
            .O(N__27459),
            .I(N__27456));
    Odrv12 I__5038 (
            .O(N__27456),
            .I(\c0.n16716 ));
    InMux I__5037 (
            .O(N__27453),
            .I(N__27444));
    InMux I__5036 (
            .O(N__27452),
            .I(N__27444));
    InMux I__5035 (
            .O(N__27451),
            .I(N__27444));
    LocalMux I__5034 (
            .O(N__27444),
            .I(\c0.FRAME_MATCHER_state_13 ));
    SRMux I__5033 (
            .O(N__27441),
            .I(N__27438));
    LocalMux I__5032 (
            .O(N__27438),
            .I(N__27435));
    Odrv4 I__5031 (
            .O(N__27435),
            .I(\c0.n8_adj_2332 ));
    InMux I__5030 (
            .O(N__27432),
            .I(N__27425));
    InMux I__5029 (
            .O(N__27431),
            .I(N__27425));
    CascadeMux I__5028 (
            .O(N__27430),
            .I(N__27422));
    LocalMux I__5027 (
            .O(N__27425),
            .I(N__27419));
    InMux I__5026 (
            .O(N__27422),
            .I(N__27416));
    Span4Mux_h I__5025 (
            .O(N__27419),
            .I(N__27413));
    LocalMux I__5024 (
            .O(N__27416),
            .I(\c0.FRAME_MATCHER_state_19 ));
    Odrv4 I__5023 (
            .O(N__27413),
            .I(\c0.FRAME_MATCHER_state_19 ));
    SRMux I__5022 (
            .O(N__27408),
            .I(N__27405));
    LocalMux I__5021 (
            .O(N__27405),
            .I(N__27402));
    Span4Mux_h I__5020 (
            .O(N__27402),
            .I(N__27399));
    Odrv4 I__5019 (
            .O(N__27399),
            .I(\c0.n8_adj_2328 ));
    InMux I__5018 (
            .O(N__27396),
            .I(N__27392));
    CascadeMux I__5017 (
            .O(N__27395),
            .I(N__27388));
    LocalMux I__5016 (
            .O(N__27392),
            .I(N__27385));
    InMux I__5015 (
            .O(N__27391),
            .I(N__27382));
    InMux I__5014 (
            .O(N__27388),
            .I(N__27379));
    Span4Mux_h I__5013 (
            .O(N__27385),
            .I(N__27374));
    LocalMux I__5012 (
            .O(N__27382),
            .I(N__27374));
    LocalMux I__5011 (
            .O(N__27379),
            .I(N__27371));
    Span4Mux_h I__5010 (
            .O(N__27374),
            .I(N__27368));
    Odrv4 I__5009 (
            .O(N__27371),
            .I(\c0.FRAME_MATCHER_state_6 ));
    Odrv4 I__5008 (
            .O(N__27368),
            .I(\c0.FRAME_MATCHER_state_6 ));
    SRMux I__5007 (
            .O(N__27363),
            .I(N__27360));
    LocalMux I__5006 (
            .O(N__27360),
            .I(N__27357));
    Span4Mux_v I__5005 (
            .O(N__27357),
            .I(N__27354));
    Odrv4 I__5004 (
            .O(N__27354),
            .I(\c0.n8_adj_2334 ));
    InMux I__5003 (
            .O(N__27351),
            .I(N__27348));
    LocalMux I__5002 (
            .O(N__27348),
            .I(N__27343));
    InMux I__5001 (
            .O(N__27347),
            .I(N__27338));
    InMux I__5000 (
            .O(N__27346),
            .I(N__27338));
    Odrv4 I__4999 (
            .O(N__27343),
            .I(\c0.FRAME_MATCHER_state_12 ));
    LocalMux I__4998 (
            .O(N__27338),
            .I(\c0.FRAME_MATCHER_state_12 ));
    SRMux I__4997 (
            .O(N__27333),
            .I(N__27330));
    LocalMux I__4996 (
            .O(N__27330),
            .I(N__27327));
    Odrv4 I__4995 (
            .O(N__27327),
            .I(\c0.n16708 ));
    InMux I__4994 (
            .O(N__27324),
            .I(N__27319));
    InMux I__4993 (
            .O(N__27323),
            .I(N__27316));
    CascadeMux I__4992 (
            .O(N__27322),
            .I(N__27313));
    LocalMux I__4991 (
            .O(N__27319),
            .I(N__27308));
    LocalMux I__4990 (
            .O(N__27316),
            .I(N__27308));
    InMux I__4989 (
            .O(N__27313),
            .I(N__27305));
    Span4Mux_h I__4988 (
            .O(N__27308),
            .I(N__27302));
    LocalMux I__4987 (
            .O(N__27305),
            .I(\c0.FRAME_MATCHER_state_14 ));
    Odrv4 I__4986 (
            .O(N__27302),
            .I(\c0.FRAME_MATCHER_state_14 ));
    SRMux I__4985 (
            .O(N__27297),
            .I(N__27294));
    LocalMux I__4984 (
            .O(N__27294),
            .I(N__27291));
    Span4Mux_h I__4983 (
            .O(N__27291),
            .I(N__27288));
    Span4Mux_v I__4982 (
            .O(N__27288),
            .I(N__27285));
    Odrv4 I__4981 (
            .O(N__27285),
            .I(\c0.n8_adj_2331 ));
    CascadeMux I__4980 (
            .O(N__27282),
            .I(N__27278));
    InMux I__4979 (
            .O(N__27281),
            .I(N__27272));
    InMux I__4978 (
            .O(N__27278),
            .I(N__27272));
    InMux I__4977 (
            .O(N__27277),
            .I(N__27269));
    LocalMux I__4976 (
            .O(N__27272),
            .I(data_in_0_6));
    LocalMux I__4975 (
            .O(N__27269),
            .I(data_in_0_6));
    InMux I__4974 (
            .O(N__27264),
            .I(N__27260));
    InMux I__4973 (
            .O(N__27263),
            .I(N__27255));
    LocalMux I__4972 (
            .O(N__27260),
            .I(N__27252));
    InMux I__4971 (
            .O(N__27259),
            .I(N__27249));
    InMux I__4970 (
            .O(N__27258),
            .I(N__27246));
    LocalMux I__4969 (
            .O(N__27255),
            .I(N__27243));
    Span4Mux_v I__4968 (
            .O(N__27252),
            .I(N__27240));
    LocalMux I__4967 (
            .O(N__27249),
            .I(N__27235));
    LocalMux I__4966 (
            .O(N__27246),
            .I(N__27235));
    Span4Mux_v I__4965 (
            .O(N__27243),
            .I(N__27232));
    Span4Mux_h I__4964 (
            .O(N__27240),
            .I(N__27227));
    Span4Mux_v I__4963 (
            .O(N__27235),
            .I(N__27227));
    Odrv4 I__4962 (
            .O(N__27232),
            .I(\c0.FRAME_MATCHER_i_15 ));
    Odrv4 I__4961 (
            .O(N__27227),
            .I(\c0.FRAME_MATCHER_i_15 ));
    InMux I__4960 (
            .O(N__27222),
            .I(N__27219));
    LocalMux I__4959 (
            .O(N__27219),
            .I(N__27216));
    Span12Mux_s8_v I__4958 (
            .O(N__27216),
            .I(N__27213));
    Odrv12 I__4957 (
            .O(N__27213),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_15 ));
    InMux I__4956 (
            .O(N__27210),
            .I(N__27207));
    LocalMux I__4955 (
            .O(N__27207),
            .I(N__27203));
    CascadeMux I__4954 (
            .O(N__27206),
            .I(N__27199));
    Span4Mux_h I__4953 (
            .O(N__27203),
            .I(N__27195));
    InMux I__4952 (
            .O(N__27202),
            .I(N__27192));
    InMux I__4951 (
            .O(N__27199),
            .I(N__27189));
    InMux I__4950 (
            .O(N__27198),
            .I(N__27186));
    Span4Mux_v I__4949 (
            .O(N__27195),
            .I(N__27179));
    LocalMux I__4948 (
            .O(N__27192),
            .I(N__27179));
    LocalMux I__4947 (
            .O(N__27189),
            .I(N__27179));
    LocalMux I__4946 (
            .O(N__27186),
            .I(\c0.FRAME_MATCHER_i_13 ));
    Odrv4 I__4945 (
            .O(N__27179),
            .I(\c0.FRAME_MATCHER_i_13 ));
    InMux I__4944 (
            .O(N__27174),
            .I(N__27171));
    LocalMux I__4943 (
            .O(N__27171),
            .I(N__27168));
    Span4Mux_v I__4942 (
            .O(N__27168),
            .I(N__27165));
    Span4Mux_h I__4941 (
            .O(N__27165),
            .I(N__27162));
    Odrv4 I__4940 (
            .O(N__27162),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_13 ));
    InMux I__4939 (
            .O(N__27159),
            .I(N__27155));
    InMux I__4938 (
            .O(N__27158),
            .I(N__27152));
    LocalMux I__4937 (
            .O(N__27155),
            .I(N__27148));
    LocalMux I__4936 (
            .O(N__27152),
            .I(N__27144));
    InMux I__4935 (
            .O(N__27151),
            .I(N__27141));
    Span4Mux_v I__4934 (
            .O(N__27148),
            .I(N__27138));
    InMux I__4933 (
            .O(N__27147),
            .I(N__27135));
    Span4Mux_h I__4932 (
            .O(N__27144),
            .I(N__27132));
    LocalMux I__4931 (
            .O(N__27141),
            .I(N__27125));
    Span4Mux_h I__4930 (
            .O(N__27138),
            .I(N__27125));
    LocalMux I__4929 (
            .O(N__27135),
            .I(N__27125));
    Span4Mux_s0_h I__4928 (
            .O(N__27132),
            .I(N__27122));
    Span4Mux_h I__4927 (
            .O(N__27125),
            .I(N__27119));
    Odrv4 I__4926 (
            .O(N__27122),
            .I(\c0.FRAME_MATCHER_i_11 ));
    Odrv4 I__4925 (
            .O(N__27119),
            .I(\c0.FRAME_MATCHER_i_11 ));
    InMux I__4924 (
            .O(N__27114),
            .I(N__27111));
    LocalMux I__4923 (
            .O(N__27111),
            .I(N__27108));
    Span4Mux_h I__4922 (
            .O(N__27108),
            .I(N__27105));
    Span4Mux_v I__4921 (
            .O(N__27105),
            .I(N__27102));
    Odrv4 I__4920 (
            .O(N__27102),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_11 ));
    InMux I__4919 (
            .O(N__27099),
            .I(N__27096));
    LocalMux I__4918 (
            .O(N__27096),
            .I(N__27092));
    CascadeMux I__4917 (
            .O(N__27095),
            .I(N__27089));
    Span4Mux_h I__4916 (
            .O(N__27092),
            .I(N__27086));
    InMux I__4915 (
            .O(N__27089),
            .I(N__27083));
    Span4Mux_h I__4914 (
            .O(N__27086),
            .I(N__27078));
    LocalMux I__4913 (
            .O(N__27083),
            .I(N__27075));
    InMux I__4912 (
            .O(N__27082),
            .I(N__27070));
    InMux I__4911 (
            .O(N__27081),
            .I(N__27070));
    Odrv4 I__4910 (
            .O(N__27078),
            .I(\c0.FRAME_MATCHER_i_7 ));
    Odrv4 I__4909 (
            .O(N__27075),
            .I(\c0.FRAME_MATCHER_i_7 ));
    LocalMux I__4908 (
            .O(N__27070),
            .I(\c0.FRAME_MATCHER_i_7 ));
    InMux I__4907 (
            .O(N__27063),
            .I(N__27060));
    LocalMux I__4906 (
            .O(N__27060),
            .I(N__27057));
    Span4Mux_h I__4905 (
            .O(N__27057),
            .I(N__27054));
    Span4Mux_h I__4904 (
            .O(N__27054),
            .I(N__27051));
    Odrv4 I__4903 (
            .O(N__27051),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_7 ));
    InMux I__4902 (
            .O(N__27048),
            .I(N__27045));
    LocalMux I__4901 (
            .O(N__27045),
            .I(N__27042));
    Span4Mux_h I__4900 (
            .O(N__27042),
            .I(N__27039));
    Span4Mux_h I__4899 (
            .O(N__27039),
            .I(N__27036));
    Odrv4 I__4898 (
            .O(N__27036),
            .I(\c0.n37 ));
    InMux I__4897 (
            .O(N__27033),
            .I(N__27030));
    LocalMux I__4896 (
            .O(N__27030),
            .I(N__27027));
    Span4Mux_h I__4895 (
            .O(N__27027),
            .I(N__27021));
    InMux I__4894 (
            .O(N__27026),
            .I(N__27016));
    InMux I__4893 (
            .O(N__27025),
            .I(N__27016));
    InMux I__4892 (
            .O(N__27024),
            .I(N__27013));
    Span4Mux_v I__4891 (
            .O(N__27021),
            .I(N__27008));
    LocalMux I__4890 (
            .O(N__27016),
            .I(N__27008));
    LocalMux I__4889 (
            .O(N__27013),
            .I(N__27005));
    Span4Mux_h I__4888 (
            .O(N__27008),
            .I(N__27002));
    Odrv4 I__4887 (
            .O(N__27005),
            .I(\c0.FRAME_MATCHER_i_28 ));
    Odrv4 I__4886 (
            .O(N__27002),
            .I(\c0.FRAME_MATCHER_i_28 ));
    InMux I__4885 (
            .O(N__26997),
            .I(N__26994));
    LocalMux I__4884 (
            .O(N__26994),
            .I(N__26991));
    Sp12to4 I__4883 (
            .O(N__26991),
            .I(N__26988));
    Span12Mux_s8_h I__4882 (
            .O(N__26988),
            .I(N__26985));
    Odrv12 I__4881 (
            .O(N__26985),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_28 ));
    CascadeMux I__4880 (
            .O(N__26982),
            .I(\c0.n17331_cascade_ ));
    InMux I__4879 (
            .O(N__26979),
            .I(N__26976));
    LocalMux I__4878 (
            .O(N__26976),
            .I(\c0.n17410 ));
    InMux I__4877 (
            .O(N__26973),
            .I(N__26970));
    LocalMux I__4876 (
            .O(N__26970),
            .I(N__26967));
    Span4Mux_s1_v I__4875 (
            .O(N__26967),
            .I(N__26964));
    Span4Mux_v I__4874 (
            .O(N__26964),
            .I(N__26959));
    InMux I__4873 (
            .O(N__26963),
            .I(N__26956));
    InMux I__4872 (
            .O(N__26962),
            .I(N__26953));
    Span4Mux_v I__4871 (
            .O(N__26959),
            .I(N__26948));
    LocalMux I__4870 (
            .O(N__26956),
            .I(N__26948));
    LocalMux I__4869 (
            .O(N__26953),
            .I(data_in_2_6));
    Odrv4 I__4868 (
            .O(N__26948),
            .I(data_in_2_6));
    InMux I__4867 (
            .O(N__26943),
            .I(N__26940));
    LocalMux I__4866 (
            .O(N__26940),
            .I(\c0.n12_adj_2355 ));
    InMux I__4865 (
            .O(N__26937),
            .I(N__26932));
    InMux I__4864 (
            .O(N__26936),
            .I(N__26927));
    InMux I__4863 (
            .O(N__26935),
            .I(N__26927));
    LocalMux I__4862 (
            .O(N__26932),
            .I(data_in_2_4));
    LocalMux I__4861 (
            .O(N__26927),
            .I(data_in_2_4));
    SRMux I__4860 (
            .O(N__26922),
            .I(N__26919));
    LocalMux I__4859 (
            .O(N__26919),
            .I(N__26916));
    Odrv12 I__4858 (
            .O(N__26916),
            .I(\c0.n4_adj_2150 ));
    InMux I__4857 (
            .O(N__26913),
            .I(N__26910));
    LocalMux I__4856 (
            .O(N__26910),
            .I(\c0.n10133 ));
    InMux I__4855 (
            .O(N__26907),
            .I(N__26904));
    LocalMux I__4854 (
            .O(N__26904),
            .I(\c0.n17406 ));
    InMux I__4853 (
            .O(N__26901),
            .I(N__26892));
    InMux I__4852 (
            .O(N__26900),
            .I(N__26892));
    InMux I__4851 (
            .O(N__26899),
            .I(N__26892));
    LocalMux I__4850 (
            .O(N__26892),
            .I(data_in_0_3));
    CascadeMux I__4849 (
            .O(N__26889),
            .I(\c0.n10133_cascade_ ));
    CascadeMux I__4848 (
            .O(N__26886),
            .I(\c0.n6_adj_2356_cascade_ ));
    CascadeMux I__4847 (
            .O(N__26883),
            .I(\c0.n10027_cascade_ ));
    InMux I__4846 (
            .O(N__26880),
            .I(N__26876));
    InMux I__4845 (
            .O(N__26879),
            .I(N__26873));
    LocalMux I__4844 (
            .O(N__26876),
            .I(data_in_0_7));
    LocalMux I__4843 (
            .O(N__26873),
            .I(data_in_0_7));
    InMux I__4842 (
            .O(N__26868),
            .I(N__26861));
    InMux I__4841 (
            .O(N__26867),
            .I(N__26861));
    InMux I__4840 (
            .O(N__26866),
            .I(N__26858));
    LocalMux I__4839 (
            .O(N__26861),
            .I(data_in_1_3));
    LocalMux I__4838 (
            .O(N__26858),
            .I(data_in_1_3));
    InMux I__4837 (
            .O(N__26853),
            .I(N__26849));
    InMux I__4836 (
            .O(N__26852),
            .I(N__26844));
    LocalMux I__4835 (
            .O(N__26849),
            .I(N__26841));
    CascadeMux I__4834 (
            .O(N__26848),
            .I(N__26836));
    InMux I__4833 (
            .O(N__26847),
            .I(N__26833));
    LocalMux I__4832 (
            .O(N__26844),
            .I(N__26830));
    Span4Mux_h I__4831 (
            .O(N__26841),
            .I(N__26827));
    InMux I__4830 (
            .O(N__26840),
            .I(N__26823));
    InMux I__4829 (
            .O(N__26839),
            .I(N__26820));
    InMux I__4828 (
            .O(N__26836),
            .I(N__26815));
    LocalMux I__4827 (
            .O(N__26833),
            .I(N__26810));
    Span4Mux_h I__4826 (
            .O(N__26830),
            .I(N__26810));
    Span4Mux_v I__4825 (
            .O(N__26827),
            .I(N__26807));
    InMux I__4824 (
            .O(N__26826),
            .I(N__26804));
    LocalMux I__4823 (
            .O(N__26823),
            .I(N__26799));
    LocalMux I__4822 (
            .O(N__26820),
            .I(N__26799));
    InMux I__4821 (
            .O(N__26819),
            .I(N__26794));
    InMux I__4820 (
            .O(N__26818),
            .I(N__26794));
    LocalMux I__4819 (
            .O(N__26815),
            .I(N__26791));
    Span4Mux_v I__4818 (
            .O(N__26810),
            .I(N__26788));
    Span4Mux_v I__4817 (
            .O(N__26807),
            .I(N__26785));
    LocalMux I__4816 (
            .O(N__26804),
            .I(N__26780));
    Span4Mux_h I__4815 (
            .O(N__26799),
            .I(N__26780));
    LocalMux I__4814 (
            .O(N__26794),
            .I(r_SM_Main_2_adj_2438));
    Odrv12 I__4813 (
            .O(N__26791),
            .I(r_SM_Main_2_adj_2438));
    Odrv4 I__4812 (
            .O(N__26788),
            .I(r_SM_Main_2_adj_2438));
    Odrv4 I__4811 (
            .O(N__26785),
            .I(r_SM_Main_2_adj_2438));
    Odrv4 I__4810 (
            .O(N__26780),
            .I(r_SM_Main_2_adj_2438));
    InMux I__4809 (
            .O(N__26769),
            .I(N__26766));
    LocalMux I__4808 (
            .O(N__26766),
            .I(N__26763));
    Span4Mux_v I__4807 (
            .O(N__26763),
            .I(N__26760));
    Span4Mux_h I__4806 (
            .O(N__26760),
            .I(N__26757));
    Odrv4 I__4805 (
            .O(N__26757),
            .I(n4_adj_2484));
    CascadeMux I__4804 (
            .O(N__26754),
            .I(N__26747));
    CascadeMux I__4803 (
            .O(N__26753),
            .I(N__26743));
    InMux I__4802 (
            .O(N__26752),
            .I(N__26735));
    InMux I__4801 (
            .O(N__26751),
            .I(N__26735));
    InMux I__4800 (
            .O(N__26750),
            .I(N__26730));
    InMux I__4799 (
            .O(N__26747),
            .I(N__26730));
    InMux I__4798 (
            .O(N__26746),
            .I(N__26727));
    InMux I__4797 (
            .O(N__26743),
            .I(N__26724));
    InMux I__4796 (
            .O(N__26742),
            .I(N__26721));
    CascadeMux I__4795 (
            .O(N__26741),
            .I(N__26717));
    CascadeMux I__4794 (
            .O(N__26740),
            .I(N__26714));
    LocalMux I__4793 (
            .O(N__26735),
            .I(N__26711));
    LocalMux I__4792 (
            .O(N__26730),
            .I(N__26708));
    LocalMux I__4791 (
            .O(N__26727),
            .I(N__26705));
    LocalMux I__4790 (
            .O(N__26724),
            .I(N__26702));
    LocalMux I__4789 (
            .O(N__26721),
            .I(N__26699));
    InMux I__4788 (
            .O(N__26720),
            .I(N__26696));
    InMux I__4787 (
            .O(N__26717),
            .I(N__26691));
    InMux I__4786 (
            .O(N__26714),
            .I(N__26691));
    Span4Mux_h I__4785 (
            .O(N__26711),
            .I(N__26686));
    Span4Mux_h I__4784 (
            .O(N__26708),
            .I(N__26686));
    Span4Mux_h I__4783 (
            .O(N__26705),
            .I(N__26679));
    Span4Mux_h I__4782 (
            .O(N__26702),
            .I(N__26679));
    Span4Mux_h I__4781 (
            .O(N__26699),
            .I(N__26679));
    LocalMux I__4780 (
            .O(N__26696),
            .I(r_SM_Main_1_adj_2439));
    LocalMux I__4779 (
            .O(N__26691),
            .I(r_SM_Main_1_adj_2439));
    Odrv4 I__4778 (
            .O(N__26686),
            .I(r_SM_Main_1_adj_2439));
    Odrv4 I__4777 (
            .O(N__26679),
            .I(r_SM_Main_1_adj_2439));
    InMux I__4776 (
            .O(N__26670),
            .I(\c0.n15977 ));
    InMux I__4775 (
            .O(N__26667),
            .I(\c0.n15978 ));
    InMux I__4774 (
            .O(N__26664),
            .I(N__26661));
    LocalMux I__4773 (
            .O(N__26661),
            .I(N__26658));
    Span4Mux_h I__4772 (
            .O(N__26658),
            .I(N__26655));
    Odrv4 I__4771 (
            .O(N__26655),
            .I(\c0.n17714 ));
    InMux I__4770 (
            .O(N__26652),
            .I(N__26649));
    LocalMux I__4769 (
            .O(N__26649),
            .I(\c0.n17589 ));
    InMux I__4768 (
            .O(N__26646),
            .I(N__26640));
    InMux I__4767 (
            .O(N__26645),
            .I(N__26640));
    LocalMux I__4766 (
            .O(N__26640),
            .I(N__26636));
    CascadeMux I__4765 (
            .O(N__26639),
            .I(N__26633));
    Span4Mux_v I__4764 (
            .O(N__26636),
            .I(N__26629));
    InMux I__4763 (
            .O(N__26633),
            .I(N__26626));
    InMux I__4762 (
            .O(N__26632),
            .I(N__26623));
    Sp12to4 I__4761 (
            .O(N__26629),
            .I(N__26618));
    LocalMux I__4760 (
            .O(N__26626),
            .I(N__26618));
    LocalMux I__4759 (
            .O(N__26623),
            .I(data_out_frame2_7_1));
    Odrv12 I__4758 (
            .O(N__26618),
            .I(data_out_frame2_7_1));
    InMux I__4757 (
            .O(N__26613),
            .I(N__26602));
    InMux I__4756 (
            .O(N__26612),
            .I(N__26602));
    CEMux I__4755 (
            .O(N__26611),
            .I(N__26593));
    CEMux I__4754 (
            .O(N__26610),
            .I(N__26590));
    CEMux I__4753 (
            .O(N__26609),
            .I(N__26568));
    CEMux I__4752 (
            .O(N__26608),
            .I(N__26551));
    CEMux I__4751 (
            .O(N__26607),
            .I(N__26548));
    LocalMux I__4750 (
            .O(N__26602),
            .I(N__26539));
    InMux I__4749 (
            .O(N__26601),
            .I(N__26531));
    InMux I__4748 (
            .O(N__26600),
            .I(N__26531));
    InMux I__4747 (
            .O(N__26599),
            .I(N__26531));
    InMux I__4746 (
            .O(N__26598),
            .I(N__26524));
    InMux I__4745 (
            .O(N__26597),
            .I(N__26524));
    InMux I__4744 (
            .O(N__26596),
            .I(N__26524));
    LocalMux I__4743 (
            .O(N__26593),
            .I(N__26519));
    LocalMux I__4742 (
            .O(N__26590),
            .I(N__26519));
    InMux I__4741 (
            .O(N__26589),
            .I(N__26501));
    InMux I__4740 (
            .O(N__26588),
            .I(N__26501));
    InMux I__4739 (
            .O(N__26587),
            .I(N__26501));
    InMux I__4738 (
            .O(N__26586),
            .I(N__26494));
    InMux I__4737 (
            .O(N__26585),
            .I(N__26494));
    InMux I__4736 (
            .O(N__26584),
            .I(N__26494));
    InMux I__4735 (
            .O(N__26583),
            .I(N__26491));
    InMux I__4734 (
            .O(N__26582),
            .I(N__26484));
    InMux I__4733 (
            .O(N__26581),
            .I(N__26484));
    InMux I__4732 (
            .O(N__26580),
            .I(N__26484));
    InMux I__4731 (
            .O(N__26579),
            .I(N__26475));
    InMux I__4730 (
            .O(N__26578),
            .I(N__26475));
    InMux I__4729 (
            .O(N__26577),
            .I(N__26475));
    InMux I__4728 (
            .O(N__26576),
            .I(N__26475));
    InMux I__4727 (
            .O(N__26575),
            .I(N__26464));
    InMux I__4726 (
            .O(N__26574),
            .I(N__26464));
    InMux I__4725 (
            .O(N__26573),
            .I(N__26464));
    InMux I__4724 (
            .O(N__26572),
            .I(N__26464));
    InMux I__4723 (
            .O(N__26571),
            .I(N__26464));
    LocalMux I__4722 (
            .O(N__26568),
            .I(N__26461));
    InMux I__4721 (
            .O(N__26567),
            .I(N__26452));
    InMux I__4720 (
            .O(N__26566),
            .I(N__26452));
    InMux I__4719 (
            .O(N__26565),
            .I(N__26452));
    CEMux I__4718 (
            .O(N__26564),
            .I(N__26449));
    InMux I__4717 (
            .O(N__26563),
            .I(N__26446));
    InMux I__4716 (
            .O(N__26562),
            .I(N__26443));
    InMux I__4715 (
            .O(N__26561),
            .I(N__26440));
    InMux I__4714 (
            .O(N__26560),
            .I(N__26433));
    InMux I__4713 (
            .O(N__26559),
            .I(N__26433));
    InMux I__4712 (
            .O(N__26558),
            .I(N__26433));
    InMux I__4711 (
            .O(N__26557),
            .I(N__26424));
    InMux I__4710 (
            .O(N__26556),
            .I(N__26424));
    InMux I__4709 (
            .O(N__26555),
            .I(N__26424));
    InMux I__4708 (
            .O(N__26554),
            .I(N__26424));
    LocalMux I__4707 (
            .O(N__26551),
            .I(N__26419));
    LocalMux I__4706 (
            .O(N__26548),
            .I(N__26419));
    CascadeMux I__4705 (
            .O(N__26547),
            .I(N__26416));
    InMux I__4704 (
            .O(N__26546),
            .I(N__26410));
    InMux I__4703 (
            .O(N__26545),
            .I(N__26410));
    CEMux I__4702 (
            .O(N__26544),
            .I(N__26407));
    CEMux I__4701 (
            .O(N__26543),
            .I(N__26404));
    CEMux I__4700 (
            .O(N__26542),
            .I(N__26401));
    Span4Mux_v I__4699 (
            .O(N__26539),
            .I(N__26398));
    InMux I__4698 (
            .O(N__26538),
            .I(N__26395));
    LocalMux I__4697 (
            .O(N__26531),
            .I(N__26390));
    LocalMux I__4696 (
            .O(N__26524),
            .I(N__26390));
    Span4Mux_v I__4695 (
            .O(N__26519),
            .I(N__26387));
    CEMux I__4694 (
            .O(N__26518),
            .I(N__26330));
    InMux I__4693 (
            .O(N__26517),
            .I(N__26327));
    InMux I__4692 (
            .O(N__26516),
            .I(N__26318));
    InMux I__4691 (
            .O(N__26515),
            .I(N__26318));
    InMux I__4690 (
            .O(N__26514),
            .I(N__26318));
    InMux I__4689 (
            .O(N__26513),
            .I(N__26318));
    InMux I__4688 (
            .O(N__26512),
            .I(N__26307));
    InMux I__4687 (
            .O(N__26511),
            .I(N__26307));
    InMux I__4686 (
            .O(N__26510),
            .I(N__26307));
    InMux I__4685 (
            .O(N__26509),
            .I(N__26307));
    InMux I__4684 (
            .O(N__26508),
            .I(N__26307));
    LocalMux I__4683 (
            .O(N__26501),
            .I(N__26304));
    LocalMux I__4682 (
            .O(N__26494),
            .I(N__26301));
    LocalMux I__4681 (
            .O(N__26491),
            .I(N__26290));
    LocalMux I__4680 (
            .O(N__26484),
            .I(N__26290));
    LocalMux I__4679 (
            .O(N__26475),
            .I(N__26290));
    LocalMux I__4678 (
            .O(N__26464),
            .I(N__26290));
    Span4Mux_v I__4677 (
            .O(N__26461),
            .I(N__26290));
    InMux I__4676 (
            .O(N__26460),
            .I(N__26285));
    InMux I__4675 (
            .O(N__26459),
            .I(N__26285));
    LocalMux I__4674 (
            .O(N__26452),
            .I(N__26282));
    LocalMux I__4673 (
            .O(N__26449),
            .I(N__26279));
    LocalMux I__4672 (
            .O(N__26446),
            .I(N__26270));
    LocalMux I__4671 (
            .O(N__26443),
            .I(N__26270));
    LocalMux I__4670 (
            .O(N__26440),
            .I(N__26270));
    LocalMux I__4669 (
            .O(N__26433),
            .I(N__26270));
    LocalMux I__4668 (
            .O(N__26424),
            .I(N__26265));
    Span4Mux_v I__4667 (
            .O(N__26419),
            .I(N__26265));
    InMux I__4666 (
            .O(N__26416),
            .I(N__26260));
    InMux I__4665 (
            .O(N__26415),
            .I(N__26260));
    LocalMux I__4664 (
            .O(N__26410),
            .I(N__26255));
    LocalMux I__4663 (
            .O(N__26407),
            .I(N__26255));
    LocalMux I__4662 (
            .O(N__26404),
            .I(N__26250));
    LocalMux I__4661 (
            .O(N__26401),
            .I(N__26250));
    Span4Mux_h I__4660 (
            .O(N__26398),
            .I(N__26241));
    LocalMux I__4659 (
            .O(N__26395),
            .I(N__26241));
    Span4Mux_v I__4658 (
            .O(N__26390),
            .I(N__26241));
    Span4Mux_s0_h I__4657 (
            .O(N__26387),
            .I(N__26241));
    InMux I__4656 (
            .O(N__26386),
            .I(N__26236));
    InMux I__4655 (
            .O(N__26385),
            .I(N__26236));
    InMux I__4654 (
            .O(N__26384),
            .I(N__26219));
    InMux I__4653 (
            .O(N__26383),
            .I(N__26219));
    InMux I__4652 (
            .O(N__26382),
            .I(N__26219));
    InMux I__4651 (
            .O(N__26381),
            .I(N__26219));
    InMux I__4650 (
            .O(N__26380),
            .I(N__26219));
    InMux I__4649 (
            .O(N__26379),
            .I(N__26219));
    InMux I__4648 (
            .O(N__26378),
            .I(N__26219));
    InMux I__4647 (
            .O(N__26377),
            .I(N__26219));
    InMux I__4646 (
            .O(N__26376),
            .I(N__26208));
    InMux I__4645 (
            .O(N__26375),
            .I(N__26208));
    InMux I__4644 (
            .O(N__26374),
            .I(N__26208));
    InMux I__4643 (
            .O(N__26373),
            .I(N__26208));
    InMux I__4642 (
            .O(N__26372),
            .I(N__26208));
    InMux I__4641 (
            .O(N__26371),
            .I(N__26193));
    InMux I__4640 (
            .O(N__26370),
            .I(N__26193));
    InMux I__4639 (
            .O(N__26369),
            .I(N__26193));
    InMux I__4638 (
            .O(N__26368),
            .I(N__26193));
    InMux I__4637 (
            .O(N__26367),
            .I(N__26193));
    InMux I__4636 (
            .O(N__26366),
            .I(N__26193));
    InMux I__4635 (
            .O(N__26365),
            .I(N__26193));
    InMux I__4634 (
            .O(N__26364),
            .I(N__26180));
    InMux I__4633 (
            .O(N__26363),
            .I(N__26180));
    InMux I__4632 (
            .O(N__26362),
            .I(N__26180));
    InMux I__4631 (
            .O(N__26361),
            .I(N__26180));
    InMux I__4630 (
            .O(N__26360),
            .I(N__26180));
    InMux I__4629 (
            .O(N__26359),
            .I(N__26180));
    InMux I__4628 (
            .O(N__26358),
            .I(N__26167));
    InMux I__4627 (
            .O(N__26357),
            .I(N__26167));
    InMux I__4626 (
            .O(N__26356),
            .I(N__26167));
    InMux I__4625 (
            .O(N__26355),
            .I(N__26167));
    InMux I__4624 (
            .O(N__26354),
            .I(N__26167));
    InMux I__4623 (
            .O(N__26353),
            .I(N__26167));
    InMux I__4622 (
            .O(N__26352),
            .I(N__26152));
    InMux I__4621 (
            .O(N__26351),
            .I(N__26152));
    InMux I__4620 (
            .O(N__26350),
            .I(N__26152));
    InMux I__4619 (
            .O(N__26349),
            .I(N__26152));
    InMux I__4618 (
            .O(N__26348),
            .I(N__26152));
    InMux I__4617 (
            .O(N__26347),
            .I(N__26152));
    InMux I__4616 (
            .O(N__26346),
            .I(N__26152));
    InMux I__4615 (
            .O(N__26345),
            .I(N__26135));
    InMux I__4614 (
            .O(N__26344),
            .I(N__26135));
    InMux I__4613 (
            .O(N__26343),
            .I(N__26135));
    InMux I__4612 (
            .O(N__26342),
            .I(N__26135));
    InMux I__4611 (
            .O(N__26341),
            .I(N__26135));
    InMux I__4610 (
            .O(N__26340),
            .I(N__26135));
    InMux I__4609 (
            .O(N__26339),
            .I(N__26135));
    InMux I__4608 (
            .O(N__26338),
            .I(N__26135));
    InMux I__4607 (
            .O(N__26337),
            .I(N__26124));
    InMux I__4606 (
            .O(N__26336),
            .I(N__26124));
    InMux I__4605 (
            .O(N__26335),
            .I(N__26124));
    InMux I__4604 (
            .O(N__26334),
            .I(N__26124));
    InMux I__4603 (
            .O(N__26333),
            .I(N__26124));
    LocalMux I__4602 (
            .O(N__26330),
            .I(N__26121));
    LocalMux I__4601 (
            .O(N__26327),
            .I(N__26118));
    LocalMux I__4600 (
            .O(N__26318),
            .I(N__26115));
    LocalMux I__4599 (
            .O(N__26307),
            .I(N__26106));
    Span4Mux_s3_h I__4598 (
            .O(N__26304),
            .I(N__26106));
    Span4Mux_v I__4597 (
            .O(N__26301),
            .I(N__26106));
    Span4Mux_v I__4596 (
            .O(N__26290),
            .I(N__26106));
    LocalMux I__4595 (
            .O(N__26285),
            .I(N__26095));
    Span4Mux_v I__4594 (
            .O(N__26282),
            .I(N__26095));
    Span4Mux_v I__4593 (
            .O(N__26279),
            .I(N__26095));
    Span4Mux_v I__4592 (
            .O(N__26270),
            .I(N__26095));
    Span4Mux_s2_h I__4591 (
            .O(N__26265),
            .I(N__26095));
    LocalMux I__4590 (
            .O(N__26260),
            .I(N__26086));
    Span4Mux_v I__4589 (
            .O(N__26255),
            .I(N__26086));
    Span4Mux_v I__4588 (
            .O(N__26250),
            .I(N__26086));
    Span4Mux_h I__4587 (
            .O(N__26241),
            .I(N__26086));
    LocalMux I__4586 (
            .O(N__26236),
            .I(n10725));
    LocalMux I__4585 (
            .O(N__26219),
            .I(n10725));
    LocalMux I__4584 (
            .O(N__26208),
            .I(n10725));
    LocalMux I__4583 (
            .O(N__26193),
            .I(n10725));
    LocalMux I__4582 (
            .O(N__26180),
            .I(n10725));
    LocalMux I__4581 (
            .O(N__26167),
            .I(n10725));
    LocalMux I__4580 (
            .O(N__26152),
            .I(n10725));
    LocalMux I__4579 (
            .O(N__26135),
            .I(n10725));
    LocalMux I__4578 (
            .O(N__26124),
            .I(n10725));
    Odrv4 I__4577 (
            .O(N__26121),
            .I(n10725));
    Odrv12 I__4576 (
            .O(N__26118),
            .I(n10725));
    Odrv4 I__4575 (
            .O(N__26115),
            .I(n10725));
    Odrv4 I__4574 (
            .O(N__26106),
            .I(n10725));
    Odrv4 I__4573 (
            .O(N__26095),
            .I(n10725));
    Odrv4 I__4572 (
            .O(N__26086),
            .I(n10725));
    InMux I__4571 (
            .O(N__26055),
            .I(N__26049));
    InMux I__4570 (
            .O(N__26054),
            .I(N__26046));
    InMux I__4569 (
            .O(N__26053),
            .I(N__26043));
    InMux I__4568 (
            .O(N__26052),
            .I(N__26039));
    LocalMux I__4567 (
            .O(N__26049),
            .I(N__26036));
    LocalMux I__4566 (
            .O(N__26046),
            .I(N__26033));
    LocalMux I__4565 (
            .O(N__26043),
            .I(N__26029));
    InMux I__4564 (
            .O(N__26042),
            .I(N__26026));
    LocalMux I__4563 (
            .O(N__26039),
            .I(N__26023));
    Span4Mux_v I__4562 (
            .O(N__26036),
            .I(N__26017));
    Span4Mux_h I__4561 (
            .O(N__26033),
            .I(N__26017));
    InMux I__4560 (
            .O(N__26032),
            .I(N__26014));
    Span4Mux_v I__4559 (
            .O(N__26029),
            .I(N__26011));
    LocalMux I__4558 (
            .O(N__26026),
            .I(N__26006));
    Span4Mux_h I__4557 (
            .O(N__26023),
            .I(N__26006));
    InMux I__4556 (
            .O(N__26022),
            .I(N__26003));
    Span4Mux_h I__4555 (
            .O(N__26017),
            .I(N__26000));
    LocalMux I__4554 (
            .O(N__26014),
            .I(N__25993));
    Span4Mux_h I__4553 (
            .O(N__26011),
            .I(N__25993));
    Span4Mux_v I__4552 (
            .O(N__26006),
            .I(N__25993));
    LocalMux I__4551 (
            .O(N__26003),
            .I(data_out_frame2_12_0));
    Odrv4 I__4550 (
            .O(N__26000),
            .I(data_out_frame2_12_0));
    Odrv4 I__4549 (
            .O(N__25993),
            .I(data_out_frame2_12_0));
    InMux I__4548 (
            .O(N__25986),
            .I(N__25978));
    InMux I__4547 (
            .O(N__25985),
            .I(N__25978));
    InMux I__4546 (
            .O(N__25984),
            .I(N__25975));
    InMux I__4545 (
            .O(N__25983),
            .I(N__25972));
    LocalMux I__4544 (
            .O(N__25978),
            .I(N__25969));
    LocalMux I__4543 (
            .O(N__25975),
            .I(N__25963));
    LocalMux I__4542 (
            .O(N__25972),
            .I(N__25963));
    Span4Mux_v I__4541 (
            .O(N__25969),
            .I(N__25959));
    InMux I__4540 (
            .O(N__25968),
            .I(N__25956));
    Span4Mux_v I__4539 (
            .O(N__25963),
            .I(N__25953));
    InMux I__4538 (
            .O(N__25962),
            .I(N__25950));
    Odrv4 I__4537 (
            .O(N__25959),
            .I(r_SM_Main_2_N_2031_1));
    LocalMux I__4536 (
            .O(N__25956),
            .I(r_SM_Main_2_N_2031_1));
    Odrv4 I__4535 (
            .O(N__25953),
            .I(r_SM_Main_2_N_2031_1));
    LocalMux I__4534 (
            .O(N__25950),
            .I(r_SM_Main_2_N_2031_1));
    InMux I__4533 (
            .O(N__25941),
            .I(N__25931));
    InMux I__4532 (
            .O(N__25940),
            .I(N__25928));
    InMux I__4531 (
            .O(N__25939),
            .I(N__25925));
    InMux I__4530 (
            .O(N__25938),
            .I(N__25920));
    InMux I__4529 (
            .O(N__25937),
            .I(N__25920));
    InMux I__4528 (
            .O(N__25936),
            .I(N__25917));
    InMux I__4527 (
            .O(N__25935),
            .I(N__25912));
    InMux I__4526 (
            .O(N__25934),
            .I(N__25912));
    LocalMux I__4525 (
            .O(N__25931),
            .I(N__25907));
    LocalMux I__4524 (
            .O(N__25928),
            .I(N__25907));
    LocalMux I__4523 (
            .O(N__25925),
            .I(N__25904));
    LocalMux I__4522 (
            .O(N__25920),
            .I(N__25901));
    LocalMux I__4521 (
            .O(N__25917),
            .I(N__25898));
    LocalMux I__4520 (
            .O(N__25912),
            .I(N__25893));
    Span4Mux_h I__4519 (
            .O(N__25907),
            .I(N__25893));
    Odrv4 I__4518 (
            .O(N__25904),
            .I(r_SM_Main_0));
    Odrv4 I__4517 (
            .O(N__25901),
            .I(r_SM_Main_0));
    Odrv4 I__4516 (
            .O(N__25898),
            .I(r_SM_Main_0));
    Odrv4 I__4515 (
            .O(N__25893),
            .I(r_SM_Main_0));
    InMux I__4514 (
            .O(N__25884),
            .I(N__25881));
    LocalMux I__4513 (
            .O(N__25881),
            .I(N__25878));
    Span4Mux_h I__4512 (
            .O(N__25878),
            .I(N__25875));
    Odrv4 I__4511 (
            .O(N__25875),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_12 ));
    CascadeMux I__4510 (
            .O(N__25872),
            .I(N__25869));
    InMux I__4509 (
            .O(N__25869),
            .I(N__25863));
    InMux I__4508 (
            .O(N__25868),
            .I(N__25858));
    InMux I__4507 (
            .O(N__25867),
            .I(N__25858));
    InMux I__4506 (
            .O(N__25866),
            .I(N__25855));
    LocalMux I__4505 (
            .O(N__25863),
            .I(N__25852));
    LocalMux I__4504 (
            .O(N__25858),
            .I(N__25849));
    LocalMux I__4503 (
            .O(N__25855),
            .I(N__25846));
    Span4Mux_h I__4502 (
            .O(N__25852),
            .I(N__25843));
    Span12Mux_v I__4501 (
            .O(N__25849),
            .I(N__25840));
    Odrv12 I__4500 (
            .O(N__25846),
            .I(\c0.FRAME_MATCHER_i_12 ));
    Odrv4 I__4499 (
            .O(N__25843),
            .I(\c0.FRAME_MATCHER_i_12 ));
    Odrv12 I__4498 (
            .O(N__25840),
            .I(\c0.FRAME_MATCHER_i_12 ));
    SRMux I__4497 (
            .O(N__25833),
            .I(N__25830));
    LocalMux I__4496 (
            .O(N__25830),
            .I(N__25827));
    Span4Mux_s2_v I__4495 (
            .O(N__25827),
            .I(N__25824));
    Span4Mux_v I__4494 (
            .O(N__25824),
            .I(N__25821));
    Odrv4 I__4493 (
            .O(N__25821),
            .I(\c0.n3_adj_2268 ));
    InMux I__4492 (
            .O(N__25818),
            .I(bfn_9_17_0_));
    InMux I__4491 (
            .O(N__25815),
            .I(\c0.n15972 ));
    InMux I__4490 (
            .O(N__25812),
            .I(\c0.n15973 ));
    InMux I__4489 (
            .O(N__25809),
            .I(\c0.n15974 ));
    InMux I__4488 (
            .O(N__25806),
            .I(N__25803));
    LocalMux I__4487 (
            .O(N__25803),
            .I(\c0.n17606 ));
    InMux I__4486 (
            .O(N__25800),
            .I(\c0.n15975 ));
    InMux I__4485 (
            .O(N__25797),
            .I(\c0.n15976 ));
    CascadeMux I__4484 (
            .O(N__25794),
            .I(N__25788));
    InMux I__4483 (
            .O(N__25793),
            .I(N__25785));
    CascadeMux I__4482 (
            .O(N__25792),
            .I(N__25782));
    InMux I__4481 (
            .O(N__25791),
            .I(N__25777));
    InMux I__4480 (
            .O(N__25788),
            .I(N__25777));
    LocalMux I__4479 (
            .O(N__25785),
            .I(N__25774));
    InMux I__4478 (
            .O(N__25782),
            .I(N__25768));
    LocalMux I__4477 (
            .O(N__25777),
            .I(N__25765));
    Span12Mux_s4_v I__4476 (
            .O(N__25774),
            .I(N__25762));
    InMux I__4475 (
            .O(N__25773),
            .I(N__25759));
    InMux I__4474 (
            .O(N__25772),
            .I(N__25754));
    InMux I__4473 (
            .O(N__25771),
            .I(N__25754));
    LocalMux I__4472 (
            .O(N__25768),
            .I(N__25749));
    Span4Mux_v I__4471 (
            .O(N__25765),
            .I(N__25749));
    Odrv12 I__4470 (
            .O(N__25762),
            .I(r_Bit_Index_1_adj_2441));
    LocalMux I__4469 (
            .O(N__25759),
            .I(r_Bit_Index_1_adj_2441));
    LocalMux I__4468 (
            .O(N__25754),
            .I(r_Bit_Index_1_adj_2441));
    Odrv4 I__4467 (
            .O(N__25749),
            .I(r_Bit_Index_1_adj_2441));
    InMux I__4466 (
            .O(N__25740),
            .I(N__25737));
    LocalMux I__4465 (
            .O(N__25737),
            .I(N__25731));
    InMux I__4464 (
            .O(N__25736),
            .I(N__25726));
    InMux I__4463 (
            .O(N__25735),
            .I(N__25721));
    InMux I__4462 (
            .O(N__25734),
            .I(N__25721));
    Span12Mux_s6_v I__4461 (
            .O(N__25731),
            .I(N__25718));
    InMux I__4460 (
            .O(N__25730),
            .I(N__25713));
    InMux I__4459 (
            .O(N__25729),
            .I(N__25713));
    LocalMux I__4458 (
            .O(N__25726),
            .I(N__25710));
    LocalMux I__4457 (
            .O(N__25721),
            .I(r_Bit_Index_0_adj_2442));
    Odrv12 I__4456 (
            .O(N__25718),
            .I(r_Bit_Index_0_adj_2442));
    LocalMux I__4455 (
            .O(N__25713),
            .I(r_Bit_Index_0_adj_2442));
    Odrv4 I__4454 (
            .O(N__25710),
            .I(r_Bit_Index_0_adj_2442));
    InMux I__4453 (
            .O(N__25701),
            .I(N__25698));
    LocalMux I__4452 (
            .O(N__25698),
            .I(N__25695));
    Span12Mux_v I__4451 (
            .O(N__25695),
            .I(N__25692));
    Odrv12 I__4450 (
            .O(N__25692),
            .I(n5266));
    IoInMux I__4449 (
            .O(N__25689),
            .I(N__25686));
    LocalMux I__4448 (
            .O(N__25686),
            .I(N__25683));
    Span4Mux_s3_v I__4447 (
            .O(N__25683),
            .I(N__25680));
    Odrv4 I__4446 (
            .O(N__25680),
            .I(tx_enable));
    CEMux I__4445 (
            .O(N__25677),
            .I(N__25673));
    CEMux I__4444 (
            .O(N__25676),
            .I(N__25669));
    LocalMux I__4443 (
            .O(N__25673),
            .I(N__25666));
    InMux I__4442 (
            .O(N__25672),
            .I(N__25663));
    LocalMux I__4441 (
            .O(N__25669),
            .I(N__25660));
    Span4Mux_v I__4440 (
            .O(N__25666),
            .I(N__25655));
    LocalMux I__4439 (
            .O(N__25663),
            .I(N__25655));
    Sp12to4 I__4438 (
            .O(N__25660),
            .I(N__25650));
    Sp12to4 I__4437 (
            .O(N__25655),
            .I(N__25650));
    Odrv12 I__4436 (
            .O(N__25650),
            .I(n10674));
    InMux I__4435 (
            .O(N__25647),
            .I(N__25644));
    LocalMux I__4434 (
            .O(N__25644),
            .I(N__25641));
    Odrv12 I__4433 (
            .O(N__25641),
            .I(\c0.n17574 ));
    InMux I__4432 (
            .O(N__25638),
            .I(N__25635));
    LocalMux I__4431 (
            .O(N__25635),
            .I(N__25632));
    Span4Mux_s2_v I__4430 (
            .O(N__25632),
            .I(N__25629));
    Odrv4 I__4429 (
            .O(N__25629),
            .I(\c0.rx.n10620 ));
    InMux I__4428 (
            .O(N__25626),
            .I(N__25620));
    InMux I__4427 (
            .O(N__25625),
            .I(N__25613));
    InMux I__4426 (
            .O(N__25624),
            .I(N__25613));
    InMux I__4425 (
            .O(N__25623),
            .I(N__25613));
    LocalMux I__4424 (
            .O(N__25620),
            .I(N__25608));
    LocalMux I__4423 (
            .O(N__25613),
            .I(N__25608));
    Span4Mux_s2_v I__4422 (
            .O(N__25608),
            .I(N__25605));
    Odrv4 I__4421 (
            .O(N__25605),
            .I(n17361));
    CascadeMux I__4420 (
            .O(N__25602),
            .I(N__25599));
    InMux I__4419 (
            .O(N__25599),
            .I(N__25595));
    InMux I__4418 (
            .O(N__25598),
            .I(N__25592));
    LocalMux I__4417 (
            .O(N__25595),
            .I(N__25588));
    LocalMux I__4416 (
            .O(N__25592),
            .I(N__25585));
    CascadeMux I__4415 (
            .O(N__25591),
            .I(N__25581));
    Span4Mux_s2_v I__4414 (
            .O(N__25588),
            .I(N__25578));
    Span4Mux_s2_v I__4413 (
            .O(N__25585),
            .I(N__25575));
    InMux I__4412 (
            .O(N__25584),
            .I(N__25570));
    InMux I__4411 (
            .O(N__25581),
            .I(N__25570));
    Odrv4 I__4410 (
            .O(N__25578),
            .I(\c0.rx.r_SM_Main_2_N_2088_2 ));
    Odrv4 I__4409 (
            .O(N__25575),
            .I(\c0.rx.r_SM_Main_2_N_2088_2 ));
    LocalMux I__4408 (
            .O(N__25570),
            .I(\c0.rx.r_SM_Main_2_N_2088_2 ));
    InMux I__4407 (
            .O(N__25563),
            .I(N__25553));
    InMux I__4406 (
            .O(N__25562),
            .I(N__25553));
    InMux I__4405 (
            .O(N__25561),
            .I(N__25553));
    CascadeMux I__4404 (
            .O(N__25560),
            .I(N__25547));
    LocalMux I__4403 (
            .O(N__25553),
            .I(N__25541));
    InMux I__4402 (
            .O(N__25552),
            .I(N__25534));
    InMux I__4401 (
            .O(N__25551),
            .I(N__25534));
    InMux I__4400 (
            .O(N__25550),
            .I(N__25534));
    InMux I__4399 (
            .O(N__25547),
            .I(N__25531));
    InMux I__4398 (
            .O(N__25546),
            .I(N__25524));
    InMux I__4397 (
            .O(N__25545),
            .I(N__25524));
    InMux I__4396 (
            .O(N__25544),
            .I(N__25524));
    Span4Mux_h I__4395 (
            .O(N__25541),
            .I(N__25521));
    LocalMux I__4394 (
            .O(N__25534),
            .I(r_SM_Main_1));
    LocalMux I__4393 (
            .O(N__25531),
            .I(r_SM_Main_1));
    LocalMux I__4392 (
            .O(N__25524),
            .I(r_SM_Main_1));
    Odrv4 I__4391 (
            .O(N__25521),
            .I(r_SM_Main_1));
    CascadeMux I__4390 (
            .O(N__25512),
            .I(\c0.rx.r_SM_Main_2_N_2088_2_cascade_ ));
    CascadeMux I__4389 (
            .O(N__25509),
            .I(N__25504));
    InMux I__4388 (
            .O(N__25508),
            .I(N__25499));
    InMux I__4387 (
            .O(N__25507),
            .I(N__25496));
    InMux I__4386 (
            .O(N__25504),
            .I(N__25489));
    InMux I__4385 (
            .O(N__25503),
            .I(N__25489));
    InMux I__4384 (
            .O(N__25502),
            .I(N__25489));
    LocalMux I__4383 (
            .O(N__25499),
            .I(N__25479));
    LocalMux I__4382 (
            .O(N__25496),
            .I(N__25479));
    LocalMux I__4381 (
            .O(N__25489),
            .I(N__25476));
    InMux I__4380 (
            .O(N__25488),
            .I(N__25469));
    InMux I__4379 (
            .O(N__25487),
            .I(N__25469));
    InMux I__4378 (
            .O(N__25486),
            .I(N__25469));
    InMux I__4377 (
            .O(N__25485),
            .I(N__25464));
    InMux I__4376 (
            .O(N__25484),
            .I(N__25464));
    Span4Mux_h I__4375 (
            .O(N__25479),
            .I(N__25461));
    Span4Mux_h I__4374 (
            .O(N__25476),
            .I(N__25458));
    LocalMux I__4373 (
            .O(N__25469),
            .I(\c0.rx.r_SM_Main_0 ));
    LocalMux I__4372 (
            .O(N__25464),
            .I(\c0.rx.r_SM_Main_0 ));
    Odrv4 I__4371 (
            .O(N__25461),
            .I(\c0.rx.r_SM_Main_0 ));
    Odrv4 I__4370 (
            .O(N__25458),
            .I(\c0.rx.r_SM_Main_0 ));
    SRMux I__4369 (
            .O(N__25449),
            .I(N__25446));
    LocalMux I__4368 (
            .O(N__25446),
            .I(N__25443));
    Span4Mux_v I__4367 (
            .O(N__25443),
            .I(N__25440));
    Odrv4 I__4366 (
            .O(N__25440),
            .I(\c0.n3_adj_2254 ));
    CascadeMux I__4365 (
            .O(N__25437),
            .I(N__25434));
    InMux I__4364 (
            .O(N__25434),
            .I(N__25426));
    InMux I__4363 (
            .O(N__25433),
            .I(N__25426));
    InMux I__4362 (
            .O(N__25432),
            .I(N__25423));
    InMux I__4361 (
            .O(N__25431),
            .I(N__25420));
    LocalMux I__4360 (
            .O(N__25426),
            .I(N__25417));
    LocalMux I__4359 (
            .O(N__25423),
            .I(N__25414));
    LocalMux I__4358 (
            .O(N__25420),
            .I(N__25411));
    Odrv4 I__4357 (
            .O(N__25417),
            .I(\c0.FRAME_MATCHER_i_18 ));
    Odrv12 I__4356 (
            .O(N__25414),
            .I(\c0.FRAME_MATCHER_i_18 ));
    Odrv4 I__4355 (
            .O(N__25411),
            .I(\c0.FRAME_MATCHER_i_18 ));
    InMux I__4354 (
            .O(N__25404),
            .I(N__25401));
    LocalMux I__4353 (
            .O(N__25401),
            .I(N__25398));
    Span4Mux_v I__4352 (
            .O(N__25398),
            .I(N__25395));
    Odrv4 I__4351 (
            .O(N__25395),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_18 ));
    SRMux I__4350 (
            .O(N__25392),
            .I(N__25389));
    LocalMux I__4349 (
            .O(N__25389),
            .I(N__25386));
    Span4Mux_v I__4348 (
            .O(N__25386),
            .I(N__25383));
    Span4Mux_h I__4347 (
            .O(N__25383),
            .I(N__25380));
    Odrv4 I__4346 (
            .O(N__25380),
            .I(\c0.n3_adj_2288 ));
    InMux I__4345 (
            .O(N__25377),
            .I(N__25374));
    LocalMux I__4344 (
            .O(N__25374),
            .I(N__25371));
    Span4Mux_h I__4343 (
            .O(N__25371),
            .I(N__25368));
    Span4Mux_h I__4342 (
            .O(N__25368),
            .I(N__25365));
    Odrv4 I__4341 (
            .O(N__25365),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_1 ));
    SRMux I__4340 (
            .O(N__25362),
            .I(N__25359));
    LocalMux I__4339 (
            .O(N__25359),
            .I(N__25356));
    Span4Mux_v I__4338 (
            .O(N__25356),
            .I(N__25353));
    Span4Mux_h I__4337 (
            .O(N__25353),
            .I(N__25350));
    Odrv4 I__4336 (
            .O(N__25350),
            .I(\c0.n3_adj_2246 ));
    CascadeMux I__4335 (
            .O(N__25347),
            .I(N__25344));
    InMux I__4334 (
            .O(N__25344),
            .I(N__25337));
    InMux I__4333 (
            .O(N__25343),
            .I(N__25337));
    CascadeMux I__4332 (
            .O(N__25342),
            .I(N__25334));
    LocalMux I__4331 (
            .O(N__25337),
            .I(N__25331));
    InMux I__4330 (
            .O(N__25334),
            .I(N__25328));
    Span4Mux_v I__4329 (
            .O(N__25331),
            .I(N__25322));
    LocalMux I__4328 (
            .O(N__25328),
            .I(N__25322));
    InMux I__4327 (
            .O(N__25327),
            .I(N__25319));
    Span4Mux_h I__4326 (
            .O(N__25322),
            .I(N__25316));
    LocalMux I__4325 (
            .O(N__25319),
            .I(\c0.FRAME_MATCHER_i_22 ));
    Odrv4 I__4324 (
            .O(N__25316),
            .I(\c0.FRAME_MATCHER_i_22 ));
    InMux I__4323 (
            .O(N__25311),
            .I(N__25308));
    LocalMux I__4322 (
            .O(N__25308),
            .I(N__25305));
    Span4Mux_v I__4321 (
            .O(N__25305),
            .I(N__25302));
    Odrv4 I__4320 (
            .O(N__25302),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_22 ));
    InMux I__4319 (
            .O(N__25299),
            .I(N__25295));
    InMux I__4318 (
            .O(N__25298),
            .I(N__25292));
    LocalMux I__4317 (
            .O(N__25295),
            .I(N__25289));
    LocalMux I__4316 (
            .O(N__25292),
            .I(N__25285));
    Span4Mux_h I__4315 (
            .O(N__25289),
            .I(N__25282));
    InMux I__4314 (
            .O(N__25288),
            .I(N__25278));
    Span4Mux_h I__4313 (
            .O(N__25285),
            .I(N__25275));
    Span4Mux_v I__4312 (
            .O(N__25282),
            .I(N__25272));
    InMux I__4311 (
            .O(N__25281),
            .I(N__25269));
    LocalMux I__4310 (
            .O(N__25278),
            .I(N__25266));
    Odrv4 I__4309 (
            .O(N__25275),
            .I(\c0.FRAME_MATCHER_i_26 ));
    Odrv4 I__4308 (
            .O(N__25272),
            .I(\c0.FRAME_MATCHER_i_26 ));
    LocalMux I__4307 (
            .O(N__25269),
            .I(\c0.FRAME_MATCHER_i_26 ));
    Odrv12 I__4306 (
            .O(N__25266),
            .I(\c0.FRAME_MATCHER_i_26 ));
    SRMux I__4305 (
            .O(N__25257),
            .I(N__25254));
    LocalMux I__4304 (
            .O(N__25254),
            .I(N__25251));
    Span4Mux_h I__4303 (
            .O(N__25251),
            .I(N__25248));
    Span4Mux_v I__4302 (
            .O(N__25248),
            .I(N__25245));
    Odrv4 I__4301 (
            .O(N__25245),
            .I(\c0.n3_adj_2238 ));
    InMux I__4300 (
            .O(N__25242),
            .I(N__25239));
    LocalMux I__4299 (
            .O(N__25239),
            .I(N__25236));
    Odrv4 I__4298 (
            .O(N__25236),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_10 ));
    InMux I__4297 (
            .O(N__25233),
            .I(N__25230));
    LocalMux I__4296 (
            .O(N__25230),
            .I(N__25227));
    Span4Mux_v I__4295 (
            .O(N__25227),
            .I(N__25224));
    Odrv4 I__4294 (
            .O(N__25224),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_26 ));
    CascadeMux I__4293 (
            .O(N__25221),
            .I(N__25215));
    InMux I__4292 (
            .O(N__25220),
            .I(N__25212));
    InMux I__4291 (
            .O(N__25219),
            .I(N__25207));
    InMux I__4290 (
            .O(N__25218),
            .I(N__25207));
    InMux I__4289 (
            .O(N__25215),
            .I(N__25204));
    LocalMux I__4288 (
            .O(N__25212),
            .I(N__25201));
    LocalMux I__4287 (
            .O(N__25207),
            .I(N__25198));
    LocalMux I__4286 (
            .O(N__25204),
            .I(N__25195));
    Span4Mux_h I__4285 (
            .O(N__25201),
            .I(N__25192));
    Span4Mux_h I__4284 (
            .O(N__25198),
            .I(N__25189));
    Odrv4 I__4283 (
            .O(N__25195),
            .I(\c0.FRAME_MATCHER_i_25 ));
    Odrv4 I__4282 (
            .O(N__25192),
            .I(\c0.FRAME_MATCHER_i_25 ));
    Odrv4 I__4281 (
            .O(N__25189),
            .I(\c0.FRAME_MATCHER_i_25 ));
    InMux I__4280 (
            .O(N__25182),
            .I(N__25179));
    LocalMux I__4279 (
            .O(N__25179),
            .I(N__25176));
    Span4Mux_v I__4278 (
            .O(N__25176),
            .I(N__25173));
    Odrv4 I__4277 (
            .O(N__25173),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_25 ));
    InMux I__4276 (
            .O(N__25170),
            .I(N__25166));
    InMux I__4275 (
            .O(N__25169),
            .I(N__25163));
    LocalMux I__4274 (
            .O(N__25166),
            .I(N__25160));
    LocalMux I__4273 (
            .O(N__25163),
            .I(N__25155));
    Span4Mux_h I__4272 (
            .O(N__25160),
            .I(N__25152));
    InMux I__4271 (
            .O(N__25159),
            .I(N__25147));
    InMux I__4270 (
            .O(N__25158),
            .I(N__25147));
    Odrv4 I__4269 (
            .O(N__25155),
            .I(\c0.FRAME_MATCHER_i_24 ));
    Odrv4 I__4268 (
            .O(N__25152),
            .I(\c0.FRAME_MATCHER_i_24 ));
    LocalMux I__4267 (
            .O(N__25147),
            .I(\c0.FRAME_MATCHER_i_24 ));
    InMux I__4266 (
            .O(N__25140),
            .I(N__25137));
    LocalMux I__4265 (
            .O(N__25137),
            .I(N__25134));
    Span4Mux_v I__4264 (
            .O(N__25134),
            .I(N__25131));
    Span4Mux_s3_h I__4263 (
            .O(N__25131),
            .I(N__25128));
    Odrv4 I__4262 (
            .O(N__25128),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_24 ));
    InMux I__4261 (
            .O(N__25125),
            .I(N__25121));
    CascadeMux I__4260 (
            .O(N__25124),
            .I(N__25116));
    LocalMux I__4259 (
            .O(N__25121),
            .I(N__25113));
    CascadeMux I__4258 (
            .O(N__25120),
            .I(N__25110));
    CascadeMux I__4257 (
            .O(N__25119),
            .I(N__25107));
    InMux I__4256 (
            .O(N__25116),
            .I(N__25104));
    Span4Mux_v I__4255 (
            .O(N__25113),
            .I(N__25101));
    InMux I__4254 (
            .O(N__25110),
            .I(N__25096));
    InMux I__4253 (
            .O(N__25107),
            .I(N__25096));
    LocalMux I__4252 (
            .O(N__25104),
            .I(N__25093));
    Span4Mux_v I__4251 (
            .O(N__25101),
            .I(N__25090));
    LocalMux I__4250 (
            .O(N__25096),
            .I(N__25087));
    Span4Mux_v I__4249 (
            .O(N__25093),
            .I(N__25082));
    Span4Mux_h I__4248 (
            .O(N__25090),
            .I(N__25082));
    Span4Mux_v I__4247 (
            .O(N__25087),
            .I(N__25079));
    Odrv4 I__4246 (
            .O(N__25082),
            .I(\c0.FRAME_MATCHER_i_23 ));
    Odrv4 I__4245 (
            .O(N__25079),
            .I(\c0.FRAME_MATCHER_i_23 ));
    InMux I__4244 (
            .O(N__25074),
            .I(N__25071));
    LocalMux I__4243 (
            .O(N__25071),
            .I(N__25068));
    Span4Mux_h I__4242 (
            .O(N__25068),
            .I(N__25065));
    Span4Mux_h I__4241 (
            .O(N__25065),
            .I(N__25062));
    Odrv4 I__4240 (
            .O(N__25062),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_23 ));
    InMux I__4239 (
            .O(N__25059),
            .I(N__25056));
    LocalMux I__4238 (
            .O(N__25056),
            .I(N__25050));
    InMux I__4237 (
            .O(N__25055),
            .I(N__25045));
    InMux I__4236 (
            .O(N__25054),
            .I(N__25045));
    InMux I__4235 (
            .O(N__25053),
            .I(N__25042));
    Span4Mux_v I__4234 (
            .O(N__25050),
            .I(N__25039));
    LocalMux I__4233 (
            .O(N__25045),
            .I(N__25036));
    LocalMux I__4232 (
            .O(N__25042),
            .I(N__25033));
    Span4Mux_h I__4231 (
            .O(N__25039),
            .I(N__25030));
    Span4Mux_h I__4230 (
            .O(N__25036),
            .I(N__25027));
    Odrv12 I__4229 (
            .O(N__25033),
            .I(\c0.FRAME_MATCHER_i_20 ));
    Odrv4 I__4228 (
            .O(N__25030),
            .I(\c0.FRAME_MATCHER_i_20 ));
    Odrv4 I__4227 (
            .O(N__25027),
            .I(\c0.FRAME_MATCHER_i_20 ));
    InMux I__4226 (
            .O(N__25020),
            .I(N__25017));
    LocalMux I__4225 (
            .O(N__25017),
            .I(N__25014));
    Span4Mux_h I__4224 (
            .O(N__25014),
            .I(N__25011));
    Odrv4 I__4223 (
            .O(N__25011),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_20 ));
    CascadeMux I__4222 (
            .O(N__25008),
            .I(N__25004));
    InMux I__4221 (
            .O(N__25007),
            .I(N__25001));
    InMux I__4220 (
            .O(N__25004),
            .I(N__24998));
    LocalMux I__4219 (
            .O(N__25001),
            .I(N__24995));
    LocalMux I__4218 (
            .O(N__24998),
            .I(N__24990));
    Span4Mux_v I__4217 (
            .O(N__24995),
            .I(N__24987));
    InMux I__4216 (
            .O(N__24994),
            .I(N__24982));
    InMux I__4215 (
            .O(N__24993),
            .I(N__24982));
    Span4Mux_h I__4214 (
            .O(N__24990),
            .I(N__24979));
    Sp12to4 I__4213 (
            .O(N__24987),
            .I(N__24974));
    LocalMux I__4212 (
            .O(N__24982),
            .I(N__24974));
    Odrv4 I__4211 (
            .O(N__24979),
            .I(\c0.FRAME_MATCHER_i_19 ));
    Odrv12 I__4210 (
            .O(N__24974),
            .I(\c0.FRAME_MATCHER_i_19 ));
    InMux I__4209 (
            .O(N__24969),
            .I(N__24966));
    LocalMux I__4208 (
            .O(N__24966),
            .I(N__24963));
    Span4Mux_h I__4207 (
            .O(N__24963),
            .I(N__24960));
    Span4Mux_h I__4206 (
            .O(N__24960),
            .I(N__24957));
    Odrv4 I__4205 (
            .O(N__24957),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_19 ));
    InMux I__4204 (
            .O(N__24954),
            .I(N__24951));
    LocalMux I__4203 (
            .O(N__24951),
            .I(N__24948));
    Span12Mux_s6_v I__4202 (
            .O(N__24948),
            .I(N__24945));
    Odrv12 I__4201 (
            .O(N__24945),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_16 ));
    InMux I__4200 (
            .O(N__24942),
            .I(N__24938));
    InMux I__4199 (
            .O(N__24941),
            .I(N__24933));
    LocalMux I__4198 (
            .O(N__24938),
            .I(N__24930));
    InMux I__4197 (
            .O(N__24937),
            .I(N__24927));
    InMux I__4196 (
            .O(N__24936),
            .I(N__24924));
    LocalMux I__4195 (
            .O(N__24933),
            .I(N__24921));
    Span4Mux_v I__4194 (
            .O(N__24930),
            .I(N__24916));
    LocalMux I__4193 (
            .O(N__24927),
            .I(N__24916));
    LocalMux I__4192 (
            .O(N__24924),
            .I(N__24912));
    Span4Mux_h I__4191 (
            .O(N__24921),
            .I(N__24909));
    Span4Mux_h I__4190 (
            .O(N__24916),
            .I(N__24906));
    InMux I__4189 (
            .O(N__24915),
            .I(N__24901));
    Span4Mux_h I__4188 (
            .O(N__24912),
            .I(N__24896));
    Span4Mux_v I__4187 (
            .O(N__24909),
            .I(N__24896));
    Span4Mux_v I__4186 (
            .O(N__24906),
            .I(N__24893));
    InMux I__4185 (
            .O(N__24905),
            .I(N__24888));
    InMux I__4184 (
            .O(N__24904),
            .I(N__24888));
    LocalMux I__4183 (
            .O(N__24901),
            .I(data_out_frame2_16_0));
    Odrv4 I__4182 (
            .O(N__24896),
            .I(data_out_frame2_16_0));
    Odrv4 I__4181 (
            .O(N__24893),
            .I(data_out_frame2_16_0));
    LocalMux I__4180 (
            .O(N__24888),
            .I(data_out_frame2_16_0));
    InMux I__4179 (
            .O(N__24879),
            .I(N__24876));
    LocalMux I__4178 (
            .O(N__24876),
            .I(N__24873));
    Span4Mux_v I__4177 (
            .O(N__24873),
            .I(N__24870));
    Span4Mux_h I__4176 (
            .O(N__24870),
            .I(N__24866));
    CascadeMux I__4175 (
            .O(N__24869),
            .I(N__24863));
    Span4Mux_v I__4174 (
            .O(N__24866),
            .I(N__24860));
    InMux I__4173 (
            .O(N__24863),
            .I(N__24857));
    Odrv4 I__4172 (
            .O(N__24860),
            .I(\c0.n17098 ));
    LocalMux I__4171 (
            .O(N__24857),
            .I(\c0.n17098 ));
    InMux I__4170 (
            .O(N__24852),
            .I(N__24847));
    InMux I__4169 (
            .O(N__24851),
            .I(N__24842));
    InMux I__4168 (
            .O(N__24850),
            .I(N__24839));
    LocalMux I__4167 (
            .O(N__24847),
            .I(N__24836));
    InMux I__4166 (
            .O(N__24846),
            .I(N__24833));
    InMux I__4165 (
            .O(N__24845),
            .I(N__24829));
    LocalMux I__4164 (
            .O(N__24842),
            .I(N__24826));
    LocalMux I__4163 (
            .O(N__24839),
            .I(N__24823));
    Span4Mux_v I__4162 (
            .O(N__24836),
            .I(N__24818));
    LocalMux I__4161 (
            .O(N__24833),
            .I(N__24818));
    InMux I__4160 (
            .O(N__24832),
            .I(N__24815));
    LocalMux I__4159 (
            .O(N__24829),
            .I(N__24812));
    Span4Mux_h I__4158 (
            .O(N__24826),
            .I(N__24805));
    Span4Mux_h I__4157 (
            .O(N__24823),
            .I(N__24805));
    Span4Mux_h I__4156 (
            .O(N__24818),
            .I(N__24805));
    LocalMux I__4155 (
            .O(N__24815),
            .I(data_out_frame2_8_3));
    Odrv4 I__4154 (
            .O(N__24812),
            .I(data_out_frame2_8_3));
    Odrv4 I__4153 (
            .O(N__24805),
            .I(data_out_frame2_8_3));
    InMux I__4152 (
            .O(N__24798),
            .I(N__24795));
    LocalMux I__4151 (
            .O(N__24795),
            .I(N__24792));
    Span4Mux_h I__4150 (
            .O(N__24792),
            .I(N__24789));
    Odrv4 I__4149 (
            .O(N__24789),
            .I(\c0.n17_adj_2321 ));
    CascadeMux I__4148 (
            .O(N__24786),
            .I(\c0.n30_cascade_ ));
    InMux I__4147 (
            .O(N__24783),
            .I(N__24779));
    InMux I__4146 (
            .O(N__24782),
            .I(N__24775));
    LocalMux I__4145 (
            .O(N__24779),
            .I(N__24771));
    InMux I__4144 (
            .O(N__24778),
            .I(N__24768));
    LocalMux I__4143 (
            .O(N__24775),
            .I(N__24765));
    InMux I__4142 (
            .O(N__24774),
            .I(N__24762));
    Span4Mux_h I__4141 (
            .O(N__24771),
            .I(N__24759));
    LocalMux I__4140 (
            .O(N__24768),
            .I(data_out_frame2_14_4));
    Odrv12 I__4139 (
            .O(N__24765),
            .I(data_out_frame2_14_4));
    LocalMux I__4138 (
            .O(N__24762),
            .I(data_out_frame2_14_4));
    Odrv4 I__4137 (
            .O(N__24759),
            .I(data_out_frame2_14_4));
    InMux I__4136 (
            .O(N__24750),
            .I(N__24745));
    InMux I__4135 (
            .O(N__24749),
            .I(N__24740));
    InMux I__4134 (
            .O(N__24748),
            .I(N__24737));
    LocalMux I__4133 (
            .O(N__24745),
            .I(N__24734));
    InMux I__4132 (
            .O(N__24744),
            .I(N__24731));
    InMux I__4131 (
            .O(N__24743),
            .I(N__24728));
    LocalMux I__4130 (
            .O(N__24740),
            .I(N__24725));
    LocalMux I__4129 (
            .O(N__24737),
            .I(N__24722));
    Span4Mux_v I__4128 (
            .O(N__24734),
            .I(N__24719));
    LocalMux I__4127 (
            .O(N__24731),
            .I(N__24716));
    LocalMux I__4126 (
            .O(N__24728),
            .I(data_out_frame2_11_0));
    Odrv4 I__4125 (
            .O(N__24725),
            .I(data_out_frame2_11_0));
    Odrv12 I__4124 (
            .O(N__24722),
            .I(data_out_frame2_11_0));
    Odrv4 I__4123 (
            .O(N__24719),
            .I(data_out_frame2_11_0));
    Odrv4 I__4122 (
            .O(N__24716),
            .I(data_out_frame2_11_0));
    InMux I__4121 (
            .O(N__24705),
            .I(N__24702));
    LocalMux I__4120 (
            .O(N__24702),
            .I(N__24699));
    Span4Mux_v I__4119 (
            .O(N__24699),
            .I(N__24695));
    InMux I__4118 (
            .O(N__24698),
            .I(N__24692));
    IoSpan4Mux I__4117 (
            .O(N__24695),
            .I(N__24689));
    LocalMux I__4116 (
            .O(N__24692),
            .I(N__24686));
    Span4Mux_s2_h I__4115 (
            .O(N__24689),
            .I(N__24681));
    Span4Mux_v I__4114 (
            .O(N__24686),
            .I(N__24681));
    Span4Mux_h I__4113 (
            .O(N__24681),
            .I(N__24678));
    Odrv4 I__4112 (
            .O(N__24678),
            .I(\c0.n17276 ));
    InMux I__4111 (
            .O(N__24675),
            .I(N__24669));
    InMux I__4110 (
            .O(N__24674),
            .I(N__24662));
    InMux I__4109 (
            .O(N__24673),
            .I(N__24662));
    InMux I__4108 (
            .O(N__24672),
            .I(N__24662));
    LocalMux I__4107 (
            .O(N__24669),
            .I(N__24657));
    LocalMux I__4106 (
            .O(N__24662),
            .I(N__24657));
    Odrv12 I__4105 (
            .O(N__24657),
            .I(n17412));
    CascadeMux I__4104 (
            .O(N__24654),
            .I(N__24648));
    InMux I__4103 (
            .O(N__24653),
            .I(N__24643));
    InMux I__4102 (
            .O(N__24652),
            .I(N__24643));
    InMux I__4101 (
            .O(N__24651),
            .I(N__24640));
    InMux I__4100 (
            .O(N__24648),
            .I(N__24637));
    LocalMux I__4099 (
            .O(N__24643),
            .I(N__24633));
    LocalMux I__4098 (
            .O(N__24640),
            .I(N__24630));
    LocalMux I__4097 (
            .O(N__24637),
            .I(N__24627));
    InMux I__4096 (
            .O(N__24636),
            .I(N__24624));
    Span4Mux_h I__4095 (
            .O(N__24633),
            .I(N__24621));
    Span4Mux_v I__4094 (
            .O(N__24630),
            .I(N__24616));
    Span4Mux_v I__4093 (
            .O(N__24627),
            .I(N__24616));
    LocalMux I__4092 (
            .O(N__24624),
            .I(data_out_frame2_9_3));
    Odrv4 I__4091 (
            .O(N__24621),
            .I(data_out_frame2_9_3));
    Odrv4 I__4090 (
            .O(N__24616),
            .I(data_out_frame2_9_3));
    InMux I__4089 (
            .O(N__24609),
            .I(N__24606));
    LocalMux I__4088 (
            .O(N__24606),
            .I(N__24603));
    Span4Mux_h I__4087 (
            .O(N__24603),
            .I(N__24600));
    Odrv4 I__4086 (
            .O(N__24600),
            .I(\c0.n6_adj_2197 ));
    InMux I__4085 (
            .O(N__24597),
            .I(N__24593));
    InMux I__4084 (
            .O(N__24596),
            .I(N__24590));
    LocalMux I__4083 (
            .O(N__24593),
            .I(N__24587));
    LocalMux I__4082 (
            .O(N__24590),
            .I(N__24584));
    Span4Mux_h I__4081 (
            .O(N__24587),
            .I(N__24579));
    Span4Mux_v I__4080 (
            .O(N__24584),
            .I(N__24576));
    InMux I__4079 (
            .O(N__24583),
            .I(N__24573));
    InMux I__4078 (
            .O(N__24582),
            .I(N__24570));
    Span4Mux_h I__4077 (
            .O(N__24579),
            .I(N__24567));
    Span4Mux_h I__4076 (
            .O(N__24576),
            .I(N__24562));
    LocalMux I__4075 (
            .O(N__24573),
            .I(N__24562));
    LocalMux I__4074 (
            .O(N__24570),
            .I(data_out_frame2_15_7));
    Odrv4 I__4073 (
            .O(N__24567),
            .I(data_out_frame2_15_7));
    Odrv4 I__4072 (
            .O(N__24562),
            .I(data_out_frame2_15_7));
    CascadeMux I__4071 (
            .O(N__24555),
            .I(N__24552));
    InMux I__4070 (
            .O(N__24552),
            .I(N__24548));
    InMux I__4069 (
            .O(N__24551),
            .I(N__24545));
    LocalMux I__4068 (
            .O(N__24548),
            .I(N__24542));
    LocalMux I__4067 (
            .O(N__24545),
            .I(N__24539));
    Span4Mux_h I__4066 (
            .O(N__24542),
            .I(N__24536));
    Span4Mux_h I__4065 (
            .O(N__24539),
            .I(N__24533));
    Odrv4 I__4064 (
            .O(N__24536),
            .I(\c0.n17123 ));
    Odrv4 I__4063 (
            .O(N__24533),
            .I(\c0.n17123 ));
    InMux I__4062 (
            .O(N__24528),
            .I(N__24522));
    InMux I__4061 (
            .O(N__24527),
            .I(N__24519));
    InMux I__4060 (
            .O(N__24526),
            .I(N__24516));
    InMux I__4059 (
            .O(N__24525),
            .I(N__24513));
    LocalMux I__4058 (
            .O(N__24522),
            .I(N__24510));
    LocalMux I__4057 (
            .O(N__24519),
            .I(N__24507));
    LocalMux I__4056 (
            .O(N__24516),
            .I(data_out_frame2_14_6));
    LocalMux I__4055 (
            .O(N__24513),
            .I(data_out_frame2_14_6));
    Odrv12 I__4054 (
            .O(N__24510),
            .I(data_out_frame2_14_6));
    Odrv4 I__4053 (
            .O(N__24507),
            .I(data_out_frame2_14_6));
    InMux I__4052 (
            .O(N__24498),
            .I(N__24495));
    LocalMux I__4051 (
            .O(N__24495),
            .I(N__24492));
    Span4Mux_v I__4050 (
            .O(N__24492),
            .I(N__24489));
    Span4Mux_h I__4049 (
            .O(N__24489),
            .I(N__24486));
    Odrv4 I__4048 (
            .O(N__24486),
            .I(\c0.n10434 ));
    InMux I__4047 (
            .O(N__24483),
            .I(N__24478));
    InMux I__4046 (
            .O(N__24482),
            .I(N__24475));
    InMux I__4045 (
            .O(N__24481),
            .I(N__24472));
    LocalMux I__4044 (
            .O(N__24478),
            .I(N__24468));
    LocalMux I__4043 (
            .O(N__24475),
            .I(N__24465));
    LocalMux I__4042 (
            .O(N__24472),
            .I(N__24461));
    InMux I__4041 (
            .O(N__24471),
            .I(N__24458));
    Span4Mux_v I__4040 (
            .O(N__24468),
            .I(N__24453));
    Span4Mux_s3_h I__4039 (
            .O(N__24465),
            .I(N__24453));
    InMux I__4038 (
            .O(N__24464),
            .I(N__24450));
    Span4Mux_h I__4037 (
            .O(N__24461),
            .I(N__24447));
    LocalMux I__4036 (
            .O(N__24458),
            .I(N__24442));
    Span4Mux_h I__4035 (
            .O(N__24453),
            .I(N__24442));
    LocalMux I__4034 (
            .O(N__24450),
            .I(data_out_frame2_16_3));
    Odrv4 I__4033 (
            .O(N__24447),
            .I(data_out_frame2_16_3));
    Odrv4 I__4032 (
            .O(N__24442),
            .I(data_out_frame2_16_3));
    InMux I__4031 (
            .O(N__24435),
            .I(N__24430));
    InMux I__4030 (
            .O(N__24434),
            .I(N__24427));
    CascadeMux I__4029 (
            .O(N__24433),
            .I(N__24423));
    LocalMux I__4028 (
            .O(N__24430),
            .I(N__24419));
    LocalMux I__4027 (
            .O(N__24427),
            .I(N__24416));
    InMux I__4026 (
            .O(N__24426),
            .I(N__24411));
    InMux I__4025 (
            .O(N__24423),
            .I(N__24411));
    InMux I__4024 (
            .O(N__24422),
            .I(N__24408));
    Span4Mux_v I__4023 (
            .O(N__24419),
            .I(N__24401));
    Span4Mux_v I__4022 (
            .O(N__24416),
            .I(N__24401));
    LocalMux I__4021 (
            .O(N__24411),
            .I(N__24401));
    LocalMux I__4020 (
            .O(N__24408),
            .I(data_out_frame2_15_3));
    Odrv4 I__4019 (
            .O(N__24401),
            .I(data_out_frame2_15_3));
    InMux I__4018 (
            .O(N__24396),
            .I(N__24393));
    LocalMux I__4017 (
            .O(N__24393),
            .I(N__24390));
    Span4Mux_s3_h I__4016 (
            .O(N__24390),
            .I(N__24387));
    Span4Mux_h I__4015 (
            .O(N__24387),
            .I(N__24384));
    Odrv4 I__4014 (
            .O(N__24384),
            .I(\c0.n10482 ));
    InMux I__4013 (
            .O(N__24381),
            .I(N__24377));
    InMux I__4012 (
            .O(N__24380),
            .I(N__24374));
    LocalMux I__4011 (
            .O(N__24377),
            .I(N__24371));
    LocalMux I__4010 (
            .O(N__24374),
            .I(N__24368));
    Span4Mux_s3_h I__4009 (
            .O(N__24371),
            .I(N__24362));
    Span4Mux_h I__4008 (
            .O(N__24368),
            .I(N__24362));
    InMux I__4007 (
            .O(N__24367),
            .I(N__24359));
    Span4Mux_v I__4006 (
            .O(N__24362),
            .I(N__24354));
    LocalMux I__4005 (
            .O(N__24359),
            .I(N__24351));
    InMux I__4004 (
            .O(N__24358),
            .I(N__24347));
    InMux I__4003 (
            .O(N__24357),
            .I(N__24344));
    Span4Mux_s3_h I__4002 (
            .O(N__24354),
            .I(N__24339));
    Span4Mux_v I__4001 (
            .O(N__24351),
            .I(N__24339));
    InMux I__4000 (
            .O(N__24350),
            .I(N__24336));
    LocalMux I__3999 (
            .O(N__24347),
            .I(data_out_frame2_8_4));
    LocalMux I__3998 (
            .O(N__24344),
            .I(data_out_frame2_8_4));
    Odrv4 I__3997 (
            .O(N__24339),
            .I(data_out_frame2_8_4));
    LocalMux I__3996 (
            .O(N__24336),
            .I(data_out_frame2_8_4));
    InMux I__3995 (
            .O(N__24327),
            .I(N__24324));
    LocalMux I__3994 (
            .O(N__24324),
            .I(N__24320));
    InMux I__3993 (
            .O(N__24323),
            .I(N__24317));
    Span4Mux_s2_h I__3992 (
            .O(N__24320),
            .I(N__24312));
    LocalMux I__3991 (
            .O(N__24317),
            .I(N__24309));
    InMux I__3990 (
            .O(N__24316),
            .I(N__24305));
    InMux I__3989 (
            .O(N__24315),
            .I(N__24302));
    Span4Mux_h I__3988 (
            .O(N__24312),
            .I(N__24299));
    Span4Mux_v I__3987 (
            .O(N__24309),
            .I(N__24296));
    InMux I__3986 (
            .O(N__24308),
            .I(N__24293));
    LocalMux I__3985 (
            .O(N__24305),
            .I(data_out_frame2_8_0));
    LocalMux I__3984 (
            .O(N__24302),
            .I(data_out_frame2_8_0));
    Odrv4 I__3983 (
            .O(N__24299),
            .I(data_out_frame2_8_0));
    Odrv4 I__3982 (
            .O(N__24296),
            .I(data_out_frame2_8_0));
    LocalMux I__3981 (
            .O(N__24293),
            .I(data_out_frame2_8_0));
    InMux I__3980 (
            .O(N__24282),
            .I(N__24279));
    LocalMux I__3979 (
            .O(N__24279),
            .I(N__24276));
    Odrv12 I__3978 (
            .O(N__24276),
            .I(\c0.n10513 ));
    CEMux I__3977 (
            .O(N__24273),
            .I(N__24266));
    CEMux I__3976 (
            .O(N__24272),
            .I(N__24261));
    CEMux I__3975 (
            .O(N__24271),
            .I(N__24258));
    CEMux I__3974 (
            .O(N__24270),
            .I(N__24255));
    CEMux I__3973 (
            .O(N__24269),
            .I(N__24251));
    LocalMux I__3972 (
            .O(N__24266),
            .I(N__24248));
    CEMux I__3971 (
            .O(N__24265),
            .I(N__24245));
    CEMux I__3970 (
            .O(N__24264),
            .I(N__24242));
    LocalMux I__3969 (
            .O(N__24261),
            .I(N__24239));
    LocalMux I__3968 (
            .O(N__24258),
            .I(N__24236));
    LocalMux I__3967 (
            .O(N__24255),
            .I(N__24233));
    CEMux I__3966 (
            .O(N__24254),
            .I(N__24230));
    LocalMux I__3965 (
            .O(N__24251),
            .I(N__24227));
    Span4Mux_v I__3964 (
            .O(N__24248),
            .I(N__24224));
    LocalMux I__3963 (
            .O(N__24245),
            .I(N__24221));
    LocalMux I__3962 (
            .O(N__24242),
            .I(N__24218));
    Span4Mux_s3_h I__3961 (
            .O(N__24239),
            .I(N__24209));
    Span4Mux_v I__3960 (
            .O(N__24236),
            .I(N__24209));
    Span4Mux_s3_h I__3959 (
            .O(N__24233),
            .I(N__24209));
    LocalMux I__3958 (
            .O(N__24230),
            .I(N__24209));
    Sp12to4 I__3957 (
            .O(N__24227),
            .I(N__24206));
    Span4Mux_h I__3956 (
            .O(N__24224),
            .I(N__24201));
    Span4Mux_v I__3955 (
            .O(N__24221),
            .I(N__24201));
    Span4Mux_v I__3954 (
            .O(N__24218),
            .I(N__24198));
    Span4Mux_h I__3953 (
            .O(N__24209),
            .I(N__24195));
    Span12Mux_v I__3952 (
            .O(N__24206),
            .I(N__24192));
    Sp12to4 I__3951 (
            .O(N__24201),
            .I(N__24189));
    Span4Mux_h I__3950 (
            .O(N__24198),
            .I(N__24184));
    Span4Mux_h I__3949 (
            .O(N__24195),
            .I(N__24184));
    Odrv12 I__3948 (
            .O(N__24192),
            .I(\c0.tx2.n9269 ));
    Odrv12 I__3947 (
            .O(N__24189),
            .I(\c0.tx2.n9269 ));
    Odrv4 I__3946 (
            .O(N__24184),
            .I(\c0.tx2.n9269 ));
    CascadeMux I__3945 (
            .O(N__24177),
            .I(N__24173));
    InMux I__3944 (
            .O(N__24176),
            .I(N__24170));
    InMux I__3943 (
            .O(N__24173),
            .I(N__24167));
    LocalMux I__3942 (
            .O(N__24170),
            .I(N__24164));
    LocalMux I__3941 (
            .O(N__24167),
            .I(N__24160));
    Span4Mux_h I__3940 (
            .O(N__24164),
            .I(N__24157));
    InMux I__3939 (
            .O(N__24163),
            .I(N__24153));
    Span4Mux_v I__3938 (
            .O(N__24160),
            .I(N__24148));
    Span4Mux_v I__3937 (
            .O(N__24157),
            .I(N__24148));
    InMux I__3936 (
            .O(N__24156),
            .I(N__24145));
    LocalMux I__3935 (
            .O(N__24153),
            .I(data_out_frame2_5_2));
    Odrv4 I__3934 (
            .O(N__24148),
            .I(data_out_frame2_5_2));
    LocalMux I__3933 (
            .O(N__24145),
            .I(data_out_frame2_5_2));
    CascadeMux I__3932 (
            .O(N__24138),
            .I(N__24134));
    InMux I__3931 (
            .O(N__24137),
            .I(N__24130));
    InMux I__3930 (
            .O(N__24134),
            .I(N__24126));
    InMux I__3929 (
            .O(N__24133),
            .I(N__24123));
    LocalMux I__3928 (
            .O(N__24130),
            .I(N__24120));
    InMux I__3927 (
            .O(N__24129),
            .I(N__24117));
    LocalMux I__3926 (
            .O(N__24126),
            .I(N__24114));
    LocalMux I__3925 (
            .O(N__24123),
            .I(data_out_frame2_10_4));
    Odrv4 I__3924 (
            .O(N__24120),
            .I(data_out_frame2_10_4));
    LocalMux I__3923 (
            .O(N__24117),
            .I(data_out_frame2_10_4));
    Odrv4 I__3922 (
            .O(N__24114),
            .I(data_out_frame2_10_4));
    InMux I__3921 (
            .O(N__24105),
            .I(N__24102));
    LocalMux I__3920 (
            .O(N__24102),
            .I(N__24099));
    Span4Mux_s2_h I__3919 (
            .O(N__24099),
            .I(N__24095));
    InMux I__3918 (
            .O(N__24098),
            .I(N__24092));
    Span4Mux_h I__3917 (
            .O(N__24095),
            .I(N__24089));
    LocalMux I__3916 (
            .O(N__24092),
            .I(N__24086));
    Odrv4 I__3915 (
            .O(N__24089),
            .I(\c0.n10456 ));
    Odrv12 I__3914 (
            .O(N__24086),
            .I(\c0.n10456 ));
    InMux I__3913 (
            .O(N__24081),
            .I(N__24074));
    InMux I__3912 (
            .O(N__24080),
            .I(N__24074));
    InMux I__3911 (
            .O(N__24079),
            .I(N__24070));
    LocalMux I__3910 (
            .O(N__24074),
            .I(N__24067));
    CascadeMux I__3909 (
            .O(N__24073),
            .I(N__24064));
    LocalMux I__3908 (
            .O(N__24070),
            .I(N__24060));
    Span4Mux_v I__3907 (
            .O(N__24067),
            .I(N__24057));
    InMux I__3906 (
            .O(N__24064),
            .I(N__24054));
    InMux I__3905 (
            .O(N__24063),
            .I(N__24051));
    Span4Mux_h I__3904 (
            .O(N__24060),
            .I(N__24048));
    Sp12to4 I__3903 (
            .O(N__24057),
            .I(N__24043));
    LocalMux I__3902 (
            .O(N__24054),
            .I(N__24043));
    LocalMux I__3901 (
            .O(N__24051),
            .I(data_out_frame2_10_5));
    Odrv4 I__3900 (
            .O(N__24048),
            .I(data_out_frame2_10_5));
    Odrv12 I__3899 (
            .O(N__24043),
            .I(data_out_frame2_10_5));
    InMux I__3898 (
            .O(N__24036),
            .I(N__24033));
    LocalMux I__3897 (
            .O(N__24033),
            .I(N__24028));
    InMux I__3896 (
            .O(N__24032),
            .I(N__24025));
    InMux I__3895 (
            .O(N__24031),
            .I(N__24021));
    Span4Mux_h I__3894 (
            .O(N__24028),
            .I(N__24018));
    LocalMux I__3893 (
            .O(N__24025),
            .I(N__24015));
    InMux I__3892 (
            .O(N__24024),
            .I(N__24012));
    LocalMux I__3891 (
            .O(N__24021),
            .I(data_out_frame2_11_3));
    Odrv4 I__3890 (
            .O(N__24018),
            .I(data_out_frame2_11_3));
    Odrv12 I__3889 (
            .O(N__24015),
            .I(data_out_frame2_11_3));
    LocalMux I__3888 (
            .O(N__24012),
            .I(data_out_frame2_11_3));
    CascadeMux I__3887 (
            .O(N__24003),
            .I(N__24000));
    InMux I__3886 (
            .O(N__24000),
            .I(N__23996));
    InMux I__3885 (
            .O(N__23999),
            .I(N__23993));
    LocalMux I__3884 (
            .O(N__23996),
            .I(N__23989));
    LocalMux I__3883 (
            .O(N__23993),
            .I(N__23986));
    InMux I__3882 (
            .O(N__23992),
            .I(N__23982));
    Span4Mux_h I__3881 (
            .O(N__23989),
            .I(N__23979));
    Span4Mux_h I__3880 (
            .O(N__23986),
            .I(N__23976));
    InMux I__3879 (
            .O(N__23985),
            .I(N__23973));
    LocalMux I__3878 (
            .O(N__23982),
            .I(data_out_frame2_14_1));
    Odrv4 I__3877 (
            .O(N__23979),
            .I(data_out_frame2_14_1));
    Odrv4 I__3876 (
            .O(N__23976),
            .I(data_out_frame2_14_1));
    LocalMux I__3875 (
            .O(N__23973),
            .I(data_out_frame2_14_1));
    InMux I__3874 (
            .O(N__23964),
            .I(N__23961));
    LocalMux I__3873 (
            .O(N__23961),
            .I(N__23955));
    InMux I__3872 (
            .O(N__23960),
            .I(N__23952));
    InMux I__3871 (
            .O(N__23959),
            .I(N__23949));
    InMux I__3870 (
            .O(N__23958),
            .I(N__23946));
    Span4Mux_h I__3869 (
            .O(N__23955),
            .I(N__23943));
    LocalMux I__3868 (
            .O(N__23952),
            .I(N__23940));
    LocalMux I__3867 (
            .O(N__23949),
            .I(data_out_frame2_15_1));
    LocalMux I__3866 (
            .O(N__23946),
            .I(data_out_frame2_15_1));
    Odrv4 I__3865 (
            .O(N__23943),
            .I(data_out_frame2_15_1));
    Odrv4 I__3864 (
            .O(N__23940),
            .I(data_out_frame2_15_1));
    InMux I__3863 (
            .O(N__23931),
            .I(N__23928));
    LocalMux I__3862 (
            .O(N__23928),
            .I(N__23925));
    Odrv4 I__3861 (
            .O(N__23925),
            .I(\c0.n18016 ));
    CascadeMux I__3860 (
            .O(N__23922),
            .I(N__23919));
    InMux I__3859 (
            .O(N__23919),
            .I(N__23911));
    InMux I__3858 (
            .O(N__23918),
            .I(N__23911));
    InMux I__3857 (
            .O(N__23917),
            .I(N__23907));
    InMux I__3856 (
            .O(N__23916),
            .I(N__23904));
    LocalMux I__3855 (
            .O(N__23911),
            .I(N__23899));
    InMux I__3854 (
            .O(N__23910),
            .I(N__23896));
    LocalMux I__3853 (
            .O(N__23907),
            .I(N__23893));
    LocalMux I__3852 (
            .O(N__23904),
            .I(N__23890));
    InMux I__3851 (
            .O(N__23903),
            .I(N__23887));
    InMux I__3850 (
            .O(N__23902),
            .I(N__23884));
    Span4Mux_v I__3849 (
            .O(N__23899),
            .I(N__23881));
    LocalMux I__3848 (
            .O(N__23896),
            .I(N__23878));
    Span4Mux_s3_h I__3847 (
            .O(N__23893),
            .I(N__23873));
    Span4Mux_v I__3846 (
            .O(N__23890),
            .I(N__23873));
    LocalMux I__3845 (
            .O(N__23887),
            .I(N__23870));
    LocalMux I__3844 (
            .O(N__23884),
            .I(data_out_frame2_12_2));
    Odrv4 I__3843 (
            .O(N__23881),
            .I(data_out_frame2_12_2));
    Odrv12 I__3842 (
            .O(N__23878),
            .I(data_out_frame2_12_2));
    Odrv4 I__3841 (
            .O(N__23873),
            .I(data_out_frame2_12_2));
    Odrv4 I__3840 (
            .O(N__23870),
            .I(data_out_frame2_12_2));
    InMux I__3839 (
            .O(N__23859),
            .I(N__23856));
    LocalMux I__3838 (
            .O(N__23856),
            .I(N__23853));
    Span4Mux_v I__3837 (
            .O(N__23853),
            .I(N__23848));
    InMux I__3836 (
            .O(N__23852),
            .I(N__23845));
    InMux I__3835 (
            .O(N__23851),
            .I(N__23841));
    Span4Mux_h I__3834 (
            .O(N__23848),
            .I(N__23836));
    LocalMux I__3833 (
            .O(N__23845),
            .I(N__23836));
    InMux I__3832 (
            .O(N__23844),
            .I(N__23833));
    LocalMux I__3831 (
            .O(N__23841),
            .I(N__23830));
    Span4Mux_h I__3830 (
            .O(N__23836),
            .I(N__23827));
    LocalMux I__3829 (
            .O(N__23833),
            .I(data_out_frame2_7_2));
    Odrv4 I__3828 (
            .O(N__23830),
            .I(data_out_frame2_7_2));
    Odrv4 I__3827 (
            .O(N__23827),
            .I(data_out_frame2_7_2));
    InMux I__3826 (
            .O(N__23820),
            .I(N__23816));
    InMux I__3825 (
            .O(N__23819),
            .I(N__23811));
    LocalMux I__3824 (
            .O(N__23816),
            .I(N__23808));
    InMux I__3823 (
            .O(N__23815),
            .I(N__23805));
    InMux I__3822 (
            .O(N__23814),
            .I(N__23802));
    LocalMux I__3821 (
            .O(N__23811),
            .I(N__23799));
    Span4Mux_v I__3820 (
            .O(N__23808),
            .I(N__23794));
    LocalMux I__3819 (
            .O(N__23805),
            .I(N__23794));
    LocalMux I__3818 (
            .O(N__23802),
            .I(data_out_frame2_6_2));
    Odrv4 I__3817 (
            .O(N__23799),
            .I(data_out_frame2_6_2));
    Odrv4 I__3816 (
            .O(N__23794),
            .I(data_out_frame2_6_2));
    InMux I__3815 (
            .O(N__23787),
            .I(N__23784));
    LocalMux I__3814 (
            .O(N__23784),
            .I(N__23781));
    Span4Mux_v I__3813 (
            .O(N__23781),
            .I(N__23778));
    Span4Mux_v I__3812 (
            .O(N__23778),
            .I(N__23775));
    Odrv4 I__3811 (
            .O(N__23775),
            .I(\c0.n5_adj_2290 ));
    CascadeMux I__3810 (
            .O(N__23772),
            .I(N__23768));
    InMux I__3809 (
            .O(N__23771),
            .I(N__23763));
    InMux I__3808 (
            .O(N__23768),
            .I(N__23763));
    LocalMux I__3807 (
            .O(N__23763),
            .I(N__23759));
    InMux I__3806 (
            .O(N__23762),
            .I(N__23756));
    Span4Mux_h I__3805 (
            .O(N__23759),
            .I(N__23751));
    LocalMux I__3804 (
            .O(N__23756),
            .I(N__23751));
    Odrv4 I__3803 (
            .O(N__23751),
            .I(\c0.n10563 ));
    CascadeMux I__3802 (
            .O(N__23748),
            .I(N__23745));
    InMux I__3801 (
            .O(N__23745),
            .I(N__23741));
    InMux I__3800 (
            .O(N__23744),
            .I(N__23738));
    LocalMux I__3799 (
            .O(N__23741),
            .I(N__23735));
    LocalMux I__3798 (
            .O(N__23738),
            .I(N__23732));
    Span4Mux_v I__3797 (
            .O(N__23735),
            .I(N__23729));
    Span4Mux_h I__3796 (
            .O(N__23732),
            .I(N__23726));
    Span4Mux_h I__3795 (
            .O(N__23729),
            .I(N__23718));
    Span4Mux_v I__3794 (
            .O(N__23726),
            .I(N__23718));
    InMux I__3793 (
            .O(N__23725),
            .I(N__23715));
    InMux I__3792 (
            .O(N__23724),
            .I(N__23712));
    InMux I__3791 (
            .O(N__23723),
            .I(N__23709));
    Span4Mux_h I__3790 (
            .O(N__23718),
            .I(N__23706));
    LocalMux I__3789 (
            .O(N__23715),
            .I(N__23703));
    LocalMux I__3788 (
            .O(N__23712),
            .I(data_out_frame2_13_5));
    LocalMux I__3787 (
            .O(N__23709),
            .I(data_out_frame2_13_5));
    Odrv4 I__3786 (
            .O(N__23706),
            .I(data_out_frame2_13_5));
    Odrv4 I__3785 (
            .O(N__23703),
            .I(data_out_frame2_13_5));
    InMux I__3784 (
            .O(N__23694),
            .I(N__23691));
    LocalMux I__3783 (
            .O(N__23691),
            .I(N__23688));
    Span4Mux_v I__3782 (
            .O(N__23688),
            .I(N__23684));
    InMux I__3781 (
            .O(N__23687),
            .I(N__23681));
    Odrv4 I__3780 (
            .O(N__23684),
            .I(\c0.n17095 ));
    LocalMux I__3779 (
            .O(N__23681),
            .I(\c0.n17095 ));
    InMux I__3778 (
            .O(N__23676),
            .I(N__23673));
    LocalMux I__3777 (
            .O(N__23673),
            .I(N__23670));
    Odrv12 I__3776 (
            .O(N__23670),
            .I(\c0.n31 ));
    InMux I__3775 (
            .O(N__23667),
            .I(N__23663));
    InMux I__3774 (
            .O(N__23666),
            .I(N__23660));
    LocalMux I__3773 (
            .O(N__23663),
            .I(N__23655));
    LocalMux I__3772 (
            .O(N__23660),
            .I(N__23655));
    Span4Mux_v I__3771 (
            .O(N__23655),
            .I(N__23649));
    InMux I__3770 (
            .O(N__23654),
            .I(N__23646));
    CascadeMux I__3769 (
            .O(N__23653),
            .I(N__23643));
    InMux I__3768 (
            .O(N__23652),
            .I(N__23640));
    Span4Mux_s3_h I__3767 (
            .O(N__23649),
            .I(N__23637));
    LocalMux I__3766 (
            .O(N__23646),
            .I(N__23634));
    InMux I__3765 (
            .O(N__23643),
            .I(N__23631));
    LocalMux I__3764 (
            .O(N__23640),
            .I(data_out_frame2_13_1));
    Odrv4 I__3763 (
            .O(N__23637),
            .I(data_out_frame2_13_1));
    Odrv12 I__3762 (
            .O(N__23634),
            .I(data_out_frame2_13_1));
    LocalMux I__3761 (
            .O(N__23631),
            .I(data_out_frame2_13_1));
    InMux I__3760 (
            .O(N__23622),
            .I(N__23618));
    InMux I__3759 (
            .O(N__23621),
            .I(N__23615));
    LocalMux I__3758 (
            .O(N__23618),
            .I(N__23609));
    LocalMux I__3757 (
            .O(N__23615),
            .I(N__23606));
    InMux I__3756 (
            .O(N__23614),
            .I(N__23603));
    InMux I__3755 (
            .O(N__23613),
            .I(N__23599));
    InMux I__3754 (
            .O(N__23612),
            .I(N__23596));
    Span4Mux_v I__3753 (
            .O(N__23609),
            .I(N__23589));
    Span4Mux_v I__3752 (
            .O(N__23606),
            .I(N__23589));
    LocalMux I__3751 (
            .O(N__23603),
            .I(N__23589));
    InMux I__3750 (
            .O(N__23602),
            .I(N__23586));
    LocalMux I__3749 (
            .O(N__23599),
            .I(data_out_frame2_12_1));
    LocalMux I__3748 (
            .O(N__23596),
            .I(data_out_frame2_12_1));
    Odrv4 I__3747 (
            .O(N__23589),
            .I(data_out_frame2_12_1));
    LocalMux I__3746 (
            .O(N__23586),
            .I(data_out_frame2_12_1));
    InMux I__3745 (
            .O(N__23577),
            .I(N__23574));
    LocalMux I__3744 (
            .O(N__23574),
            .I(N__23571));
    Span4Mux_v I__3743 (
            .O(N__23571),
            .I(N__23568));
    Odrv4 I__3742 (
            .O(N__23568),
            .I(\c0.n18019 ));
    InMux I__3741 (
            .O(N__23565),
            .I(N__23558));
    InMux I__3740 (
            .O(N__23564),
            .I(N__23558));
    CascadeMux I__3739 (
            .O(N__23563),
            .I(N__23555));
    LocalMux I__3738 (
            .O(N__23558),
            .I(N__23551));
    InMux I__3737 (
            .O(N__23555),
            .I(N__23548));
    InMux I__3736 (
            .O(N__23554),
            .I(N__23543));
    Span4Mux_h I__3735 (
            .O(N__23551),
            .I(N__23540));
    LocalMux I__3734 (
            .O(N__23548),
            .I(N__23537));
    InMux I__3733 (
            .O(N__23547),
            .I(N__23532));
    InMux I__3732 (
            .O(N__23546),
            .I(N__23532));
    LocalMux I__3731 (
            .O(N__23543),
            .I(data_out_frame2_12_3));
    Odrv4 I__3730 (
            .O(N__23540),
            .I(data_out_frame2_12_3));
    Odrv12 I__3729 (
            .O(N__23537),
            .I(data_out_frame2_12_3));
    LocalMux I__3728 (
            .O(N__23532),
            .I(data_out_frame2_12_3));
    InMux I__3727 (
            .O(N__23523),
            .I(N__23519));
    CascadeMux I__3726 (
            .O(N__23522),
            .I(N__23516));
    LocalMux I__3725 (
            .O(N__23519),
            .I(N__23513));
    InMux I__3724 (
            .O(N__23516),
            .I(N__23510));
    Span4Mux_v I__3723 (
            .O(N__23513),
            .I(N__23505));
    LocalMux I__3722 (
            .O(N__23510),
            .I(N__23505));
    Span4Mux_h I__3721 (
            .O(N__23505),
            .I(N__23500));
    InMux I__3720 (
            .O(N__23504),
            .I(N__23495));
    InMux I__3719 (
            .O(N__23503),
            .I(N__23495));
    Odrv4 I__3718 (
            .O(N__23500),
            .I(data_out_frame2_5_3));
    LocalMux I__3717 (
            .O(N__23495),
            .I(data_out_frame2_5_3));
    InMux I__3716 (
            .O(N__23490),
            .I(N__23487));
    LocalMux I__3715 (
            .O(N__23487),
            .I(\c0.n18142 ));
    InMux I__3714 (
            .O(N__23484),
            .I(N__23479));
    CascadeMux I__3713 (
            .O(N__23483),
            .I(N__23476));
    CascadeMux I__3712 (
            .O(N__23482),
            .I(N__23472));
    LocalMux I__3711 (
            .O(N__23479),
            .I(N__23469));
    InMux I__3710 (
            .O(N__23476),
            .I(N__23462));
    InMux I__3709 (
            .O(N__23475),
            .I(N__23462));
    InMux I__3708 (
            .O(N__23472),
            .I(N__23462));
    Span4Mux_h I__3707 (
            .O(N__23469),
            .I(N__23459));
    LocalMux I__3706 (
            .O(N__23462),
            .I(data_out_frame2_8_7));
    Odrv4 I__3705 (
            .O(N__23459),
            .I(data_out_frame2_8_7));
    InMux I__3704 (
            .O(N__23454),
            .I(N__23450));
    InMux I__3703 (
            .O(N__23453),
            .I(N__23444));
    LocalMux I__3702 (
            .O(N__23450),
            .I(N__23441));
    CascadeMux I__3701 (
            .O(N__23449),
            .I(N__23438));
    InMux I__3700 (
            .O(N__23448),
            .I(N__23435));
    InMux I__3699 (
            .O(N__23447),
            .I(N__23432));
    LocalMux I__3698 (
            .O(N__23444),
            .I(N__23429));
    Span12Mux_v I__3697 (
            .O(N__23441),
            .I(N__23426));
    InMux I__3696 (
            .O(N__23438),
            .I(N__23423));
    LocalMux I__3695 (
            .O(N__23435),
            .I(data_out_frame2_9_7));
    LocalMux I__3694 (
            .O(N__23432),
            .I(data_out_frame2_9_7));
    Odrv4 I__3693 (
            .O(N__23429),
            .I(data_out_frame2_9_7));
    Odrv12 I__3692 (
            .O(N__23426),
            .I(data_out_frame2_9_7));
    LocalMux I__3691 (
            .O(N__23423),
            .I(data_out_frame2_9_7));
    InMux I__3690 (
            .O(N__23412),
            .I(N__23409));
    LocalMux I__3689 (
            .O(N__23409),
            .I(N__23406));
    Span4Mux_s2_h I__3688 (
            .O(N__23406),
            .I(N__23403));
    Span4Mux_h I__3687 (
            .O(N__23403),
            .I(N__23400));
    Odrv4 I__3686 (
            .O(N__23400),
            .I(\c0.n18145 ));
    InMux I__3685 (
            .O(N__23397),
            .I(N__23393));
    InMux I__3684 (
            .O(N__23396),
            .I(N__23390));
    LocalMux I__3683 (
            .O(N__23393),
            .I(N__23385));
    LocalMux I__3682 (
            .O(N__23390),
            .I(N__23382));
    InMux I__3681 (
            .O(N__23389),
            .I(N__23378));
    CascadeMux I__3680 (
            .O(N__23388),
            .I(N__23375));
    Span4Mux_v I__3679 (
            .O(N__23385),
            .I(N__23370));
    Span4Mux_v I__3678 (
            .O(N__23382),
            .I(N__23370));
    InMux I__3677 (
            .O(N__23381),
            .I(N__23367));
    LocalMux I__3676 (
            .O(N__23378),
            .I(N__23364));
    InMux I__3675 (
            .O(N__23375),
            .I(N__23361));
    Span4Mux_h I__3674 (
            .O(N__23370),
            .I(N__23358));
    LocalMux I__3673 (
            .O(N__23367),
            .I(data_out_frame2_5_1));
    Odrv12 I__3672 (
            .O(N__23364),
            .I(data_out_frame2_5_1));
    LocalMux I__3671 (
            .O(N__23361),
            .I(data_out_frame2_5_1));
    Odrv4 I__3670 (
            .O(N__23358),
            .I(data_out_frame2_5_1));
    InMux I__3669 (
            .O(N__23349),
            .I(N__23346));
    LocalMux I__3668 (
            .O(N__23346),
            .I(N__23343));
    Span12Mux_v I__3667 (
            .O(N__23343),
            .I(N__23340));
    Odrv12 I__3666 (
            .O(N__23340),
            .I(\c0.n6_adj_2142 ));
    InMux I__3665 (
            .O(N__23337),
            .I(N__23334));
    LocalMux I__3664 (
            .O(N__23334),
            .I(N__23331));
    Span4Mux_h I__3663 (
            .O(N__23331),
            .I(N__23328));
    Span4Mux_h I__3662 (
            .O(N__23328),
            .I(N__23325));
    Odrv4 I__3661 (
            .O(N__23325),
            .I(\c0.n18064 ));
    InMux I__3660 (
            .O(N__23322),
            .I(N__23319));
    LocalMux I__3659 (
            .O(N__23319),
            .I(\c0.n18067 ));
    InMux I__3658 (
            .O(N__23316),
            .I(N__23313));
    LocalMux I__3657 (
            .O(N__23313),
            .I(N__23310));
    Odrv4 I__3656 (
            .O(N__23310),
            .I(n8191));
    InMux I__3655 (
            .O(N__23307),
            .I(N__23304));
    LocalMux I__3654 (
            .O(N__23304),
            .I(N__23300));
    InMux I__3653 (
            .O(N__23303),
            .I(N__23297));
    Span4Mux_h I__3652 (
            .O(N__23300),
            .I(N__23292));
    LocalMux I__3651 (
            .O(N__23297),
            .I(N__23289));
    InMux I__3650 (
            .O(N__23296),
            .I(N__23286));
    InMux I__3649 (
            .O(N__23295),
            .I(N__23283));
    Span4Mux_v I__3648 (
            .O(N__23292),
            .I(N__23280));
    Span4Mux_v I__3647 (
            .O(N__23289),
            .I(N__23275));
    LocalMux I__3646 (
            .O(N__23286),
            .I(N__23275));
    LocalMux I__3645 (
            .O(N__23283),
            .I(data_out_frame2_6_1));
    Odrv4 I__3644 (
            .O(N__23280),
            .I(data_out_frame2_6_1));
    Odrv4 I__3643 (
            .O(N__23275),
            .I(data_out_frame2_6_1));
    InMux I__3642 (
            .O(N__23268),
            .I(N__23265));
    LocalMux I__3641 (
            .O(N__23265),
            .I(\c0.n5_adj_2289 ));
    InMux I__3640 (
            .O(N__23262),
            .I(N__23256));
    InMux I__3639 (
            .O(N__23261),
            .I(N__23250));
    InMux I__3638 (
            .O(N__23260),
            .I(N__23250));
    InMux I__3637 (
            .O(N__23259),
            .I(N__23247));
    LocalMux I__3636 (
            .O(N__23256),
            .I(N__23244));
    InMux I__3635 (
            .O(N__23255),
            .I(N__23241));
    LocalMux I__3634 (
            .O(N__23250),
            .I(N__23234));
    LocalMux I__3633 (
            .O(N__23247),
            .I(N__23234));
    Span4Mux_v I__3632 (
            .O(N__23244),
            .I(N__23229));
    LocalMux I__3631 (
            .O(N__23241),
            .I(N__23229));
    InMux I__3630 (
            .O(N__23240),
            .I(N__23226));
    InMux I__3629 (
            .O(N__23239),
            .I(N__23223));
    Span4Mux_v I__3628 (
            .O(N__23234),
            .I(N__23218));
    Span4Mux_h I__3627 (
            .O(N__23229),
            .I(N__23218));
    LocalMux I__3626 (
            .O(N__23226),
            .I(data_out_frame2_11_7));
    LocalMux I__3625 (
            .O(N__23223),
            .I(data_out_frame2_11_7));
    Odrv4 I__3624 (
            .O(N__23218),
            .I(data_out_frame2_11_7));
    CascadeMux I__3623 (
            .O(N__23211),
            .I(\c0.n10413_cascade_ ));
    InMux I__3622 (
            .O(N__23208),
            .I(N__23202));
    InMux I__3621 (
            .O(N__23207),
            .I(N__23202));
    LocalMux I__3620 (
            .O(N__23202),
            .I(N__23199));
    Span4Mux_s2_h I__3619 (
            .O(N__23199),
            .I(N__23196));
    Span4Mux_h I__3618 (
            .O(N__23196),
            .I(N__23193));
    Odrv4 I__3617 (
            .O(N__23193),
            .I(\c0.n17282 ));
    InMux I__3616 (
            .O(N__23190),
            .I(N__23187));
    LocalMux I__3615 (
            .O(N__23187),
            .I(N__23181));
    InMux I__3614 (
            .O(N__23186),
            .I(N__23177));
    InMux I__3613 (
            .O(N__23185),
            .I(N__23174));
    InMux I__3612 (
            .O(N__23184),
            .I(N__23171));
    Span4Mux_h I__3611 (
            .O(N__23181),
            .I(N__23168));
    InMux I__3610 (
            .O(N__23180),
            .I(N__23165));
    LocalMux I__3609 (
            .O(N__23177),
            .I(N__23160));
    LocalMux I__3608 (
            .O(N__23174),
            .I(N__23160));
    LocalMux I__3607 (
            .O(N__23171),
            .I(data_out_frame2_10_6));
    Odrv4 I__3606 (
            .O(N__23168),
            .I(data_out_frame2_10_6));
    LocalMux I__3605 (
            .O(N__23165),
            .I(data_out_frame2_10_6));
    Odrv12 I__3604 (
            .O(N__23160),
            .I(data_out_frame2_10_6));
    CascadeMux I__3603 (
            .O(N__23151),
            .I(N__23147));
    InMux I__3602 (
            .O(N__23150),
            .I(N__23144));
    InMux I__3601 (
            .O(N__23147),
            .I(N__23141));
    LocalMux I__3600 (
            .O(N__23144),
            .I(N__23138));
    LocalMux I__3599 (
            .O(N__23141),
            .I(N__23131));
    Span4Mux_v I__3598 (
            .O(N__23138),
            .I(N__23131));
    InMux I__3597 (
            .O(N__23137),
            .I(N__23128));
    InMux I__3596 (
            .O(N__23136),
            .I(N__23125));
    Sp12to4 I__3595 (
            .O(N__23131),
            .I(N__23120));
    LocalMux I__3594 (
            .O(N__23128),
            .I(N__23115));
    LocalMux I__3593 (
            .O(N__23125),
            .I(N__23115));
    InMux I__3592 (
            .O(N__23124),
            .I(N__23110));
    InMux I__3591 (
            .O(N__23123),
            .I(N__23110));
    Odrv12 I__3590 (
            .O(N__23120),
            .I(data_out_frame2_11_6));
    Odrv4 I__3589 (
            .O(N__23115),
            .I(data_out_frame2_11_6));
    LocalMux I__3588 (
            .O(N__23110),
            .I(data_out_frame2_11_6));
    InMux I__3587 (
            .O(N__23103),
            .I(N__23100));
    LocalMux I__3586 (
            .O(N__23100),
            .I(\c0.n18124 ));
    InMux I__3585 (
            .O(N__23097),
            .I(N__23094));
    LocalMux I__3584 (
            .O(N__23094),
            .I(N__23091));
    Span4Mux_h I__3583 (
            .O(N__23091),
            .I(N__23088));
    Odrv4 I__3582 (
            .O(N__23088),
            .I(\c0.data_out_frame2_19_0 ));
    InMux I__3581 (
            .O(N__23085),
            .I(N__23081));
    InMux I__3580 (
            .O(N__23084),
            .I(N__23078));
    LocalMux I__3579 (
            .O(N__23081),
            .I(data_out_frame2_18_0));
    LocalMux I__3578 (
            .O(N__23078),
            .I(data_out_frame2_18_0));
    InMux I__3577 (
            .O(N__23073),
            .I(N__23070));
    LocalMux I__3576 (
            .O(N__23070),
            .I(N__23067));
    Odrv4 I__3575 (
            .O(N__23067),
            .I(\c0.n18160 ));
    CascadeMux I__3574 (
            .O(N__23064),
            .I(\c0.tx2.n13614_cascade_ ));
    InMux I__3573 (
            .O(N__23061),
            .I(N__23058));
    LocalMux I__3572 (
            .O(N__23058),
            .I(N__23055));
    Span4Mux_v I__3571 (
            .O(N__23055),
            .I(N__23052));
    Span4Mux_h I__3570 (
            .O(N__23052),
            .I(N__23049));
    Odrv4 I__3569 (
            .O(N__23049),
            .I(\c0.n17587 ));
    CascadeMux I__3568 (
            .O(N__23046),
            .I(N__23042));
    InMux I__3567 (
            .O(N__23045),
            .I(N__23039));
    InMux I__3566 (
            .O(N__23042),
            .I(N__23036));
    LocalMux I__3565 (
            .O(N__23039),
            .I(N__23031));
    LocalMux I__3564 (
            .O(N__23036),
            .I(N__23031));
    Span4Mux_h I__3563 (
            .O(N__23031),
            .I(N__23028));
    Odrv4 I__3562 (
            .O(N__23028),
            .I(\c0.n17107 ));
    InMux I__3561 (
            .O(N__23025),
            .I(N__23020));
    InMux I__3560 (
            .O(N__23024),
            .I(N__23016));
    CascadeMux I__3559 (
            .O(N__23023),
            .I(N__23013));
    LocalMux I__3558 (
            .O(N__23020),
            .I(N__23009));
    InMux I__3557 (
            .O(N__23019),
            .I(N__23006));
    LocalMux I__3556 (
            .O(N__23016),
            .I(N__23003));
    InMux I__3555 (
            .O(N__23013),
            .I(N__23000));
    InMux I__3554 (
            .O(N__23012),
            .I(N__22997));
    Span4Mux_h I__3553 (
            .O(N__23009),
            .I(N__22994));
    LocalMux I__3552 (
            .O(N__23006),
            .I(N__22991));
    Span4Mux_h I__3551 (
            .O(N__23003),
            .I(N__22988));
    LocalMux I__3550 (
            .O(N__23000),
            .I(N__22985));
    LocalMux I__3549 (
            .O(N__22997),
            .I(data_out_frame2_15_6));
    Odrv4 I__3548 (
            .O(N__22994),
            .I(data_out_frame2_15_6));
    Odrv12 I__3547 (
            .O(N__22991),
            .I(data_out_frame2_15_6));
    Odrv4 I__3546 (
            .O(N__22988),
            .I(data_out_frame2_15_6));
    Odrv4 I__3545 (
            .O(N__22985),
            .I(data_out_frame2_15_6));
    InMux I__3544 (
            .O(N__22974),
            .I(N__22969));
    InMux I__3543 (
            .O(N__22973),
            .I(N__22966));
    InMux I__3542 (
            .O(N__22972),
            .I(N__22963));
    LocalMux I__3541 (
            .O(N__22969),
            .I(N__22959));
    LocalMux I__3540 (
            .O(N__22966),
            .I(N__22954));
    LocalMux I__3539 (
            .O(N__22963),
            .I(N__22954));
    InMux I__3538 (
            .O(N__22962),
            .I(N__22951));
    Span4Mux_v I__3537 (
            .O(N__22959),
            .I(N__22946));
    Span4Mux_v I__3536 (
            .O(N__22954),
            .I(N__22946));
    LocalMux I__3535 (
            .O(N__22951),
            .I(data_out_frame2_12_6));
    Odrv4 I__3534 (
            .O(N__22946),
            .I(data_out_frame2_12_6));
    CascadeMux I__3533 (
            .O(N__22941),
            .I(\c0.n18118_cascade_ ));
    InMux I__3532 (
            .O(N__22938),
            .I(N__22934));
    InMux I__3531 (
            .O(N__22937),
            .I(N__22931));
    LocalMux I__3530 (
            .O(N__22934),
            .I(N__22928));
    LocalMux I__3529 (
            .O(N__22931),
            .I(N__22922));
    Span4Mux_h I__3528 (
            .O(N__22928),
            .I(N__22922));
    InMux I__3527 (
            .O(N__22927),
            .I(N__22918));
    Span4Mux_v I__3526 (
            .O(N__22922),
            .I(N__22915));
    InMux I__3525 (
            .O(N__22921),
            .I(N__22912));
    LocalMux I__3524 (
            .O(N__22918),
            .I(data_out_frame2_13_6));
    Odrv4 I__3523 (
            .O(N__22915),
            .I(data_out_frame2_13_6));
    LocalMux I__3522 (
            .O(N__22912),
            .I(data_out_frame2_13_6));
    CascadeMux I__3521 (
            .O(N__22905),
            .I(N__22902));
    InMux I__3520 (
            .O(N__22902),
            .I(N__22899));
    LocalMux I__3519 (
            .O(N__22899),
            .I(N__22896));
    Span4Mux_h I__3518 (
            .O(N__22896),
            .I(N__22893));
    Odrv4 I__3517 (
            .O(N__22893),
            .I(\c0.n18121 ));
    InMux I__3516 (
            .O(N__22890),
            .I(N__22887));
    LocalMux I__3515 (
            .O(N__22887),
            .I(N__22884));
    Odrv4 I__3514 (
            .O(N__22884),
            .I(\c0.tx2.n13614 ));
    InMux I__3513 (
            .O(N__22881),
            .I(N__22875));
    InMux I__3512 (
            .O(N__22880),
            .I(N__22875));
    LocalMux I__3511 (
            .O(N__22875),
            .I(n10976));
    CascadeMux I__3510 (
            .O(N__22872),
            .I(n10976_cascade_));
    InMux I__3509 (
            .O(N__22869),
            .I(N__22864));
    InMux I__3508 (
            .O(N__22868),
            .I(N__22859));
    InMux I__3507 (
            .O(N__22867),
            .I(N__22859));
    LocalMux I__3506 (
            .O(N__22864),
            .I(r_Bit_Index_2_adj_2440));
    LocalMux I__3505 (
            .O(N__22859),
            .I(r_Bit_Index_2_adj_2440));
    InMux I__3504 (
            .O(N__22854),
            .I(N__22849));
    InMux I__3503 (
            .O(N__22853),
            .I(N__22844));
    InMux I__3502 (
            .O(N__22852),
            .I(N__22844));
    LocalMux I__3501 (
            .O(N__22849),
            .I(\c0.rx.r_SM_Main_2_N_2094_0 ));
    LocalMux I__3500 (
            .O(N__22844),
            .I(\c0.rx.r_SM_Main_2_N_2094_0 ));
    InMux I__3499 (
            .O(N__22839),
            .I(N__22836));
    LocalMux I__3498 (
            .O(N__22836),
            .I(\c0.rx.n6_adj_2130 ));
    InMux I__3497 (
            .O(N__22833),
            .I(N__22830));
    LocalMux I__3496 (
            .O(N__22830),
            .I(\c0.n18247 ));
    CascadeMux I__3495 (
            .O(N__22827),
            .I(N__22824));
    InMux I__3494 (
            .O(N__22824),
            .I(N__22821));
    LocalMux I__3493 (
            .O(N__22821),
            .I(N__22818));
    Span4Mux_h I__3492 (
            .O(N__22818),
            .I(N__22815));
    Odrv4 I__3491 (
            .O(N__22815),
            .I(\c0.n22_adj_2372 ));
    InMux I__3490 (
            .O(N__22812),
            .I(N__22809));
    LocalMux I__3489 (
            .O(N__22809),
            .I(\c0.tx2.r_Tx_Data_2 ));
    InMux I__3488 (
            .O(N__22806),
            .I(N__22803));
    LocalMux I__3487 (
            .O(N__22803),
            .I(N__22800));
    Span4Mux_h I__3486 (
            .O(N__22800),
            .I(N__22797));
    Odrv4 I__3485 (
            .O(N__22797),
            .I(\c0.n17620 ));
    InMux I__3484 (
            .O(N__22794),
            .I(N__22791));
    LocalMux I__3483 (
            .O(N__22791),
            .I(N__22788));
    Span12Mux_v I__3482 (
            .O(N__22788),
            .I(N__22785));
    Odrv12 I__3481 (
            .O(N__22785),
            .I(\c0.tx2.r_Tx_Data_6 ));
    CascadeMux I__3480 (
            .O(N__22782),
            .I(N__22779));
    InMux I__3479 (
            .O(N__22779),
            .I(N__22776));
    LocalMux I__3478 (
            .O(N__22776),
            .I(N__22773));
    Span4Mux_h I__3477 (
            .O(N__22773),
            .I(N__22770));
    Span4Mux_h I__3476 (
            .O(N__22770),
            .I(N__22767));
    Odrv4 I__3475 (
            .O(N__22767),
            .I(\c0.tx2.r_Tx_Data_7 ));
    InMux I__3474 (
            .O(N__22764),
            .I(N__22761));
    LocalMux I__3473 (
            .O(N__22761),
            .I(N__22758));
    Span4Mux_v I__3472 (
            .O(N__22758),
            .I(N__22755));
    Span4Mux_h I__3471 (
            .O(N__22755),
            .I(N__22752));
    Odrv4 I__3470 (
            .O(N__22752),
            .I(\c0.tx2.r_Tx_Data_4 ));
    CascadeMux I__3469 (
            .O(N__22749),
            .I(\c0.tx2.n18082_cascade_ ));
    InMux I__3468 (
            .O(N__22746),
            .I(N__22743));
    LocalMux I__3467 (
            .O(N__22743),
            .I(N__22740));
    Span4Mux_h I__3466 (
            .O(N__22740),
            .I(N__22737));
    Span4Mux_h I__3465 (
            .O(N__22737),
            .I(N__22734));
    Odrv4 I__3464 (
            .O(N__22734),
            .I(\c0.tx2.r_Tx_Data_5 ));
    CascadeMux I__3463 (
            .O(N__22731),
            .I(\c0.tx2.n18085_cascade_ ));
    InMux I__3462 (
            .O(N__22728),
            .I(N__22725));
    LocalMux I__3461 (
            .O(N__22725),
            .I(\c0.tx2.n18235 ));
    CascadeMux I__3460 (
            .O(N__22722),
            .I(\c0.tx2.o_Tx_Serial_N_2062_cascade_ ));
    InMux I__3459 (
            .O(N__22719),
            .I(N__22716));
    LocalMux I__3458 (
            .O(N__22716),
            .I(N__22713));
    Span4Mux_v I__3457 (
            .O(N__22713),
            .I(N__22710));
    Odrv4 I__3456 (
            .O(N__22710),
            .I(n3));
    InMux I__3455 (
            .O(N__22707),
            .I(N__22704));
    LocalMux I__3454 (
            .O(N__22704),
            .I(N__22701));
    Odrv4 I__3453 (
            .O(N__22701),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_27 ));
    CascadeMux I__3452 (
            .O(N__22698),
            .I(N__22695));
    InMux I__3451 (
            .O(N__22695),
            .I(N__22690));
    InMux I__3450 (
            .O(N__22694),
            .I(N__22687));
    CascadeMux I__3449 (
            .O(N__22693),
            .I(N__22684));
    LocalMux I__3448 (
            .O(N__22690),
            .I(N__22680));
    LocalMux I__3447 (
            .O(N__22687),
            .I(N__22677));
    InMux I__3446 (
            .O(N__22684),
            .I(N__22672));
    InMux I__3445 (
            .O(N__22683),
            .I(N__22672));
    Sp12to4 I__3444 (
            .O(N__22680),
            .I(N__22669));
    Span4Mux_h I__3443 (
            .O(N__22677),
            .I(N__22666));
    LocalMux I__3442 (
            .O(N__22672),
            .I(\c0.FRAME_MATCHER_i_27 ));
    Odrv12 I__3441 (
            .O(N__22669),
            .I(\c0.FRAME_MATCHER_i_27 ));
    Odrv4 I__3440 (
            .O(N__22666),
            .I(\c0.FRAME_MATCHER_i_27 ));
    SRMux I__3439 (
            .O(N__22659),
            .I(N__22656));
    LocalMux I__3438 (
            .O(N__22656),
            .I(N__22653));
    Span4Mux_v I__3437 (
            .O(N__22653),
            .I(N__22650));
    Span4Mux_s2_v I__3436 (
            .O(N__22650),
            .I(N__22647));
    Odrv4 I__3435 (
            .O(N__22647),
            .I(\c0.n3_adj_2236 ));
    InMux I__3434 (
            .O(N__22644),
            .I(N__22641));
    LocalMux I__3433 (
            .O(N__22641),
            .I(N__22638));
    Span4Mux_v I__3432 (
            .O(N__22638),
            .I(N__22635));
    Odrv4 I__3431 (
            .O(N__22635),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_9 ));
    InMux I__3430 (
            .O(N__22632),
            .I(N__22627));
    InMux I__3429 (
            .O(N__22631),
            .I(N__22621));
    InMux I__3428 (
            .O(N__22630),
            .I(N__22621));
    LocalMux I__3427 (
            .O(N__22627),
            .I(N__22618));
    InMux I__3426 (
            .O(N__22626),
            .I(N__22615));
    LocalMux I__3425 (
            .O(N__22621),
            .I(N__22612));
    Span4Mux_h I__3424 (
            .O(N__22618),
            .I(N__22609));
    LocalMux I__3423 (
            .O(N__22615),
            .I(N__22606));
    Odrv4 I__3422 (
            .O(N__22612),
            .I(\c0.FRAME_MATCHER_i_9 ));
    Odrv4 I__3421 (
            .O(N__22609),
            .I(\c0.FRAME_MATCHER_i_9 ));
    Odrv12 I__3420 (
            .O(N__22606),
            .I(\c0.FRAME_MATCHER_i_9 ));
    SRMux I__3419 (
            .O(N__22599),
            .I(N__22596));
    LocalMux I__3418 (
            .O(N__22596),
            .I(N__22593));
    Span4Mux_h I__3417 (
            .O(N__22593),
            .I(N__22590));
    Odrv4 I__3416 (
            .O(N__22590),
            .I(\c0.n3_adj_2274 ));
    InMux I__3415 (
            .O(N__22587),
            .I(N__22584));
    LocalMux I__3414 (
            .O(N__22584),
            .I(\c0.rx.n17636 ));
    InMux I__3413 (
            .O(N__22581),
            .I(N__22578));
    LocalMux I__3412 (
            .O(N__22578),
            .I(n17707));
    InMux I__3411 (
            .O(N__22575),
            .I(N__22571));
    InMux I__3410 (
            .O(N__22574),
            .I(N__22568));
    LocalMux I__3409 (
            .O(N__22571),
            .I(N__22565));
    LocalMux I__3408 (
            .O(N__22568),
            .I(\c0.rx.r_Clock_Count_2 ));
    Odrv4 I__3407 (
            .O(N__22565),
            .I(\c0.rx.r_Clock_Count_2 ));
    InMux I__3406 (
            .O(N__22560),
            .I(N__22556));
    InMux I__3405 (
            .O(N__22559),
            .I(N__22553));
    LocalMux I__3404 (
            .O(N__22556),
            .I(N__22550));
    LocalMux I__3403 (
            .O(N__22553),
            .I(\c0.rx.r_Clock_Count_0 ));
    Odrv4 I__3402 (
            .O(N__22550),
            .I(\c0.rx.r_Clock_Count_0 ));
    CascadeMux I__3401 (
            .O(N__22545),
            .I(N__22542));
    InMux I__3400 (
            .O(N__22542),
            .I(N__22538));
    InMux I__3399 (
            .O(N__22541),
            .I(N__22535));
    LocalMux I__3398 (
            .O(N__22538),
            .I(N__22532));
    LocalMux I__3397 (
            .O(N__22535),
            .I(\c0.rx.r_Clock_Count_3 ));
    Odrv4 I__3396 (
            .O(N__22532),
            .I(\c0.rx.r_Clock_Count_3 ));
    InMux I__3395 (
            .O(N__22527),
            .I(N__22524));
    LocalMux I__3394 (
            .O(N__22524),
            .I(\c0.rx.n6 ));
    CascadeMux I__3393 (
            .O(N__22521),
            .I(\c0.rx.n17022_cascade_ ));
    CascadeMux I__3392 (
            .O(N__22518),
            .I(\c0.rx.r_SM_Main_2_N_2094_0_cascade_ ));
    CascadeMux I__3391 (
            .O(N__22515),
            .I(\c0.rx.n17380_cascade_ ));
    InMux I__3390 (
            .O(N__22512),
            .I(N__22509));
    LocalMux I__3389 (
            .O(N__22509),
            .I(\c0.rx.n17635 ));
    InMux I__3388 (
            .O(N__22506),
            .I(N__22503));
    LocalMux I__3387 (
            .O(N__22503),
            .I(N__22500));
    Odrv4 I__3386 (
            .O(N__22500),
            .I(\c0.n40 ));
    InMux I__3385 (
            .O(N__22497),
            .I(N__22494));
    LocalMux I__3384 (
            .O(N__22494),
            .I(N__22491));
    Span4Mux_h I__3383 (
            .O(N__22491),
            .I(N__22488));
    Odrv4 I__3382 (
            .O(N__22488),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_24 ));
    SRMux I__3381 (
            .O(N__22485),
            .I(N__22482));
    LocalMux I__3380 (
            .O(N__22482),
            .I(N__22479));
    Odrv4 I__3379 (
            .O(N__22479),
            .I(\c0.n3_adj_2242 ));
    SRMux I__3378 (
            .O(N__22476),
            .I(N__22473));
    LocalMux I__3377 (
            .O(N__22473),
            .I(N__22470));
    Span4Mux_v I__3376 (
            .O(N__22470),
            .I(N__22467));
    Odrv4 I__3375 (
            .O(N__22467),
            .I(\c0.n3_adj_2240 ));
    SRMux I__3374 (
            .O(N__22464),
            .I(N__22461));
    LocalMux I__3373 (
            .O(N__22461),
            .I(N__22458));
    Span4Mux_h I__3372 (
            .O(N__22458),
            .I(N__22455));
    Odrv4 I__3371 (
            .O(N__22455),
            .I(\c0.n3_adj_2234 ));
    SRMux I__3370 (
            .O(N__22452),
            .I(N__22449));
    LocalMux I__3369 (
            .O(N__22449),
            .I(N__22446));
    Span4Mux_h I__3368 (
            .O(N__22446),
            .I(N__22443));
    Odrv4 I__3367 (
            .O(N__22443),
            .I(\c0.n3_adj_2230 ));
    CascadeMux I__3366 (
            .O(N__22440),
            .I(\c0.n10009_cascade_ ));
    SRMux I__3365 (
            .O(N__22437),
            .I(N__22434));
    LocalMux I__3364 (
            .O(N__22434),
            .I(N__22431));
    Span4Mux_v I__3363 (
            .O(N__22431),
            .I(N__22428));
    Odrv4 I__3362 (
            .O(N__22428),
            .I(\c0.n3_adj_2181 ));
    InMux I__3361 (
            .O(N__22425),
            .I(N__22422));
    LocalMux I__3360 (
            .O(N__22422),
            .I(N__22419));
    Odrv4 I__3359 (
            .O(N__22419),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_18 ));
    InMux I__3358 (
            .O(N__22416),
            .I(N__22413));
    LocalMux I__3357 (
            .O(N__22413),
            .I(N__22410));
    Odrv4 I__3356 (
            .O(N__22410),
            .I(\c0.n42 ));
    CascadeMux I__3355 (
            .O(N__22407),
            .I(\c0.n41_adj_2376_cascade_ ));
    InMux I__3354 (
            .O(N__22404),
            .I(N__22401));
    LocalMux I__3353 (
            .O(N__22401),
            .I(\c0.n39_adj_2377 ));
    InMux I__3352 (
            .O(N__22398),
            .I(N__22395));
    LocalMux I__3351 (
            .O(N__22395),
            .I(N__22392));
    Span4Mux_h I__3350 (
            .O(N__22392),
            .I(N__22389));
    Odrv4 I__3349 (
            .O(N__22389),
            .I(\c0.n43_adj_2380 ));
    CascadeMux I__3348 (
            .O(N__22386),
            .I(\c0.n48_adj_2379_cascade_ ));
    InMux I__3347 (
            .O(N__22383),
            .I(N__22380));
    LocalMux I__3346 (
            .O(N__22380),
            .I(\c0.n44_adj_2378 ));
    CascadeMux I__3345 (
            .O(N__22377),
            .I(\c0.n9995_cascade_ ));
    InMux I__3344 (
            .O(N__22374),
            .I(N__22370));
    InMux I__3343 (
            .O(N__22373),
            .I(N__22367));
    LocalMux I__3342 (
            .O(N__22370),
            .I(\c0.n9995 ));
    LocalMux I__3341 (
            .O(N__22367),
            .I(\c0.n9995 ));
    InMux I__3340 (
            .O(N__22362),
            .I(N__22359));
    LocalMux I__3339 (
            .O(N__22359),
            .I(N__22356));
    Odrv4 I__3338 (
            .O(N__22356),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_2 ));
    SRMux I__3337 (
            .O(N__22353),
            .I(N__22350));
    LocalMux I__3336 (
            .O(N__22350),
            .I(N__22347));
    Odrv4 I__3335 (
            .O(N__22347),
            .I(\c0.n3_adj_2286 ));
    SRMux I__3334 (
            .O(N__22344),
            .I(N__22341));
    LocalMux I__3333 (
            .O(N__22341),
            .I(N__22338));
    Span4Mux_v I__3332 (
            .O(N__22338),
            .I(N__22335));
    Odrv4 I__3331 (
            .O(N__22335),
            .I(\c0.n3_adj_2226 ));
    InMux I__3330 (
            .O(N__22332),
            .I(N__22329));
    LocalMux I__3329 (
            .O(N__22329),
            .I(N__22326));
    Odrv4 I__3328 (
            .O(N__22326),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_2 ));
    InMux I__3327 (
            .O(N__22323),
            .I(N__22319));
    InMux I__3326 (
            .O(N__22322),
            .I(N__22316));
    LocalMux I__3325 (
            .O(N__22319),
            .I(N__22313));
    LocalMux I__3324 (
            .O(N__22316),
            .I(\c0.tx2.r_Clock_Count_3 ));
    Odrv4 I__3323 (
            .O(N__22313),
            .I(\c0.tx2.r_Clock_Count_3 ));
    InMux I__3322 (
            .O(N__22308),
            .I(\c0.tx2.n16134 ));
    CascadeMux I__3321 (
            .O(N__22305),
            .I(N__22301));
    InMux I__3320 (
            .O(N__22304),
            .I(N__22298));
    InMux I__3319 (
            .O(N__22301),
            .I(N__22295));
    LocalMux I__3318 (
            .O(N__22298),
            .I(\c0.tx2.r_Clock_Count_4 ));
    LocalMux I__3317 (
            .O(N__22295),
            .I(\c0.tx2.r_Clock_Count_4 ));
    InMux I__3316 (
            .O(N__22290),
            .I(\c0.tx2.n16135 ));
    CascadeMux I__3315 (
            .O(N__22287),
            .I(N__22284));
    InMux I__3314 (
            .O(N__22284),
            .I(N__22277));
    InMux I__3313 (
            .O(N__22283),
            .I(N__22277));
    InMux I__3312 (
            .O(N__22282),
            .I(N__22274));
    LocalMux I__3311 (
            .O(N__22277),
            .I(N__22271));
    LocalMux I__3310 (
            .O(N__22274),
            .I(\c0.tx2.r_Clock_Count_5 ));
    Odrv4 I__3309 (
            .O(N__22271),
            .I(\c0.tx2.r_Clock_Count_5 ));
    InMux I__3308 (
            .O(N__22266),
            .I(\c0.tx2.n16136 ));
    InMux I__3307 (
            .O(N__22263),
            .I(N__22259));
    InMux I__3306 (
            .O(N__22262),
            .I(N__22256));
    LocalMux I__3305 (
            .O(N__22259),
            .I(\c0.tx2.r_Clock_Count_6 ));
    LocalMux I__3304 (
            .O(N__22256),
            .I(\c0.tx2.r_Clock_Count_6 ));
    InMux I__3303 (
            .O(N__22251),
            .I(\c0.tx2.n16137 ));
    InMux I__3302 (
            .O(N__22248),
            .I(N__22244));
    InMux I__3301 (
            .O(N__22247),
            .I(N__22241));
    LocalMux I__3300 (
            .O(N__22244),
            .I(\c0.tx2.r_Clock_Count_7 ));
    LocalMux I__3299 (
            .O(N__22241),
            .I(\c0.tx2.r_Clock_Count_7 ));
    InMux I__3298 (
            .O(N__22236),
            .I(\c0.tx2.n16138 ));
    InMux I__3297 (
            .O(N__22233),
            .I(bfn_6_25_0_));
    InMux I__3296 (
            .O(N__22230),
            .I(N__22226));
    InMux I__3295 (
            .O(N__22229),
            .I(N__22223));
    LocalMux I__3294 (
            .O(N__22226),
            .I(N__22220));
    LocalMux I__3293 (
            .O(N__22223),
            .I(\c0.tx2.r_Clock_Count_8 ));
    Odrv4 I__3292 (
            .O(N__22220),
            .I(\c0.tx2.r_Clock_Count_8 ));
    SRMux I__3291 (
            .O(N__22215),
            .I(N__22211));
    SRMux I__3290 (
            .O(N__22214),
            .I(N__22208));
    LocalMux I__3289 (
            .O(N__22211),
            .I(N__22205));
    LocalMux I__3288 (
            .O(N__22208),
            .I(N__22202));
    Span4Mux_h I__3287 (
            .O(N__22205),
            .I(N__22199));
    Odrv4 I__3286 (
            .O(N__22202),
            .I(\c0.tx2.n10852 ));
    Odrv4 I__3285 (
            .O(N__22199),
            .I(\c0.tx2.n10852 ));
    InMux I__3284 (
            .O(N__22194),
            .I(N__22189));
    InMux I__3283 (
            .O(N__22193),
            .I(N__22186));
    CascadeMux I__3282 (
            .O(N__22192),
            .I(N__22183));
    LocalMux I__3281 (
            .O(N__22189),
            .I(N__22177));
    LocalMux I__3280 (
            .O(N__22186),
            .I(N__22177));
    InMux I__3279 (
            .O(N__22183),
            .I(N__22174));
    InMux I__3278 (
            .O(N__22182),
            .I(N__22171));
    Span4Mux_v I__3277 (
            .O(N__22177),
            .I(N__22166));
    LocalMux I__3276 (
            .O(N__22174),
            .I(N__22166));
    LocalMux I__3275 (
            .O(N__22171),
            .I(N__22163));
    Span4Mux_h I__3274 (
            .O(N__22166),
            .I(N__22160));
    Span4Mux_v I__3273 (
            .O(N__22163),
            .I(N__22157));
    Span4Mux_s0_h I__3272 (
            .O(N__22160),
            .I(N__22154));
    Span4Mux_h I__3271 (
            .O(N__22157),
            .I(N__22151));
    Odrv4 I__3270 (
            .O(N__22154),
            .I(\c0.FRAME_MATCHER_i_8 ));
    Odrv4 I__3269 (
            .O(N__22151),
            .I(\c0.FRAME_MATCHER_i_8 ));
    CascadeMux I__3268 (
            .O(N__22146),
            .I(N__22142));
    InMux I__3267 (
            .O(N__22145),
            .I(N__22139));
    InMux I__3266 (
            .O(N__22142),
            .I(N__22136));
    LocalMux I__3265 (
            .O(N__22139),
            .I(\c0.tx2.n10 ));
    LocalMux I__3264 (
            .O(N__22136),
            .I(\c0.tx2.n10 ));
    IoInMux I__3263 (
            .O(N__22131),
            .I(N__22128));
    LocalMux I__3262 (
            .O(N__22128),
            .I(N__22125));
    IoSpan4Mux I__3261 (
            .O(N__22125),
            .I(N__22122));
    Span4Mux_s2_h I__3260 (
            .O(N__22122),
            .I(N__22118));
    InMux I__3259 (
            .O(N__22121),
            .I(N__22115));
    Span4Mux_v I__3258 (
            .O(N__22118),
            .I(N__22109));
    LocalMux I__3257 (
            .O(N__22115),
            .I(N__22109));
    InMux I__3256 (
            .O(N__22114),
            .I(N__22106));
    Span4Mux_v I__3255 (
            .O(N__22109),
            .I(N__22103));
    LocalMux I__3254 (
            .O(N__22106),
            .I(N__22100));
    Odrv4 I__3253 (
            .O(N__22103),
            .I(tx2_o));
    Odrv4 I__3252 (
            .O(N__22100),
            .I(tx2_o));
    InMux I__3251 (
            .O(N__22095),
            .I(N__22090));
    InMux I__3250 (
            .O(N__22094),
            .I(N__22087));
    InMux I__3249 (
            .O(N__22093),
            .I(N__22084));
    LocalMux I__3248 (
            .O(N__22090),
            .I(N__22081));
    LocalMux I__3247 (
            .O(N__22087),
            .I(data_out_frame2_14_7));
    LocalMux I__3246 (
            .O(N__22084),
            .I(data_out_frame2_14_7));
    Odrv4 I__3245 (
            .O(N__22081),
            .I(data_out_frame2_14_7));
    InMux I__3244 (
            .O(N__22074),
            .I(N__22071));
    LocalMux I__3243 (
            .O(N__22071),
            .I(\c0.tx2.n17322 ));
    InMux I__3242 (
            .O(N__22068),
            .I(N__22062));
    InMux I__3241 (
            .O(N__22067),
            .I(N__22062));
    LocalMux I__3240 (
            .O(N__22062),
            .I(\c0.tx2.n17018 ));
    InMux I__3239 (
            .O(N__22059),
            .I(N__22055));
    InMux I__3238 (
            .O(N__22058),
            .I(N__22052));
    LocalMux I__3237 (
            .O(N__22055),
            .I(\c0.tx2.r_Clock_Count_0 ));
    LocalMux I__3236 (
            .O(N__22052),
            .I(\c0.tx2.r_Clock_Count_0 ));
    InMux I__3235 (
            .O(N__22047),
            .I(bfn_6_24_0_));
    InMux I__3234 (
            .O(N__22044),
            .I(N__22037));
    InMux I__3233 (
            .O(N__22043),
            .I(N__22037));
    InMux I__3232 (
            .O(N__22042),
            .I(N__22034));
    LocalMux I__3231 (
            .O(N__22037),
            .I(N__22031));
    LocalMux I__3230 (
            .O(N__22034),
            .I(\c0.tx2.r_Clock_Count_1 ));
    Odrv4 I__3229 (
            .O(N__22031),
            .I(\c0.tx2.r_Clock_Count_1 ));
    InMux I__3228 (
            .O(N__22026),
            .I(\c0.tx2.n16132 ));
    InMux I__3227 (
            .O(N__22023),
            .I(N__22019));
    InMux I__3226 (
            .O(N__22022),
            .I(N__22016));
    LocalMux I__3225 (
            .O(N__22019),
            .I(\c0.tx2.r_Clock_Count_2 ));
    LocalMux I__3224 (
            .O(N__22016),
            .I(\c0.tx2.r_Clock_Count_2 ));
    InMux I__3223 (
            .O(N__22011),
            .I(\c0.tx2.n16133 ));
    CascadeMux I__3222 (
            .O(N__22008),
            .I(\c0.tx2.n13748_cascade_ ));
    InMux I__3221 (
            .O(N__22005),
            .I(N__22002));
    LocalMux I__3220 (
            .O(N__22002),
            .I(N__21998));
    InMux I__3219 (
            .O(N__22001),
            .I(N__21995));
    Span4Mux_h I__3218 (
            .O(N__21998),
            .I(N__21992));
    LocalMux I__3217 (
            .O(N__21995),
            .I(N__21987));
    Span4Mux_v I__3216 (
            .O(N__21992),
            .I(N__21987));
    Odrv4 I__3215 (
            .O(N__21987),
            .I(data_out_frame2_18_7));
    CascadeMux I__3214 (
            .O(N__21984),
            .I(N__21981));
    InMux I__3213 (
            .O(N__21981),
            .I(N__21978));
    LocalMux I__3212 (
            .O(N__21978),
            .I(N__21974));
    InMux I__3211 (
            .O(N__21977),
            .I(N__21971));
    Span4Mux_h I__3210 (
            .O(N__21974),
            .I(N__21968));
    LocalMux I__3209 (
            .O(N__21971),
            .I(data_out_frame2_17_2));
    Odrv4 I__3208 (
            .O(N__21968),
            .I(data_out_frame2_17_2));
    InMux I__3207 (
            .O(N__21963),
            .I(N__21959));
    InMux I__3206 (
            .O(N__21962),
            .I(N__21952));
    LocalMux I__3205 (
            .O(N__21959),
            .I(N__21949));
    InMux I__3204 (
            .O(N__21958),
            .I(N__21946));
    InMux I__3203 (
            .O(N__21957),
            .I(N__21943));
    InMux I__3202 (
            .O(N__21956),
            .I(N__21940));
    InMux I__3201 (
            .O(N__21955),
            .I(N__21937));
    LocalMux I__3200 (
            .O(N__21952),
            .I(N__21934));
    Span4Mux_v I__3199 (
            .O(N__21949),
            .I(N__21931));
    LocalMux I__3198 (
            .O(N__21946),
            .I(N__21928));
    LocalMux I__3197 (
            .O(N__21943),
            .I(N__21925));
    LocalMux I__3196 (
            .O(N__21940),
            .I(N__21922));
    LocalMux I__3195 (
            .O(N__21937),
            .I(N__21919));
    Span4Mux_v I__3194 (
            .O(N__21934),
            .I(N__21914));
    Span4Mux_v I__3193 (
            .O(N__21931),
            .I(N__21914));
    Span12Mux_v I__3192 (
            .O(N__21928),
            .I(N__21911));
    Span4Mux_h I__3191 (
            .O(N__21925),
            .I(N__21906));
    Span4Mux_h I__3190 (
            .O(N__21922),
            .I(N__21906));
    Odrv4 I__3189 (
            .O(N__21919),
            .I(data_out_frame2_7_5));
    Odrv4 I__3188 (
            .O(N__21914),
            .I(data_out_frame2_7_5));
    Odrv12 I__3187 (
            .O(N__21911),
            .I(data_out_frame2_7_5));
    Odrv4 I__3186 (
            .O(N__21906),
            .I(data_out_frame2_7_5));
    InMux I__3185 (
            .O(N__21897),
            .I(N__21890));
    InMux I__3184 (
            .O(N__21896),
            .I(N__21887));
    InMux I__3183 (
            .O(N__21895),
            .I(N__21882));
    InMux I__3182 (
            .O(N__21894),
            .I(N__21882));
    InMux I__3181 (
            .O(N__21893),
            .I(N__21879));
    LocalMux I__3180 (
            .O(N__21890),
            .I(data_out_frame2_11_4));
    LocalMux I__3179 (
            .O(N__21887),
            .I(data_out_frame2_11_4));
    LocalMux I__3178 (
            .O(N__21882),
            .I(data_out_frame2_11_4));
    LocalMux I__3177 (
            .O(N__21879),
            .I(data_out_frame2_11_4));
    InMux I__3176 (
            .O(N__21870),
            .I(N__21861));
    InMux I__3175 (
            .O(N__21869),
            .I(N__21861));
    InMux I__3174 (
            .O(N__21868),
            .I(N__21857));
    CascadeMux I__3173 (
            .O(N__21867),
            .I(N__21854));
    InMux I__3172 (
            .O(N__21866),
            .I(N__21851));
    LocalMux I__3171 (
            .O(N__21861),
            .I(N__21848));
    InMux I__3170 (
            .O(N__21860),
            .I(N__21845));
    LocalMux I__3169 (
            .O(N__21857),
            .I(N__21842));
    InMux I__3168 (
            .O(N__21854),
            .I(N__21839));
    LocalMux I__3167 (
            .O(N__21851),
            .I(data_out_frame2_11_5));
    Odrv12 I__3166 (
            .O(N__21848),
            .I(data_out_frame2_11_5));
    LocalMux I__3165 (
            .O(N__21845),
            .I(data_out_frame2_11_5));
    Odrv4 I__3164 (
            .O(N__21842),
            .I(data_out_frame2_11_5));
    LocalMux I__3163 (
            .O(N__21839),
            .I(data_out_frame2_11_5));
    InMux I__3162 (
            .O(N__21828),
            .I(N__21825));
    LocalMux I__3161 (
            .O(N__21825),
            .I(N__21821));
    InMux I__3160 (
            .O(N__21824),
            .I(N__21817));
    Span4Mux_s1_h I__3159 (
            .O(N__21821),
            .I(N__21814));
    InMux I__3158 (
            .O(N__21820),
            .I(N__21811));
    LocalMux I__3157 (
            .O(N__21817),
            .I(N__21808));
    Span4Mux_h I__3156 (
            .O(N__21814),
            .I(N__21805));
    LocalMux I__3155 (
            .O(N__21811),
            .I(N__21800));
    Span4Mux_v I__3154 (
            .O(N__21808),
            .I(N__21800));
    Odrv4 I__3153 (
            .O(N__21805),
            .I(\c0.n10359 ));
    Odrv4 I__3152 (
            .O(N__21800),
            .I(\c0.n10359 ));
    InMux I__3151 (
            .O(N__21795),
            .I(N__21791));
    InMux I__3150 (
            .O(N__21794),
            .I(N__21788));
    LocalMux I__3149 (
            .O(N__21791),
            .I(N__21784));
    LocalMux I__3148 (
            .O(N__21788),
            .I(N__21780));
    CascadeMux I__3147 (
            .O(N__21787),
            .I(N__21777));
    Span4Mux_s2_h I__3146 (
            .O(N__21784),
            .I(N__21774));
    InMux I__3145 (
            .O(N__21783),
            .I(N__21771));
    Span4Mux_h I__3144 (
            .O(N__21780),
            .I(N__21768));
    InMux I__3143 (
            .O(N__21777),
            .I(N__21765));
    Span4Mux_h I__3142 (
            .O(N__21774),
            .I(N__21762));
    LocalMux I__3141 (
            .O(N__21771),
            .I(data_out_frame2_5_4));
    Odrv4 I__3140 (
            .O(N__21768),
            .I(data_out_frame2_5_4));
    LocalMux I__3139 (
            .O(N__21765),
            .I(data_out_frame2_5_4));
    Odrv4 I__3138 (
            .O(N__21762),
            .I(data_out_frame2_5_4));
    InMux I__3137 (
            .O(N__21753),
            .I(N__21749));
    InMux I__3136 (
            .O(N__21752),
            .I(N__21746));
    LocalMux I__3135 (
            .O(N__21749),
            .I(N__21742));
    LocalMux I__3134 (
            .O(N__21746),
            .I(N__21737));
    InMux I__3133 (
            .O(N__21745),
            .I(N__21734));
    Span4Mux_h I__3132 (
            .O(N__21742),
            .I(N__21731));
    InMux I__3131 (
            .O(N__21741),
            .I(N__21726));
    InMux I__3130 (
            .O(N__21740),
            .I(N__21726));
    Odrv4 I__3129 (
            .O(N__21737),
            .I(data_out_frame2_10_7));
    LocalMux I__3128 (
            .O(N__21734),
            .I(data_out_frame2_10_7));
    Odrv4 I__3127 (
            .O(N__21731),
            .I(data_out_frame2_10_7));
    LocalMux I__3126 (
            .O(N__21726),
            .I(data_out_frame2_10_7));
    CascadeMux I__3125 (
            .O(N__21717),
            .I(N__21714));
    InMux I__3124 (
            .O(N__21714),
            .I(N__21710));
    InMux I__3123 (
            .O(N__21713),
            .I(N__21707));
    LocalMux I__3122 (
            .O(N__21710),
            .I(N__21704));
    LocalMux I__3121 (
            .O(N__21707),
            .I(data_out_frame2_17_0));
    Odrv4 I__3120 (
            .O(N__21704),
            .I(data_out_frame2_17_0));
    CascadeMux I__3119 (
            .O(N__21699),
            .I(N__21696));
    InMux I__3118 (
            .O(N__21696),
            .I(N__21693));
    LocalMux I__3117 (
            .O(N__21693),
            .I(N__21690));
    Odrv12 I__3116 (
            .O(N__21690),
            .I(\c0.n18163 ));
    InMux I__3115 (
            .O(N__21687),
            .I(N__21684));
    LocalMux I__3114 (
            .O(N__21684),
            .I(\c0.n18208 ));
    InMux I__3113 (
            .O(N__21681),
            .I(N__21677));
    InMux I__3112 (
            .O(N__21680),
            .I(N__21674));
    LocalMux I__3111 (
            .O(N__21677),
            .I(N__21671));
    LocalMux I__3110 (
            .O(N__21674),
            .I(data_out_frame2_17_3));
    Odrv4 I__3109 (
            .O(N__21671),
            .I(data_out_frame2_17_3));
    InMux I__3108 (
            .O(N__21666),
            .I(N__21661));
    InMux I__3107 (
            .O(N__21665),
            .I(N__21657));
    InMux I__3106 (
            .O(N__21664),
            .I(N__21654));
    LocalMux I__3105 (
            .O(N__21661),
            .I(N__21651));
    InMux I__3104 (
            .O(N__21660),
            .I(N__21648));
    LocalMux I__3103 (
            .O(N__21657),
            .I(N__21645));
    LocalMux I__3102 (
            .O(N__21654),
            .I(N__21642));
    Span4Mux_h I__3101 (
            .O(N__21651),
            .I(N__21639));
    LocalMux I__3100 (
            .O(N__21648),
            .I(data_out_frame2_14_2));
    Odrv12 I__3099 (
            .O(N__21645),
            .I(data_out_frame2_14_2));
    Odrv4 I__3098 (
            .O(N__21642),
            .I(data_out_frame2_14_2));
    Odrv4 I__3097 (
            .O(N__21639),
            .I(data_out_frame2_14_2));
    InMux I__3096 (
            .O(N__21630),
            .I(N__21627));
    LocalMux I__3095 (
            .O(N__21627),
            .I(N__21624));
    Span4Mux_h I__3094 (
            .O(N__21624),
            .I(N__21621));
    Span4Mux_h I__3093 (
            .O(N__21621),
            .I(N__21618));
    Odrv4 I__3092 (
            .O(N__21618),
            .I(\c0.n10_adj_2207 ));
    CascadeMux I__3091 (
            .O(N__21615),
            .I(N__21612));
    InMux I__3090 (
            .O(N__21612),
            .I(N__21609));
    LocalMux I__3089 (
            .O(N__21609),
            .I(N__21606));
    Span4Mux_h I__3088 (
            .O(N__21606),
            .I(N__21603));
    Odrv4 I__3087 (
            .O(N__21603),
            .I(\c0.n18061 ));
    CascadeMux I__3086 (
            .O(N__21600),
            .I(\c0.n18256_cascade_ ));
    InMux I__3085 (
            .O(N__21597),
            .I(N__21594));
    LocalMux I__3084 (
            .O(N__21594),
            .I(\c0.n6_adj_2139 ));
    InMux I__3083 (
            .O(N__21591),
            .I(N__21588));
    LocalMux I__3082 (
            .O(N__21588),
            .I(\c0.n22_adj_2371 ));
    CascadeMux I__3081 (
            .O(N__21585),
            .I(\c0.n18259_cascade_ ));
    InMux I__3080 (
            .O(N__21582),
            .I(N__21579));
    LocalMux I__3079 (
            .O(N__21579),
            .I(N__21576));
    Odrv4 I__3078 (
            .O(N__21576),
            .I(\c0.tx2.r_Tx_Data_3 ));
    InMux I__3077 (
            .O(N__21573),
            .I(N__21568));
    InMux I__3076 (
            .O(N__21572),
            .I(N__21565));
    InMux I__3075 (
            .O(N__21571),
            .I(N__21561));
    LocalMux I__3074 (
            .O(N__21568),
            .I(N__21558));
    LocalMux I__3073 (
            .O(N__21565),
            .I(N__21555));
    InMux I__3072 (
            .O(N__21564),
            .I(N__21552));
    LocalMux I__3071 (
            .O(N__21561),
            .I(N__21547));
    Span4Mux_v I__3070 (
            .O(N__21558),
            .I(N__21547));
    Span4Mux_h I__3069 (
            .O(N__21555),
            .I(N__21544));
    LocalMux I__3068 (
            .O(N__21552),
            .I(data_out_frame2_10_1));
    Odrv4 I__3067 (
            .O(N__21547),
            .I(data_out_frame2_10_1));
    Odrv4 I__3066 (
            .O(N__21544),
            .I(data_out_frame2_10_1));
    InMux I__3065 (
            .O(N__21537),
            .I(N__21534));
    LocalMux I__3064 (
            .O(N__21534),
            .I(N__21531));
    Span4Mux_h I__3063 (
            .O(N__21531),
            .I(N__21528));
    Odrv4 I__3062 (
            .O(N__21528),
            .I(\c0.n17203 ));
    InMux I__3061 (
            .O(N__21525),
            .I(N__21519));
    InMux I__3060 (
            .O(N__21524),
            .I(N__21516));
    InMux I__3059 (
            .O(N__21523),
            .I(N__21513));
    InMux I__3058 (
            .O(N__21522),
            .I(N__21510));
    LocalMux I__3057 (
            .O(N__21519),
            .I(N__21506));
    LocalMux I__3056 (
            .O(N__21516),
            .I(N__21503));
    LocalMux I__3055 (
            .O(N__21513),
            .I(N__21500));
    LocalMux I__3054 (
            .O(N__21510),
            .I(N__21497));
    InMux I__3053 (
            .O(N__21509),
            .I(N__21494));
    Span4Mux_h I__3052 (
            .O(N__21506),
            .I(N__21491));
    Span4Mux_v I__3051 (
            .O(N__21503),
            .I(N__21486));
    Span4Mux_h I__3050 (
            .O(N__21500),
            .I(N__21486));
    Span4Mux_h I__3049 (
            .O(N__21497),
            .I(N__21483));
    LocalMux I__3048 (
            .O(N__21494),
            .I(data_out_frame2_8_6));
    Odrv4 I__3047 (
            .O(N__21491),
            .I(data_out_frame2_8_6));
    Odrv4 I__3046 (
            .O(N__21486),
            .I(data_out_frame2_8_6));
    Odrv4 I__3045 (
            .O(N__21483),
            .I(data_out_frame2_8_6));
    CascadeMux I__3044 (
            .O(N__21474),
            .I(N__21471));
    InMux I__3043 (
            .O(N__21471),
            .I(N__21468));
    LocalMux I__3042 (
            .O(N__21468),
            .I(N__21464));
    InMux I__3041 (
            .O(N__21467),
            .I(N__21461));
    Span4Mux_v I__3040 (
            .O(N__21464),
            .I(N__21458));
    LocalMux I__3039 (
            .O(N__21461),
            .I(N__21453));
    Span4Mux_v I__3038 (
            .O(N__21458),
            .I(N__21450));
    InMux I__3037 (
            .O(N__21457),
            .I(N__21447));
    InMux I__3036 (
            .O(N__21456),
            .I(N__21444));
    Span4Mux_s3_h I__3035 (
            .O(N__21453),
            .I(N__21441));
    Span4Mux_h I__3034 (
            .O(N__21450),
            .I(N__21436));
    LocalMux I__3033 (
            .O(N__21447),
            .I(N__21436));
    LocalMux I__3032 (
            .O(N__21444),
            .I(data_out_frame2_9_6));
    Odrv4 I__3031 (
            .O(N__21441),
            .I(data_out_frame2_9_6));
    Odrv4 I__3030 (
            .O(N__21436),
            .I(data_out_frame2_9_6));
    InMux I__3029 (
            .O(N__21429),
            .I(N__21426));
    LocalMux I__3028 (
            .O(N__21426),
            .I(N__21423));
    Span4Mux_v I__3027 (
            .O(N__21423),
            .I(N__21420));
    Odrv4 I__3026 (
            .O(N__21420),
            .I(\c0.n18127 ));
    InMux I__3025 (
            .O(N__21417),
            .I(N__21413));
    InMux I__3024 (
            .O(N__21416),
            .I(N__21410));
    LocalMux I__3023 (
            .O(N__21413),
            .I(data_out_frame2_18_3));
    LocalMux I__3022 (
            .O(N__21410),
            .I(data_out_frame2_18_3));
    InMux I__3021 (
            .O(N__21405),
            .I(N__21402));
    LocalMux I__3020 (
            .O(N__21402),
            .I(\c0.n22_adj_2387 ));
    InMux I__3019 (
            .O(N__21399),
            .I(N__21396));
    LocalMux I__3018 (
            .O(N__21396),
            .I(\c0.tx2.r_Tx_Data_0 ));
    InMux I__3017 (
            .O(N__21393),
            .I(N__21390));
    LocalMux I__3016 (
            .O(N__21390),
            .I(N__21387));
    Odrv12 I__3015 (
            .O(N__21387),
            .I(\c0.n18157 ));
    InMux I__3014 (
            .O(N__21384),
            .I(N__21381));
    LocalMux I__3013 (
            .O(N__21381),
            .I(\c0.n17603 ));
    CascadeMux I__3012 (
            .O(N__21378),
            .I(\c0.n18226_cascade_ ));
    InMux I__3011 (
            .O(N__21375),
            .I(N__21372));
    LocalMux I__3010 (
            .O(N__21372),
            .I(\c0.n18229 ));
    CascadeMux I__3009 (
            .O(N__21369),
            .I(N__21365));
    InMux I__3008 (
            .O(N__21368),
            .I(N__21361));
    InMux I__3007 (
            .O(N__21365),
            .I(N__21354));
    InMux I__3006 (
            .O(N__21364),
            .I(N__21354));
    LocalMux I__3005 (
            .O(N__21361),
            .I(N__21350));
    InMux I__3004 (
            .O(N__21360),
            .I(N__21347));
    InMux I__3003 (
            .O(N__21359),
            .I(N__21344));
    LocalMux I__3002 (
            .O(N__21354),
            .I(N__21341));
    InMux I__3001 (
            .O(N__21353),
            .I(N__21338));
    Span4Mux_v I__3000 (
            .O(N__21350),
            .I(N__21335));
    LocalMux I__2999 (
            .O(N__21347),
            .I(data_out_frame2_10_0));
    LocalMux I__2998 (
            .O(N__21344),
            .I(data_out_frame2_10_0));
    Odrv4 I__2997 (
            .O(N__21341),
            .I(data_out_frame2_10_0));
    LocalMux I__2996 (
            .O(N__21338),
            .I(data_out_frame2_10_0));
    Odrv4 I__2995 (
            .O(N__21335),
            .I(data_out_frame2_10_0));
    CascadeMux I__2994 (
            .O(N__21324),
            .I(\c0.n18148_cascade_ ));
    CascadeMux I__2993 (
            .O(N__21321),
            .I(N__21318));
    InMux I__2992 (
            .O(N__21318),
            .I(N__21315));
    LocalMux I__2991 (
            .O(N__21315),
            .I(\c0.n18151 ));
    InMux I__2990 (
            .O(N__21312),
            .I(N__21308));
    InMux I__2989 (
            .O(N__21311),
            .I(N__21305));
    LocalMux I__2988 (
            .O(N__21308),
            .I(N__21301));
    LocalMux I__2987 (
            .O(N__21305),
            .I(N__21297));
    CascadeMux I__2986 (
            .O(N__21304),
            .I(N__21294));
    Span4Mux_h I__2985 (
            .O(N__21301),
            .I(N__21290));
    InMux I__2984 (
            .O(N__21300),
            .I(N__21287));
    Span4Mux_v I__2983 (
            .O(N__21297),
            .I(N__21284));
    InMux I__2982 (
            .O(N__21294),
            .I(N__21279));
    InMux I__2981 (
            .O(N__21293),
            .I(N__21279));
    Span4Mux_v I__2980 (
            .O(N__21290),
            .I(N__21274));
    LocalMux I__2979 (
            .O(N__21287),
            .I(N__21274));
    Odrv4 I__2978 (
            .O(N__21284),
            .I(data_out_frame2_5_0));
    LocalMux I__2977 (
            .O(N__21279),
            .I(data_out_frame2_5_0));
    Odrv4 I__2976 (
            .O(N__21274),
            .I(data_out_frame2_5_0));
    CascadeMux I__2975 (
            .O(N__21267),
            .I(N__21264));
    InMux I__2974 (
            .O(N__21264),
            .I(N__21261));
    LocalMux I__2973 (
            .O(N__21261),
            .I(N__21258));
    Span4Mux_h I__2972 (
            .O(N__21258),
            .I(N__21255));
    Span4Mux_v I__2971 (
            .O(N__21255),
            .I(N__21252));
    Span4Mux_h I__2970 (
            .O(N__21252),
            .I(N__21249));
    Odrv4 I__2969 (
            .O(N__21249),
            .I(\c0.n5_adj_2217 ));
    InMux I__2968 (
            .O(N__21246),
            .I(N__21243));
    LocalMux I__2967 (
            .O(N__21243),
            .I(\c0.n6_adj_2143 ));
    CascadeMux I__2966 (
            .O(N__21240),
            .I(N__21237));
    InMux I__2965 (
            .O(N__21237),
            .I(N__21234));
    LocalMux I__2964 (
            .O(N__21234),
            .I(N__21231));
    Odrv12 I__2963 (
            .O(N__21231),
            .I(\c0.data_out_frame2_19_3 ));
    CascadeMux I__2962 (
            .O(N__21228),
            .I(\c0.n18052_cascade_ ));
    InMux I__2961 (
            .O(N__21225),
            .I(N__21222));
    LocalMux I__2960 (
            .O(N__21222),
            .I(N__21219));
    Odrv12 I__2959 (
            .O(N__21219),
            .I(\c0.data_out_frame2_20_3 ));
    CascadeMux I__2958 (
            .O(N__21216),
            .I(\c0.n18055_cascade_ ));
    InMux I__2957 (
            .O(N__21213),
            .I(N__21207));
    InMux I__2956 (
            .O(N__21212),
            .I(N__21204));
    InMux I__2955 (
            .O(N__21211),
            .I(N__21200));
    InMux I__2954 (
            .O(N__21210),
            .I(N__21196));
    LocalMux I__2953 (
            .O(N__21207),
            .I(N__21191));
    LocalMux I__2952 (
            .O(N__21204),
            .I(N__21188));
    InMux I__2951 (
            .O(N__21203),
            .I(N__21185));
    LocalMux I__2950 (
            .O(N__21200),
            .I(N__21182));
    InMux I__2949 (
            .O(N__21199),
            .I(N__21179));
    LocalMux I__2948 (
            .O(N__21196),
            .I(N__21176));
    InMux I__2947 (
            .O(N__21195),
            .I(N__21173));
    InMux I__2946 (
            .O(N__21194),
            .I(N__21170));
    Span4Mux_v I__2945 (
            .O(N__21191),
            .I(N__21167));
    Span4Mux_s3_h I__2944 (
            .O(N__21188),
            .I(N__21162));
    LocalMux I__2943 (
            .O(N__21185),
            .I(N__21162));
    Span4Mux_v I__2942 (
            .O(N__21182),
            .I(N__21153));
    LocalMux I__2941 (
            .O(N__21179),
            .I(N__21153));
    Span4Mux_v I__2940 (
            .O(N__21176),
            .I(N__21153));
    LocalMux I__2939 (
            .O(N__21173),
            .I(N__21153));
    LocalMux I__2938 (
            .O(N__21170),
            .I(N__21150));
    Span4Mux_s3_h I__2937 (
            .O(N__21167),
            .I(N__21145));
    Span4Mux_v I__2936 (
            .O(N__21162),
            .I(N__21145));
    Span4Mux_h I__2935 (
            .O(N__21153),
            .I(N__21142));
    Odrv12 I__2934 (
            .O(N__21150),
            .I(\c0.n9157 ));
    Odrv4 I__2933 (
            .O(N__21145),
            .I(\c0.n9157 ));
    Odrv4 I__2932 (
            .O(N__21142),
            .I(\c0.n9157 ));
    CascadeMux I__2931 (
            .O(N__21135),
            .I(n17708_cascade_));
    InMux I__2930 (
            .O(N__21132),
            .I(N__21128));
    InMux I__2929 (
            .O(N__21131),
            .I(N__21125));
    LocalMux I__2928 (
            .O(N__21128),
            .I(n5244));
    LocalMux I__2927 (
            .O(N__21125),
            .I(n5244));
    InMux I__2926 (
            .O(N__21120),
            .I(N__21116));
    InMux I__2925 (
            .O(N__21119),
            .I(N__21113));
    LocalMux I__2924 (
            .O(N__21116),
            .I(n11018));
    LocalMux I__2923 (
            .O(N__21113),
            .I(n11018));
    InMux I__2922 (
            .O(N__21108),
            .I(N__21105));
    LocalMux I__2921 (
            .O(N__21105),
            .I(\c0.data_out_frame2_20_0 ));
    InMux I__2920 (
            .O(N__21102),
            .I(N__21099));
    LocalMux I__2919 (
            .O(N__21099),
            .I(N__21096));
    Span4Mux_h I__2918 (
            .O(N__21096),
            .I(N__21093));
    Span4Mux_v I__2917 (
            .O(N__21093),
            .I(N__21090));
    Odrv4 I__2916 (
            .O(N__21090),
            .I(\c0.n18049 ));
    CascadeMux I__2915 (
            .O(N__21087),
            .I(N__21084));
    InMux I__2914 (
            .O(N__21084),
            .I(N__21081));
    LocalMux I__2913 (
            .O(N__21081),
            .I(N__21078));
    Span4Mux_h I__2912 (
            .O(N__21078),
            .I(N__21075));
    Odrv4 I__2911 (
            .O(N__21075),
            .I(\c0.n18043 ));
    InMux I__2910 (
            .O(N__21072),
            .I(N__21069));
    LocalMux I__2909 (
            .O(N__21069),
            .I(N__21066));
    Span4Mux_h I__2908 (
            .O(N__21066),
            .I(N__21063));
    Odrv4 I__2907 (
            .O(N__21063),
            .I(\c0.n17586 ));
    CascadeMux I__2906 (
            .O(N__21060),
            .I(\c0.n18244_cascade_ ));
    InMux I__2905 (
            .O(N__21057),
            .I(N__21054));
    LocalMux I__2904 (
            .O(N__21054),
            .I(\c0.n6_adj_2140 ));
    InMux I__2903 (
            .O(N__21051),
            .I(N__21048));
    LocalMux I__2902 (
            .O(N__21048),
            .I(N__21045));
    Odrv12 I__2901 (
            .O(N__21045),
            .I(\c0.tx2.r_Tx_Data_1 ));
    CascadeMux I__2900 (
            .O(N__21042),
            .I(\c0.tx2.n18232_cascade_ ));
    CascadeMux I__2899 (
            .O(N__21039),
            .I(N__21036));
    InMux I__2898 (
            .O(N__21036),
            .I(N__21033));
    LocalMux I__2897 (
            .O(N__21033),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_31 ));
    InMux I__2896 (
            .O(N__21030),
            .I(N__21027));
    LocalMux I__2895 (
            .O(N__21027),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_25 ));
    InMux I__2894 (
            .O(N__21024),
            .I(N__21021));
    LocalMux I__2893 (
            .O(N__21021),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_26 ));
    SRMux I__2892 (
            .O(N__21018),
            .I(N__21015));
    LocalMux I__2891 (
            .O(N__21015),
            .I(N__21012));
    Odrv4 I__2890 (
            .O(N__21012),
            .I(\c0.rx.n10845 ));
    InMux I__2889 (
            .O(N__21009),
            .I(N__21006));
    LocalMux I__2888 (
            .O(N__21006),
            .I(n1));
    InMux I__2887 (
            .O(N__21003),
            .I(N__20999));
    InMux I__2886 (
            .O(N__21002),
            .I(N__20996));
    LocalMux I__2885 (
            .O(N__20999),
            .I(\c0.rx.r_Clock_Count_4 ));
    LocalMux I__2884 (
            .O(N__20996),
            .I(\c0.rx.r_Clock_Count_4 ));
    InMux I__2883 (
            .O(N__20991),
            .I(N__20987));
    InMux I__2882 (
            .O(N__20990),
            .I(N__20984));
    LocalMux I__2881 (
            .O(N__20987),
            .I(\c0.rx.r_Clock_Count_1 ));
    LocalMux I__2880 (
            .O(N__20984),
            .I(\c0.rx.r_Clock_Count_1 ));
    CEMux I__2879 (
            .O(N__20979),
            .I(N__20976));
    LocalMux I__2878 (
            .O(N__20976),
            .I(N__20973));
    Span4Mux_h I__2877 (
            .O(N__20973),
            .I(N__20970));
    Odrv4 I__2876 (
            .O(N__20970),
            .I(\c0.rx.n10656 ));
    SRMux I__2875 (
            .O(N__20967),
            .I(N__20964));
    LocalMux I__2874 (
            .O(N__20964),
            .I(N__20961));
    Span4Mux_s1_h I__2873 (
            .O(N__20961),
            .I(N__20958));
    Span4Mux_h I__2872 (
            .O(N__20958),
            .I(N__20955));
    Odrv4 I__2871 (
            .O(N__20955),
            .I(\c0.n3_adj_2244 ));
    CascadeMux I__2870 (
            .O(N__20952),
            .I(N__20949));
    InMux I__2869 (
            .O(N__20949),
            .I(N__20943));
    InMux I__2868 (
            .O(N__20948),
            .I(N__20936));
    InMux I__2867 (
            .O(N__20947),
            .I(N__20936));
    InMux I__2866 (
            .O(N__20946),
            .I(N__20936));
    LocalMux I__2865 (
            .O(N__20943),
            .I(N__20933));
    LocalMux I__2864 (
            .O(N__20936),
            .I(N__20930));
    Span4Mux_h I__2863 (
            .O(N__20933),
            .I(N__20927));
    Span12Mux_h I__2862 (
            .O(N__20930),
            .I(N__20924));
    Odrv4 I__2861 (
            .O(N__20927),
            .I(\c0.FRAME_MATCHER_i_21 ));
    Odrv12 I__2860 (
            .O(N__20924),
            .I(\c0.FRAME_MATCHER_i_21 ));
    InMux I__2859 (
            .O(N__20919),
            .I(N__20916));
    LocalMux I__2858 (
            .O(N__20916),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_21 ));
    InMux I__2857 (
            .O(N__20913),
            .I(N__20910));
    LocalMux I__2856 (
            .O(N__20910),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_27 ));
    SRMux I__2855 (
            .O(N__20907),
            .I(N__20904));
    LocalMux I__2854 (
            .O(N__20904),
            .I(N__20901));
    Span4Mux_v I__2853 (
            .O(N__20901),
            .I(N__20898));
    Span4Mux_h I__2852 (
            .O(N__20898),
            .I(N__20895));
    Odrv4 I__2851 (
            .O(N__20895),
            .I(\c0.n3_adj_2276 ));
    InMux I__2850 (
            .O(N__20892),
            .I(N__20889));
    LocalMux I__2849 (
            .O(N__20889),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_8 ));
    InMux I__2848 (
            .O(N__20886),
            .I(N__20883));
    LocalMux I__2847 (
            .O(N__20883),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_9 ));
    InMux I__2846 (
            .O(N__20880),
            .I(N__20874));
    InMux I__2845 (
            .O(N__20879),
            .I(N__20867));
    InMux I__2844 (
            .O(N__20878),
            .I(N__20867));
    InMux I__2843 (
            .O(N__20877),
            .I(N__20867));
    LocalMux I__2842 (
            .O(N__20874),
            .I(\c0.FRAME_MATCHER_i_6 ));
    LocalMux I__2841 (
            .O(N__20867),
            .I(\c0.FRAME_MATCHER_i_6 ));
    InMux I__2840 (
            .O(N__20862),
            .I(N__20859));
    LocalMux I__2839 (
            .O(N__20859),
            .I(\c0.n41 ));
    SRMux I__2838 (
            .O(N__20856),
            .I(N__20853));
    LocalMux I__2837 (
            .O(N__20853),
            .I(N__20850));
    Span4Mux_s1_h I__2836 (
            .O(N__20850),
            .I(N__20847));
    Span4Mux_h I__2835 (
            .O(N__20847),
            .I(N__20844));
    Odrv4 I__2834 (
            .O(N__20844),
            .I(\c0.n3_adj_2261 ));
    SRMux I__2833 (
            .O(N__20841),
            .I(N__20838));
    LocalMux I__2832 (
            .O(N__20838),
            .I(N__20835));
    Span4Mux_s1_h I__2831 (
            .O(N__20835),
            .I(N__20832));
    Span4Mux_h I__2830 (
            .O(N__20832),
            .I(N__20829));
    Odrv4 I__2829 (
            .O(N__20829),
            .I(\c0.n3_adj_2270 ));
    SRMux I__2828 (
            .O(N__20826),
            .I(N__20823));
    LocalMux I__2827 (
            .O(N__20823),
            .I(N__20820));
    Span4Mux_s2_h I__2826 (
            .O(N__20820),
            .I(N__20817));
    Odrv4 I__2825 (
            .O(N__20817),
            .I(\c0.n3_adj_2252 ));
    InMux I__2824 (
            .O(N__20814),
            .I(N__20811));
    LocalMux I__2823 (
            .O(N__20811),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_17 ));
    SRMux I__2822 (
            .O(N__20808),
            .I(N__20805));
    LocalMux I__2821 (
            .O(N__20805),
            .I(N__20802));
    Odrv4 I__2820 (
            .O(N__20802),
            .I(\c0.n3_adj_2257 ));
    InMux I__2819 (
            .O(N__20799),
            .I(N__20793));
    InMux I__2818 (
            .O(N__20798),
            .I(N__20786));
    InMux I__2817 (
            .O(N__20797),
            .I(N__20786));
    InMux I__2816 (
            .O(N__20796),
            .I(N__20786));
    LocalMux I__2815 (
            .O(N__20793),
            .I(\c0.FRAME_MATCHER_i_17 ));
    LocalMux I__2814 (
            .O(N__20786),
            .I(\c0.FRAME_MATCHER_i_17 ));
    InMux I__2813 (
            .O(N__20781),
            .I(N__20778));
    LocalMux I__2812 (
            .O(N__20778),
            .I(N__20775));
    Span4Mux_v I__2811 (
            .O(N__20775),
            .I(N__20772));
    Odrv4 I__2810 (
            .O(N__20772),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_17 ));
    SRMux I__2809 (
            .O(N__20769),
            .I(N__20766));
    LocalMux I__2808 (
            .O(N__20766),
            .I(N__20763));
    Span12Mux_s4_h I__2807 (
            .O(N__20763),
            .I(N__20760));
    Odrv12 I__2806 (
            .O(N__20760),
            .I(\c0.n3_adj_2248 ));
    SRMux I__2805 (
            .O(N__20757),
            .I(N__20754));
    LocalMux I__2804 (
            .O(N__20754),
            .I(N__20751));
    Span4Mux_s1_h I__2803 (
            .O(N__20751),
            .I(N__20748));
    Span4Mux_h I__2802 (
            .O(N__20748),
            .I(N__20745));
    Odrv4 I__2801 (
            .O(N__20745),
            .I(\c0.n3_adj_2250 ));
    InMux I__2800 (
            .O(N__20742),
            .I(n16005));
    InMux I__2799 (
            .O(N__20739),
            .I(n16006));
    InMux I__2798 (
            .O(N__20736),
            .I(n16007));
    InMux I__2797 (
            .O(N__20733),
            .I(n16008));
    InMux I__2796 (
            .O(N__20730),
            .I(n16009));
    InMux I__2795 (
            .O(N__20727),
            .I(N__20724));
    LocalMux I__2794 (
            .O(N__20724),
            .I(\c0.n3 ));
    CascadeMux I__2793 (
            .O(N__20721),
            .I(\c0.n26_adj_2373_cascade_ ));
    SRMux I__2792 (
            .O(N__20718),
            .I(N__20715));
    LocalMux I__2791 (
            .O(N__20715),
            .I(N__20712));
    Sp12to4 I__2790 (
            .O(N__20712),
            .I(N__20709));
    Odrv12 I__2789 (
            .O(N__20709),
            .I(\c0.n3_adj_2280 ));
    InMux I__2788 (
            .O(N__20706),
            .I(n15996));
    InMux I__2787 (
            .O(N__20703),
            .I(n15997));
    InMux I__2786 (
            .O(N__20700),
            .I(n15998));
    InMux I__2785 (
            .O(N__20697),
            .I(n15999));
    InMux I__2784 (
            .O(N__20694),
            .I(n16000));
    InMux I__2783 (
            .O(N__20691),
            .I(n16001));
    InMux I__2782 (
            .O(N__20688),
            .I(bfn_5_26_0_));
    InMux I__2781 (
            .O(N__20685),
            .I(n16003));
    InMux I__2780 (
            .O(N__20682),
            .I(n16004));
    InMux I__2779 (
            .O(N__20679),
            .I(n15987));
    InMux I__2778 (
            .O(N__20676),
            .I(n15988));
    InMux I__2777 (
            .O(N__20673),
            .I(n15989));
    InMux I__2776 (
            .O(N__20670),
            .I(n15990));
    InMux I__2775 (
            .O(N__20667),
            .I(n15991));
    InMux I__2774 (
            .O(N__20664),
            .I(n15992));
    InMux I__2773 (
            .O(N__20661),
            .I(n15993));
    InMux I__2772 (
            .O(N__20658),
            .I(bfn_5_25_0_));
    InMux I__2771 (
            .O(N__20655),
            .I(n15995));
    InMux I__2770 (
            .O(N__20652),
            .I(bfn_5_23_0_));
    InMux I__2769 (
            .O(N__20649),
            .I(n15979));
    InMux I__2768 (
            .O(N__20646),
            .I(n15980));
    InMux I__2767 (
            .O(N__20643),
            .I(n15981));
    InMux I__2766 (
            .O(N__20640),
            .I(n15982));
    InMux I__2765 (
            .O(N__20637),
            .I(n15983));
    InMux I__2764 (
            .O(N__20634),
            .I(n15984));
    InMux I__2763 (
            .O(N__20631),
            .I(n15985));
    InMux I__2762 (
            .O(N__20628),
            .I(bfn_5_24_0_));
    CascadeMux I__2761 (
            .O(N__20625),
            .I(N__20621));
    InMux I__2760 (
            .O(N__20624),
            .I(N__20616));
    InMux I__2759 (
            .O(N__20621),
            .I(N__20613));
    InMux I__2758 (
            .O(N__20620),
            .I(N__20609));
    InMux I__2757 (
            .O(N__20619),
            .I(N__20606));
    LocalMux I__2756 (
            .O(N__20616),
            .I(N__20601));
    LocalMux I__2755 (
            .O(N__20613),
            .I(N__20601));
    InMux I__2754 (
            .O(N__20612),
            .I(N__20598));
    LocalMux I__2753 (
            .O(N__20609),
            .I(N__20595));
    LocalMux I__2752 (
            .O(N__20606),
            .I(N__20592));
    Span4Mux_h I__2751 (
            .O(N__20601),
            .I(N__20589));
    LocalMux I__2750 (
            .O(N__20598),
            .I(data_out_frame2_15_2));
    Odrv4 I__2749 (
            .O(N__20595),
            .I(data_out_frame2_15_2));
    Odrv4 I__2748 (
            .O(N__20592),
            .I(data_out_frame2_15_2));
    Odrv4 I__2747 (
            .O(N__20589),
            .I(data_out_frame2_15_2));
    InMux I__2746 (
            .O(N__20580),
            .I(N__20577));
    LocalMux I__2745 (
            .O(N__20577),
            .I(N__20573));
    InMux I__2744 (
            .O(N__20576),
            .I(N__20570));
    Span4Mux_s3_h I__2743 (
            .O(N__20573),
            .I(N__20567));
    LocalMux I__2742 (
            .O(N__20570),
            .I(data_out_frame2_18_2));
    Odrv4 I__2741 (
            .O(N__20567),
            .I(data_out_frame2_18_2));
    InMux I__2740 (
            .O(N__20562),
            .I(N__20558));
    InMux I__2739 (
            .O(N__20561),
            .I(N__20554));
    LocalMux I__2738 (
            .O(N__20558),
            .I(N__20551));
    InMux I__2737 (
            .O(N__20557),
            .I(N__20548));
    LocalMux I__2736 (
            .O(N__20554),
            .I(N__20544));
    Span4Mux_v I__2735 (
            .O(N__20551),
            .I(N__20539));
    LocalMux I__2734 (
            .O(N__20548),
            .I(N__20539));
    InMux I__2733 (
            .O(N__20547),
            .I(N__20536));
    Span4Mux_h I__2732 (
            .O(N__20544),
            .I(N__20531));
    Span4Mux_h I__2731 (
            .O(N__20539),
            .I(N__20531));
    LocalMux I__2730 (
            .O(N__20536),
            .I(data_out_frame2_16_5));
    Odrv4 I__2729 (
            .O(N__20531),
            .I(data_out_frame2_16_5));
    CascadeMux I__2728 (
            .O(N__20526),
            .I(N__20522));
    InMux I__2727 (
            .O(N__20525),
            .I(N__20518));
    InMux I__2726 (
            .O(N__20522),
            .I(N__20514));
    InMux I__2725 (
            .O(N__20521),
            .I(N__20510));
    LocalMux I__2724 (
            .O(N__20518),
            .I(N__20507));
    InMux I__2723 (
            .O(N__20517),
            .I(N__20504));
    LocalMux I__2722 (
            .O(N__20514),
            .I(N__20501));
    InMux I__2721 (
            .O(N__20513),
            .I(N__20498));
    LocalMux I__2720 (
            .O(N__20510),
            .I(N__20495));
    Span4Mux_s2_h I__2719 (
            .O(N__20507),
            .I(N__20490));
    LocalMux I__2718 (
            .O(N__20504),
            .I(N__20490));
    Span4Mux_h I__2717 (
            .O(N__20501),
            .I(N__20487));
    LocalMux I__2716 (
            .O(N__20498),
            .I(data_out_frame2_15_4));
    Odrv12 I__2715 (
            .O(N__20495),
            .I(data_out_frame2_15_4));
    Odrv4 I__2714 (
            .O(N__20490),
            .I(data_out_frame2_15_4));
    Odrv4 I__2713 (
            .O(N__20487),
            .I(data_out_frame2_15_4));
    InMux I__2712 (
            .O(N__20478),
            .I(N__20475));
    LocalMux I__2711 (
            .O(N__20475),
            .I(N__20471));
    InMux I__2710 (
            .O(N__20474),
            .I(N__20468));
    Odrv4 I__2709 (
            .O(N__20471),
            .I(\c0.n17156 ));
    LocalMux I__2708 (
            .O(N__20468),
            .I(\c0.n17156 ));
    CascadeMux I__2707 (
            .O(N__20463),
            .I(\c0.n6_adj_2182_cascade_ ));
    InMux I__2706 (
            .O(N__20460),
            .I(N__20457));
    LocalMux I__2705 (
            .O(N__20457),
            .I(N__20454));
    Span4Mux_v I__2704 (
            .O(N__20454),
            .I(N__20450));
    InMux I__2703 (
            .O(N__20453),
            .I(N__20447));
    Odrv4 I__2702 (
            .O(N__20450),
            .I(\c0.n10229 ));
    LocalMux I__2701 (
            .O(N__20447),
            .I(\c0.n10229 ));
    CascadeMux I__2700 (
            .O(N__20442),
            .I(n10725_cascade_));
    CascadeMux I__2699 (
            .O(N__20439),
            .I(N__20435));
    CascadeMux I__2698 (
            .O(N__20438),
            .I(N__20432));
    InMux I__2697 (
            .O(N__20435),
            .I(N__20428));
    InMux I__2696 (
            .O(N__20432),
            .I(N__20425));
    InMux I__2695 (
            .O(N__20431),
            .I(N__20421));
    LocalMux I__2694 (
            .O(N__20428),
            .I(N__20418));
    LocalMux I__2693 (
            .O(N__20425),
            .I(N__20415));
    InMux I__2692 (
            .O(N__20424),
            .I(N__20412));
    LocalMux I__2691 (
            .O(N__20421),
            .I(N__20409));
    Span4Mux_s1_h I__2690 (
            .O(N__20418),
            .I(N__20404));
    Span4Mux_v I__2689 (
            .O(N__20415),
            .I(N__20404));
    LocalMux I__2688 (
            .O(N__20412),
            .I(data_out_frame2_12_7));
    Odrv4 I__2687 (
            .O(N__20409),
            .I(data_out_frame2_12_7));
    Odrv4 I__2686 (
            .O(N__20404),
            .I(data_out_frame2_12_7));
    CascadeMux I__2685 (
            .O(N__20397),
            .I(N__20392));
    CascadeMux I__2684 (
            .O(N__20396),
            .I(N__20389));
    InMux I__2683 (
            .O(N__20395),
            .I(N__20386));
    InMux I__2682 (
            .O(N__20392),
            .I(N__20383));
    InMux I__2681 (
            .O(N__20389),
            .I(N__20380));
    LocalMux I__2680 (
            .O(N__20386),
            .I(N__20376));
    LocalMux I__2679 (
            .O(N__20383),
            .I(N__20373));
    LocalMux I__2678 (
            .O(N__20380),
            .I(N__20370));
    InMux I__2677 (
            .O(N__20379),
            .I(N__20367));
    Span4Mux_h I__2676 (
            .O(N__20376),
            .I(N__20364));
    Span4Mux_v I__2675 (
            .O(N__20373),
            .I(N__20359));
    Span4Mux_s1_h I__2674 (
            .O(N__20370),
            .I(N__20359));
    LocalMux I__2673 (
            .O(N__20367),
            .I(data_out_frame2_10_3));
    Odrv4 I__2672 (
            .O(N__20364),
            .I(data_out_frame2_10_3));
    Odrv4 I__2671 (
            .O(N__20359),
            .I(data_out_frame2_10_3));
    InMux I__2670 (
            .O(N__20352),
            .I(N__20349));
    LocalMux I__2669 (
            .O(N__20349),
            .I(N__20346));
    Span4Mux_h I__2668 (
            .O(N__20346),
            .I(N__20343));
    Odrv4 I__2667 (
            .O(N__20343),
            .I(\c0.n18106 ));
    InMux I__2666 (
            .O(N__20340),
            .I(N__20336));
    InMux I__2665 (
            .O(N__20339),
            .I(N__20333));
    LocalMux I__2664 (
            .O(N__20336),
            .I(N__20327));
    LocalMux I__2663 (
            .O(N__20333),
            .I(N__20327));
    InMux I__2662 (
            .O(N__20332),
            .I(N__20324));
    Span4Mux_v I__2661 (
            .O(N__20327),
            .I(N__20319));
    LocalMux I__2660 (
            .O(N__20324),
            .I(N__20316));
    InMux I__2659 (
            .O(N__20323),
            .I(N__20313));
    InMux I__2658 (
            .O(N__20322),
            .I(N__20310));
    Span4Mux_s2_h I__2657 (
            .O(N__20319),
            .I(N__20307));
    Span4Mux_h I__2656 (
            .O(N__20316),
            .I(N__20304));
    LocalMux I__2655 (
            .O(N__20313),
            .I(N__20301));
    LocalMux I__2654 (
            .O(N__20310),
            .I(data_out_frame2_16_2));
    Odrv4 I__2653 (
            .O(N__20307),
            .I(data_out_frame2_16_2));
    Odrv4 I__2652 (
            .O(N__20304),
            .I(data_out_frame2_16_2));
    Odrv4 I__2651 (
            .O(N__20301),
            .I(data_out_frame2_16_2));
    CascadeMux I__2650 (
            .O(N__20292),
            .I(N__20289));
    InMux I__2649 (
            .O(N__20289),
            .I(N__20285));
    InMux I__2648 (
            .O(N__20288),
            .I(N__20281));
    LocalMux I__2647 (
            .O(N__20285),
            .I(N__20278));
    InMux I__2646 (
            .O(N__20284),
            .I(N__20275));
    LocalMux I__2645 (
            .O(N__20281),
            .I(N__20272));
    Odrv4 I__2644 (
            .O(N__20278),
            .I(\c0.n10263 ));
    LocalMux I__2643 (
            .O(N__20275),
            .I(\c0.n10263 ));
    Odrv4 I__2642 (
            .O(N__20272),
            .I(\c0.n10263 ));
    InMux I__2641 (
            .O(N__20265),
            .I(N__20262));
    LocalMux I__2640 (
            .O(N__20262),
            .I(N__20259));
    Odrv4 I__2639 (
            .O(N__20259),
            .I(\c0.n15_adj_2205 ));
    InMux I__2638 (
            .O(N__20256),
            .I(N__20253));
    LocalMux I__2637 (
            .O(N__20253),
            .I(N__20250));
    Span4Mux_v I__2636 (
            .O(N__20250),
            .I(N__20247));
    Span4Mux_h I__2635 (
            .O(N__20247),
            .I(N__20244));
    Odrv4 I__2634 (
            .O(N__20244),
            .I(\c0.n5_adj_2337 ));
    InMux I__2633 (
            .O(N__20241),
            .I(N__20235));
    InMux I__2632 (
            .O(N__20240),
            .I(N__20235));
    LocalMux I__2631 (
            .O(N__20235),
            .I(N__20231));
    InMux I__2630 (
            .O(N__20234),
            .I(N__20226));
    Span4Mux_s3_h I__2629 (
            .O(N__20231),
            .I(N__20223));
    InMux I__2628 (
            .O(N__20230),
            .I(N__20220));
    InMux I__2627 (
            .O(N__20229),
            .I(N__20217));
    LocalMux I__2626 (
            .O(N__20226),
            .I(data_out_frame2_10_2));
    Odrv4 I__2625 (
            .O(N__20223),
            .I(data_out_frame2_10_2));
    LocalMux I__2624 (
            .O(N__20220),
            .I(data_out_frame2_10_2));
    LocalMux I__2623 (
            .O(N__20217),
            .I(data_out_frame2_10_2));
    InMux I__2622 (
            .O(N__20208),
            .I(N__20204));
    InMux I__2621 (
            .O(N__20207),
            .I(N__20201));
    LocalMux I__2620 (
            .O(N__20204),
            .I(N__20198));
    LocalMux I__2619 (
            .O(N__20201),
            .I(N__20195));
    Span4Mux_s3_h I__2618 (
            .O(N__20198),
            .I(N__20190));
    Span4Mux_v I__2617 (
            .O(N__20195),
            .I(N__20190));
    Odrv4 I__2616 (
            .O(N__20190),
            .I(\c0.n10492 ));
    CascadeMux I__2615 (
            .O(N__20187),
            .I(N__20184));
    InMux I__2614 (
            .O(N__20184),
            .I(N__20179));
    InMux I__2613 (
            .O(N__20183),
            .I(N__20174));
    InMux I__2612 (
            .O(N__20182),
            .I(N__20174));
    LocalMux I__2611 (
            .O(N__20179),
            .I(N__20171));
    LocalMux I__2610 (
            .O(N__20174),
            .I(N__20168));
    Span4Mux_s2_h I__2609 (
            .O(N__20171),
            .I(N__20161));
    Span4Mux_h I__2608 (
            .O(N__20168),
            .I(N__20161));
    InMux I__2607 (
            .O(N__20167),
            .I(N__20158));
    InMux I__2606 (
            .O(N__20166),
            .I(N__20155));
    Span4Mux_v I__2605 (
            .O(N__20161),
            .I(N__20152));
    LocalMux I__2604 (
            .O(N__20158),
            .I(data_out_frame2_12_5));
    LocalMux I__2603 (
            .O(N__20155),
            .I(data_out_frame2_12_5));
    Odrv4 I__2602 (
            .O(N__20152),
            .I(data_out_frame2_12_5));
    InMux I__2601 (
            .O(N__20145),
            .I(N__20142));
    LocalMux I__2600 (
            .O(N__20142),
            .I(N__20139));
    Span4Mux_v I__2599 (
            .O(N__20139),
            .I(N__20135));
    InMux I__2598 (
            .O(N__20138),
            .I(N__20132));
    Span4Mux_s1_h I__2597 (
            .O(N__20135),
            .I(N__20129));
    LocalMux I__2596 (
            .O(N__20132),
            .I(\c0.n17255 ));
    Odrv4 I__2595 (
            .O(N__20129),
            .I(\c0.n17255 ));
    InMux I__2594 (
            .O(N__20124),
            .I(N__20120));
    InMux I__2593 (
            .O(N__20123),
            .I(N__20117));
    LocalMux I__2592 (
            .O(N__20120),
            .I(N__20114));
    LocalMux I__2591 (
            .O(N__20117),
            .I(N__20110));
    Span4Mux_v I__2590 (
            .O(N__20114),
            .I(N__20107));
    InMux I__2589 (
            .O(N__20113),
            .I(N__20103));
    Span4Mux_v I__2588 (
            .O(N__20110),
            .I(N__20098));
    Span4Mux_s2_h I__2587 (
            .O(N__20107),
            .I(N__20098));
    InMux I__2586 (
            .O(N__20106),
            .I(N__20095));
    LocalMux I__2585 (
            .O(N__20103),
            .I(data_out_frame2_16_4));
    Odrv4 I__2584 (
            .O(N__20098),
            .I(data_out_frame2_16_4));
    LocalMux I__2583 (
            .O(N__20095),
            .I(data_out_frame2_16_4));
    CascadeMux I__2582 (
            .O(N__20088),
            .I(N__20084));
    InMux I__2581 (
            .O(N__20087),
            .I(N__20081));
    InMux I__2580 (
            .O(N__20084),
            .I(N__20077));
    LocalMux I__2579 (
            .O(N__20081),
            .I(N__20074));
    CascadeMux I__2578 (
            .O(N__20080),
            .I(N__20071));
    LocalMux I__2577 (
            .O(N__20077),
            .I(N__20068));
    Span4Mux_v I__2576 (
            .O(N__20074),
            .I(N__20065));
    InMux I__2575 (
            .O(N__20071),
            .I(N__20061));
    Span4Mux_h I__2574 (
            .O(N__20068),
            .I(N__20058));
    Span4Mux_h I__2573 (
            .O(N__20065),
            .I(N__20055));
    InMux I__2572 (
            .O(N__20064),
            .I(N__20052));
    LocalMux I__2571 (
            .O(N__20061),
            .I(data_out_frame2_11_1));
    Odrv4 I__2570 (
            .O(N__20058),
            .I(data_out_frame2_11_1));
    Odrv4 I__2569 (
            .O(N__20055),
            .I(data_out_frame2_11_1));
    LocalMux I__2568 (
            .O(N__20052),
            .I(data_out_frame2_11_1));
    InMux I__2567 (
            .O(N__20043),
            .I(N__20040));
    LocalMux I__2566 (
            .O(N__20040),
            .I(N__20037));
    Odrv4 I__2565 (
            .O(N__20037),
            .I(\c0.n17288 ));
    InMux I__2564 (
            .O(N__20034),
            .I(N__20031));
    LocalMux I__2563 (
            .O(N__20031),
            .I(N__20027));
    InMux I__2562 (
            .O(N__20030),
            .I(N__20023));
    Span4Mux_v I__2561 (
            .O(N__20027),
            .I(N__20020));
    CascadeMux I__2560 (
            .O(N__20026),
            .I(N__20016));
    LocalMux I__2559 (
            .O(N__20023),
            .I(N__20013));
    Sp12to4 I__2558 (
            .O(N__20020),
            .I(N__20008));
    InMux I__2557 (
            .O(N__20019),
            .I(N__20005));
    InMux I__2556 (
            .O(N__20016),
            .I(N__20002));
    Span4Mux_s2_h I__2555 (
            .O(N__20013),
            .I(N__19999));
    InMux I__2554 (
            .O(N__20012),
            .I(N__19994));
    InMux I__2553 (
            .O(N__20011),
            .I(N__19994));
    Span12Mux_h I__2552 (
            .O(N__20008),
            .I(N__19989));
    LocalMux I__2551 (
            .O(N__20005),
            .I(N__19989));
    LocalMux I__2550 (
            .O(N__20002),
            .I(data_out_frame2_12_4));
    Odrv4 I__2549 (
            .O(N__19999),
            .I(data_out_frame2_12_4));
    LocalMux I__2548 (
            .O(N__19994),
            .I(data_out_frame2_12_4));
    Odrv12 I__2547 (
            .O(N__19989),
            .I(data_out_frame2_12_4));
    CascadeMux I__2546 (
            .O(N__19980),
            .I(\c0.n17288_cascade_ ));
    InMux I__2545 (
            .O(N__19977),
            .I(N__19974));
    LocalMux I__2544 (
            .O(N__19974),
            .I(\c0.n14_adj_2292 ));
    CascadeMux I__2543 (
            .O(N__19971),
            .I(N__19967));
    InMux I__2542 (
            .O(N__19970),
            .I(N__19964));
    InMux I__2541 (
            .O(N__19967),
            .I(N__19961));
    LocalMux I__2540 (
            .O(N__19964),
            .I(\c0.n17294 ));
    LocalMux I__2539 (
            .O(N__19961),
            .I(\c0.n17294 ));
    CascadeMux I__2538 (
            .O(N__19956),
            .I(\c0.n10428_cascade_ ));
    InMux I__2537 (
            .O(N__19953),
            .I(N__19950));
    LocalMux I__2536 (
            .O(N__19950),
            .I(N__19947));
    Span4Mux_h I__2535 (
            .O(N__19947),
            .I(N__19944));
    Odrv4 I__2534 (
            .O(N__19944),
            .I(\c0.n12_adj_2178 ));
    CascadeMux I__2533 (
            .O(N__19941),
            .I(N__19938));
    InMux I__2532 (
            .O(N__19938),
            .I(N__19935));
    LocalMux I__2531 (
            .O(N__19935),
            .I(N__19932));
    Span4Mux_h I__2530 (
            .O(N__19932),
            .I(N__19929));
    Odrv4 I__2529 (
            .O(N__19929),
            .I(\c0.n10504 ));
    InMux I__2528 (
            .O(N__19926),
            .I(N__19923));
    LocalMux I__2527 (
            .O(N__19923),
            .I(N__19919));
    InMux I__2526 (
            .O(N__19922),
            .I(N__19916));
    Span4Mux_v I__2525 (
            .O(N__19919),
            .I(N__19913));
    LocalMux I__2524 (
            .O(N__19916),
            .I(N__19908));
    Span4Mux_s3_h I__2523 (
            .O(N__19913),
            .I(N__19908));
    Odrv4 I__2522 (
            .O(N__19908),
            .I(data_out_frame2_17_1));
    InMux I__2521 (
            .O(N__19905),
            .I(N__19900));
    InMux I__2520 (
            .O(N__19904),
            .I(N__19897));
    CascadeMux I__2519 (
            .O(N__19903),
            .I(N__19894));
    LocalMux I__2518 (
            .O(N__19900),
            .I(N__19891));
    LocalMux I__2517 (
            .O(N__19897),
            .I(N__19888));
    InMux I__2516 (
            .O(N__19894),
            .I(N__19885));
    Span4Mux_v I__2515 (
            .O(N__19891),
            .I(N__19881));
    Span4Mux_v I__2514 (
            .O(N__19888),
            .I(N__19875));
    LocalMux I__2513 (
            .O(N__19885),
            .I(N__19875));
    InMux I__2512 (
            .O(N__19884),
            .I(N__19872));
    Span4Mux_s2_h I__2511 (
            .O(N__19881),
            .I(N__19869));
    InMux I__2510 (
            .O(N__19880),
            .I(N__19866));
    Span4Mux_v I__2509 (
            .O(N__19875),
            .I(N__19863));
    LocalMux I__2508 (
            .O(N__19872),
            .I(N__19858));
    Sp12to4 I__2507 (
            .O(N__19869),
            .I(N__19858));
    LocalMux I__2506 (
            .O(N__19866),
            .I(N__19855));
    Odrv4 I__2505 (
            .O(N__19863),
            .I(data_out_frame2_9_4));
    Odrv12 I__2504 (
            .O(N__19858),
            .I(data_out_frame2_9_4));
    Odrv4 I__2503 (
            .O(N__19855),
            .I(data_out_frame2_9_4));
    InMux I__2502 (
            .O(N__19848),
            .I(N__19845));
    LocalMux I__2501 (
            .O(N__19845),
            .I(N__19842));
    Span4Mux_h I__2500 (
            .O(N__19842),
            .I(N__19839));
    Odrv4 I__2499 (
            .O(N__19839),
            .I(\c0.n17568 ));
    InMux I__2498 (
            .O(N__19836),
            .I(N__19833));
    LocalMux I__2497 (
            .O(N__19833),
            .I(\c0.n10554 ));
    InMux I__2496 (
            .O(N__19830),
            .I(N__19826));
    InMux I__2495 (
            .O(N__19829),
            .I(N__19823));
    LocalMux I__2494 (
            .O(N__19826),
            .I(N__19820));
    LocalMux I__2493 (
            .O(N__19823),
            .I(N__19812));
    Span4Mux_v I__2492 (
            .O(N__19820),
            .I(N__19812));
    InMux I__2491 (
            .O(N__19819),
            .I(N__19809));
    InMux I__2490 (
            .O(N__19818),
            .I(N__19806));
    InMux I__2489 (
            .O(N__19817),
            .I(N__19803));
    Span4Mux_h I__2488 (
            .O(N__19812),
            .I(N__19796));
    LocalMux I__2487 (
            .O(N__19809),
            .I(N__19796));
    LocalMux I__2486 (
            .O(N__19806),
            .I(N__19796));
    LocalMux I__2485 (
            .O(N__19803),
            .I(data_out_frame2_5_6));
    Odrv4 I__2484 (
            .O(N__19796),
            .I(data_out_frame2_5_6));
    CascadeMux I__2483 (
            .O(N__19791),
            .I(\c0.n14_adj_2188_cascade_ ));
    InMux I__2482 (
            .O(N__19788),
            .I(N__19785));
    LocalMux I__2481 (
            .O(N__19785),
            .I(N__19782));
    Span4Mux_h I__2480 (
            .O(N__19782),
            .I(N__19779));
    Span4Mux_v I__2479 (
            .O(N__19779),
            .I(N__19776));
    Odrv4 I__2478 (
            .O(N__19776),
            .I(\c0.n15_adj_2185 ));
    CascadeMux I__2477 (
            .O(N__19773),
            .I(N__19770));
    InMux I__2476 (
            .O(N__19770),
            .I(N__19767));
    LocalMux I__2475 (
            .O(N__19767),
            .I(\c0.data_out_frame2_20_2 ));
    InMux I__2474 (
            .O(N__19764),
            .I(N__19759));
    InMux I__2473 (
            .O(N__19763),
            .I(N__19756));
    InMux I__2472 (
            .O(N__19762),
            .I(N__19753));
    LocalMux I__2471 (
            .O(N__19759),
            .I(N__19749));
    LocalMux I__2470 (
            .O(N__19756),
            .I(N__19746));
    LocalMux I__2469 (
            .O(N__19753),
            .I(N__19743));
    InMux I__2468 (
            .O(N__19752),
            .I(N__19740));
    Span4Mux_h I__2467 (
            .O(N__19749),
            .I(N__19737));
    Span4Mux_s3_h I__2466 (
            .O(N__19746),
            .I(N__19734));
    Span4Mux_s3_h I__2465 (
            .O(N__19743),
            .I(N__19731));
    LocalMux I__2464 (
            .O(N__19740),
            .I(data_out_frame2_7_4));
    Odrv4 I__2463 (
            .O(N__19737),
            .I(data_out_frame2_7_4));
    Odrv4 I__2462 (
            .O(N__19734),
            .I(data_out_frame2_7_4));
    Odrv4 I__2461 (
            .O(N__19731),
            .I(data_out_frame2_7_4));
    InMux I__2460 (
            .O(N__19722),
            .I(N__19719));
    LocalMux I__2459 (
            .O(N__19719),
            .I(\c0.n17240 ));
    CascadeMux I__2458 (
            .O(N__19716),
            .I(\c0.n17240_cascade_ ));
    InMux I__2457 (
            .O(N__19713),
            .I(N__19710));
    LocalMux I__2456 (
            .O(N__19710),
            .I(N__19707));
    Span12Mux_v I__2455 (
            .O(N__19707),
            .I(N__19704));
    Odrv12 I__2454 (
            .O(N__19704),
            .I(\c0.n14_adj_2206 ));
    CascadeMux I__2453 (
            .O(N__19701),
            .I(N__19698));
    InMux I__2452 (
            .O(N__19698),
            .I(N__19695));
    LocalMux I__2451 (
            .O(N__19695),
            .I(N__19692));
    Span12Mux_v I__2450 (
            .O(N__19692),
            .I(N__19689));
    Odrv12 I__2449 (
            .O(N__19689),
            .I(\c0.n17439 ));
    CascadeMux I__2448 (
            .O(N__19686),
            .I(N__19683));
    InMux I__2447 (
            .O(N__19683),
            .I(N__19680));
    LocalMux I__2446 (
            .O(N__19680),
            .I(\c0.n17249 ));
    CascadeMux I__2445 (
            .O(N__19677),
            .I(N__19674));
    InMux I__2444 (
            .O(N__19674),
            .I(N__19671));
    LocalMux I__2443 (
            .O(N__19671),
            .I(N__19668));
    Span12Mux_v I__2442 (
            .O(N__19668),
            .I(N__19665));
    Odrv12 I__2441 (
            .O(N__19665),
            .I(\c0.data_out_frame2_19_5 ));
    InMux I__2440 (
            .O(N__19662),
            .I(N__19658));
    InMux I__2439 (
            .O(N__19661),
            .I(N__19655));
    LocalMux I__2438 (
            .O(N__19658),
            .I(N__19652));
    LocalMux I__2437 (
            .O(N__19655),
            .I(N__19649));
    Span4Mux_h I__2436 (
            .O(N__19652),
            .I(N__19646));
    Span4Mux_h I__2435 (
            .O(N__19649),
            .I(N__19643));
    Odrv4 I__2434 (
            .O(N__19646),
            .I(\c0.n17116 ));
    Odrv4 I__2433 (
            .O(N__19643),
            .I(\c0.n17116 ));
    InMux I__2432 (
            .O(N__19638),
            .I(N__19635));
    LocalMux I__2431 (
            .O(N__19635),
            .I(N__19632));
    Span4Mux_h I__2430 (
            .O(N__19632),
            .I(N__19628));
    CascadeMux I__2429 (
            .O(N__19631),
            .I(N__19625));
    Span4Mux_h I__2428 (
            .O(N__19628),
            .I(N__19622));
    InMux I__2427 (
            .O(N__19625),
            .I(N__19619));
    Odrv4 I__2426 (
            .O(N__19622),
            .I(\c0.n17234 ));
    LocalMux I__2425 (
            .O(N__19619),
            .I(\c0.n17234 ));
    InMux I__2424 (
            .O(N__19614),
            .I(N__19611));
    LocalMux I__2423 (
            .O(N__19611),
            .I(\c0.n15_adj_2291 ));
    InMux I__2422 (
            .O(N__19608),
            .I(\c0.rx.n16125 ));
    InMux I__2421 (
            .O(N__19605),
            .I(\c0.rx.n16126 ));
    InMux I__2420 (
            .O(N__19602),
            .I(\c0.rx.n16127 ));
    InMux I__2419 (
            .O(N__19599),
            .I(\c0.rx.n16128 ));
    InMux I__2418 (
            .O(N__19596),
            .I(\c0.rx.n16129 ));
    InMux I__2417 (
            .O(N__19593),
            .I(\c0.rx.n16130 ));
    InMux I__2416 (
            .O(N__19590),
            .I(\c0.rx.n16131 ));
    InMux I__2415 (
            .O(N__19587),
            .I(N__19583));
    InMux I__2414 (
            .O(N__19586),
            .I(N__19580));
    LocalMux I__2413 (
            .O(N__19583),
            .I(N__19577));
    LocalMux I__2412 (
            .O(N__19580),
            .I(N__19572));
    Span4Mux_v I__2411 (
            .O(N__19577),
            .I(N__19572));
    Odrv4 I__2410 (
            .O(N__19572),
            .I(data_out_frame2_18_1));
    InMux I__2409 (
            .O(N__19569),
            .I(N__19566));
    LocalMux I__2408 (
            .O(N__19566),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_31 ));
    CascadeMux I__2407 (
            .O(N__19563),
            .I(n5244_cascade_));
    CascadeMux I__2406 (
            .O(N__19560),
            .I(n11018_cascade_));
    CascadeMux I__2405 (
            .O(N__19557),
            .I(N__19538));
    CascadeMux I__2404 (
            .O(N__19556),
            .I(N__19534));
    CascadeMux I__2403 (
            .O(N__19555),
            .I(N__19530));
    CascadeMux I__2402 (
            .O(N__19554),
            .I(N__19526));
    CascadeMux I__2401 (
            .O(N__19553),
            .I(N__19523));
    CascadeMux I__2400 (
            .O(N__19552),
            .I(N__19520));
    CascadeMux I__2399 (
            .O(N__19551),
            .I(N__19516));
    CascadeMux I__2398 (
            .O(N__19550),
            .I(N__19512));
    CascadeMux I__2397 (
            .O(N__19549),
            .I(N__19508));
    CascadeMux I__2396 (
            .O(N__19548),
            .I(N__19503));
    CascadeMux I__2395 (
            .O(N__19547),
            .I(N__19499));
    CascadeMux I__2394 (
            .O(N__19546),
            .I(N__19495));
    CascadeMux I__2393 (
            .O(N__19545),
            .I(N__19491));
    CascadeMux I__2392 (
            .O(N__19544),
            .I(N__19487));
    CascadeMux I__2391 (
            .O(N__19543),
            .I(N__19483));
    CascadeMux I__2390 (
            .O(N__19542),
            .I(N__19479));
    CascadeMux I__2389 (
            .O(N__19541),
            .I(N__19475));
    InMux I__2388 (
            .O(N__19538),
            .I(N__19472));
    InMux I__2387 (
            .O(N__19537),
            .I(N__19457));
    InMux I__2386 (
            .O(N__19534),
            .I(N__19457));
    InMux I__2385 (
            .O(N__19533),
            .I(N__19457));
    InMux I__2384 (
            .O(N__19530),
            .I(N__19457));
    InMux I__2383 (
            .O(N__19529),
            .I(N__19457));
    InMux I__2382 (
            .O(N__19526),
            .I(N__19457));
    InMux I__2381 (
            .O(N__19523),
            .I(N__19457));
    InMux I__2380 (
            .O(N__19520),
            .I(N__19440));
    InMux I__2379 (
            .O(N__19519),
            .I(N__19440));
    InMux I__2378 (
            .O(N__19516),
            .I(N__19440));
    InMux I__2377 (
            .O(N__19515),
            .I(N__19440));
    InMux I__2376 (
            .O(N__19512),
            .I(N__19440));
    InMux I__2375 (
            .O(N__19511),
            .I(N__19440));
    InMux I__2374 (
            .O(N__19508),
            .I(N__19440));
    InMux I__2373 (
            .O(N__19507),
            .I(N__19440));
    InMux I__2372 (
            .O(N__19506),
            .I(N__19423));
    InMux I__2371 (
            .O(N__19503),
            .I(N__19423));
    InMux I__2370 (
            .O(N__19502),
            .I(N__19423));
    InMux I__2369 (
            .O(N__19499),
            .I(N__19423));
    InMux I__2368 (
            .O(N__19498),
            .I(N__19423));
    InMux I__2367 (
            .O(N__19495),
            .I(N__19423));
    InMux I__2366 (
            .O(N__19494),
            .I(N__19423));
    InMux I__2365 (
            .O(N__19491),
            .I(N__19423));
    InMux I__2364 (
            .O(N__19490),
            .I(N__19406));
    InMux I__2363 (
            .O(N__19487),
            .I(N__19406));
    InMux I__2362 (
            .O(N__19486),
            .I(N__19406));
    InMux I__2361 (
            .O(N__19483),
            .I(N__19406));
    InMux I__2360 (
            .O(N__19482),
            .I(N__19406));
    InMux I__2359 (
            .O(N__19479),
            .I(N__19406));
    InMux I__2358 (
            .O(N__19478),
            .I(N__19406));
    InMux I__2357 (
            .O(N__19475),
            .I(N__19406));
    LocalMux I__2356 (
            .O(N__19472),
            .I(N__19397));
    LocalMux I__2355 (
            .O(N__19457),
            .I(N__19397));
    LocalMux I__2354 (
            .O(N__19440),
            .I(N__19397));
    LocalMux I__2353 (
            .O(N__19423),
            .I(N__19397));
    LocalMux I__2352 (
            .O(N__19406),
            .I(\c0.n18008 ));
    Odrv12 I__2351 (
            .O(N__19397),
            .I(\c0.n18008 ));
    CascadeMux I__2350 (
            .O(N__19392),
            .I(n13692_cascade_));
    InMux I__2349 (
            .O(N__19389),
            .I(bfn_4_32_0_));
    InMux I__2348 (
            .O(N__19386),
            .I(N__19383));
    LocalMux I__2347 (
            .O(N__19383),
            .I(N__19380));
    Span4Mux_s3_h I__2346 (
            .O(N__19380),
            .I(N__19377));
    Odrv4 I__2345 (
            .O(N__19377),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_23 ));
    InMux I__2344 (
            .O(N__19374),
            .I(\c0.n16101 ));
    InMux I__2343 (
            .O(N__19371),
            .I(bfn_4_30_0_));
    InMux I__2342 (
            .O(N__19368),
            .I(\c0.n16103 ));
    InMux I__2341 (
            .O(N__19365),
            .I(\c0.n16104 ));
    InMux I__2340 (
            .O(N__19362),
            .I(\c0.n16105 ));
    InMux I__2339 (
            .O(N__19359),
            .I(N__19356));
    LocalMux I__2338 (
            .O(N__19356),
            .I(N__19353));
    Odrv4 I__2337 (
            .O(N__19353),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_28 ));
    InMux I__2336 (
            .O(N__19350),
            .I(\c0.n16106 ));
    InMux I__2335 (
            .O(N__19347),
            .I(N__19344));
    LocalMux I__2334 (
            .O(N__19344),
            .I(N__19341));
    Span4Mux_s3_v I__2333 (
            .O(N__19341),
            .I(N__19338));
    Odrv4 I__2332 (
            .O(N__19338),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_29 ));
    CascadeMux I__2331 (
            .O(N__19335),
            .I(N__19332));
    InMux I__2330 (
            .O(N__19332),
            .I(N__19329));
    LocalMux I__2329 (
            .O(N__19329),
            .I(N__19323));
    InMux I__2328 (
            .O(N__19328),
            .I(N__19316));
    InMux I__2327 (
            .O(N__19327),
            .I(N__19316));
    InMux I__2326 (
            .O(N__19326),
            .I(N__19316));
    Odrv4 I__2325 (
            .O(N__19323),
            .I(\c0.FRAME_MATCHER_i_29 ));
    LocalMux I__2324 (
            .O(N__19316),
            .I(\c0.FRAME_MATCHER_i_29 ));
    InMux I__2323 (
            .O(N__19311),
            .I(N__19308));
    LocalMux I__2322 (
            .O(N__19308),
            .I(N__19305));
    Odrv4 I__2321 (
            .O(N__19305),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_29 ));
    InMux I__2320 (
            .O(N__19302),
            .I(\c0.n16107 ));
    InMux I__2319 (
            .O(N__19299),
            .I(N__19296));
    LocalMux I__2318 (
            .O(N__19296),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_30 ));
    InMux I__2317 (
            .O(N__19293),
            .I(\c0.n16108 ));
    InMux I__2316 (
            .O(N__19290),
            .I(\c0.n16109 ));
    InMux I__2315 (
            .O(N__19287),
            .I(N__19284));
    LocalMux I__2314 (
            .O(N__19284),
            .I(N__19281));
    Odrv4 I__2313 (
            .O(N__19281),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_14 ));
    InMux I__2312 (
            .O(N__19278),
            .I(\c0.n16092 ));
    InMux I__2311 (
            .O(N__19275),
            .I(N__19272));
    LocalMux I__2310 (
            .O(N__19272),
            .I(N__19269));
    Span4Mux_s3_h I__2309 (
            .O(N__19269),
            .I(N__19266));
    Odrv4 I__2308 (
            .O(N__19266),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_15 ));
    InMux I__2307 (
            .O(N__19263),
            .I(\c0.n16093 ));
    InMux I__2306 (
            .O(N__19260),
            .I(bfn_4_29_0_));
    InMux I__2305 (
            .O(N__19257),
            .I(\c0.n16095 ));
    InMux I__2304 (
            .O(N__19254),
            .I(\c0.n16096 ));
    InMux I__2303 (
            .O(N__19251),
            .I(N__19248));
    LocalMux I__2302 (
            .O(N__19248),
            .I(N__19245));
    Span4Mux_v I__2301 (
            .O(N__19245),
            .I(N__19242));
    Odrv4 I__2300 (
            .O(N__19242),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_19 ));
    InMux I__2299 (
            .O(N__19239),
            .I(\c0.n16097 ));
    InMux I__2298 (
            .O(N__19236),
            .I(N__19233));
    LocalMux I__2297 (
            .O(N__19233),
            .I(N__19230));
    Span4Mux_v I__2296 (
            .O(N__19230),
            .I(N__19227));
    Odrv4 I__2295 (
            .O(N__19227),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_20 ));
    InMux I__2294 (
            .O(N__19224),
            .I(\c0.n16098 ));
    InMux I__2293 (
            .O(N__19221),
            .I(N__19218));
    LocalMux I__2292 (
            .O(N__19218),
            .I(N__19215));
    Odrv4 I__2291 (
            .O(N__19215),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_21 ));
    InMux I__2290 (
            .O(N__19212),
            .I(\c0.n16099 ));
    InMux I__2289 (
            .O(N__19209),
            .I(N__19206));
    LocalMux I__2288 (
            .O(N__19206),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_22 ));
    InMux I__2287 (
            .O(N__19203),
            .I(\c0.n16100 ));
    InMux I__2286 (
            .O(N__19200),
            .I(\c0.n16084 ));
    InMux I__2285 (
            .O(N__19197),
            .I(N__19194));
    LocalMux I__2284 (
            .O(N__19194),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_7 ));
    InMux I__2283 (
            .O(N__19191),
            .I(\c0.n16085 ));
    InMux I__2282 (
            .O(N__19188),
            .I(N__19185));
    LocalMux I__2281 (
            .O(N__19185),
            .I(N__19182));
    Span4Mux_v I__2280 (
            .O(N__19182),
            .I(N__19179));
    Odrv4 I__2279 (
            .O(N__19179),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_8 ));
    InMux I__2278 (
            .O(N__19176),
            .I(bfn_4_28_0_));
    InMux I__2277 (
            .O(N__19173),
            .I(\c0.n16087 ));
    InMux I__2276 (
            .O(N__19170),
            .I(\c0.n16088 ));
    InMux I__2275 (
            .O(N__19167),
            .I(N__19164));
    LocalMux I__2274 (
            .O(N__19164),
            .I(N__19161));
    Span4Mux_v I__2273 (
            .O(N__19161),
            .I(N__19158));
    Odrv4 I__2272 (
            .O(N__19158),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_11 ));
    InMux I__2271 (
            .O(N__19155),
            .I(\c0.n16089 ));
    InMux I__2270 (
            .O(N__19152),
            .I(N__19149));
    LocalMux I__2269 (
            .O(N__19149),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_12 ));
    InMux I__2268 (
            .O(N__19146),
            .I(\c0.n16090 ));
    InMux I__2267 (
            .O(N__19143),
            .I(N__19140));
    LocalMux I__2266 (
            .O(N__19140),
            .I(N__19137));
    Odrv4 I__2265 (
            .O(N__19137),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_13 ));
    InMux I__2264 (
            .O(N__19134),
            .I(\c0.n16091 ));
    SRMux I__2263 (
            .O(N__19131),
            .I(N__19128));
    LocalMux I__2262 (
            .O(N__19128),
            .I(N__19125));
    Span4Mux_s3_h I__2261 (
            .O(N__19125),
            .I(N__19122));
    Odrv4 I__2260 (
            .O(N__19122),
            .I(\c0.n3_adj_2179 ));
    InMux I__2259 (
            .O(N__19119),
            .I(N__19116));
    LocalMux I__2258 (
            .O(N__19116),
            .I(N__19113));
    Odrv4 I__2257 (
            .O(N__19113),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_0 ));
    InMux I__2256 (
            .O(N__19110),
            .I(bfn_4_27_0_));
    InMux I__2255 (
            .O(N__19107),
            .I(N__19104));
    LocalMux I__2254 (
            .O(N__19104),
            .I(N__19101));
    Span4Mux_h I__2253 (
            .O(N__19101),
            .I(N__19098));
    Odrv4 I__2252 (
            .O(N__19098),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_1 ));
    InMux I__2251 (
            .O(N__19095),
            .I(\c0.n16079 ));
    InMux I__2250 (
            .O(N__19092),
            .I(\c0.n16080 ));
    InMux I__2249 (
            .O(N__19089),
            .I(N__19086));
    LocalMux I__2248 (
            .O(N__19086),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_3 ));
    CascadeMux I__2247 (
            .O(N__19083),
            .I(N__19080));
    InMux I__2246 (
            .O(N__19080),
            .I(N__19076));
    InMux I__2245 (
            .O(N__19079),
            .I(N__19071));
    LocalMux I__2244 (
            .O(N__19076),
            .I(N__19068));
    InMux I__2243 (
            .O(N__19075),
            .I(N__19063));
    InMux I__2242 (
            .O(N__19074),
            .I(N__19063));
    LocalMux I__2241 (
            .O(N__19071),
            .I(\c0.FRAME_MATCHER_i_3 ));
    Odrv4 I__2240 (
            .O(N__19068),
            .I(\c0.FRAME_MATCHER_i_3 ));
    LocalMux I__2239 (
            .O(N__19063),
            .I(\c0.FRAME_MATCHER_i_3 ));
    InMux I__2238 (
            .O(N__19056),
            .I(N__19053));
    LocalMux I__2237 (
            .O(N__19053),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_3 ));
    InMux I__2236 (
            .O(N__19050),
            .I(\c0.n16081 ));
    InMux I__2235 (
            .O(N__19047),
            .I(N__19044));
    LocalMux I__2234 (
            .O(N__19044),
            .I(\c0.FRAME_MATCHER_i_31_N_1310_4 ));
    InMux I__2233 (
            .O(N__19041),
            .I(N__19035));
    InMux I__2232 (
            .O(N__19040),
            .I(N__19032));
    InMux I__2231 (
            .O(N__19039),
            .I(N__19027));
    InMux I__2230 (
            .O(N__19038),
            .I(N__19027));
    LocalMux I__2229 (
            .O(N__19035),
            .I(N__19024));
    LocalMux I__2228 (
            .O(N__19032),
            .I(N__19019));
    LocalMux I__2227 (
            .O(N__19027),
            .I(N__19019));
    Span4Mux_h I__2226 (
            .O(N__19024),
            .I(N__19016));
    Span4Mux_h I__2225 (
            .O(N__19019),
            .I(N__19013));
    Odrv4 I__2224 (
            .O(N__19016),
            .I(\c0.FRAME_MATCHER_i_4 ));
    Odrv4 I__2223 (
            .O(N__19013),
            .I(\c0.FRAME_MATCHER_i_4 ));
    InMux I__2222 (
            .O(N__19008),
            .I(N__19005));
    LocalMux I__2221 (
            .O(N__19005),
            .I(N__19002));
    Span4Mux_s3_h I__2220 (
            .O(N__19002),
            .I(N__18999));
    Odrv4 I__2219 (
            .O(N__18999),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_4 ));
    InMux I__2218 (
            .O(N__18996),
            .I(\c0.n16082 ));
    InMux I__2217 (
            .O(N__18993),
            .I(N__18990));
    LocalMux I__2216 (
            .O(N__18990),
            .I(\c0.n43 ));
    CascadeMux I__2215 (
            .O(N__18987),
            .I(N__18984));
    InMux I__2214 (
            .O(N__18984),
            .I(N__18978));
    InMux I__2213 (
            .O(N__18983),
            .I(N__18971));
    InMux I__2212 (
            .O(N__18982),
            .I(N__18971));
    InMux I__2211 (
            .O(N__18981),
            .I(N__18971));
    LocalMux I__2210 (
            .O(N__18978),
            .I(\c0.FRAME_MATCHER_i_5 ));
    LocalMux I__2209 (
            .O(N__18971),
            .I(\c0.FRAME_MATCHER_i_5 ));
    InMux I__2208 (
            .O(N__18966),
            .I(N__18963));
    LocalMux I__2207 (
            .O(N__18963),
            .I(\c0.FRAME_MATCHER_i_31_N_1278_5 ));
    InMux I__2206 (
            .O(N__18960),
            .I(\c0.n16083 ));
    InMux I__2205 (
            .O(N__18957),
            .I(N__18953));
    InMux I__2204 (
            .O(N__18956),
            .I(N__18947));
    LocalMux I__2203 (
            .O(N__18953),
            .I(N__18944));
    CascadeMux I__2202 (
            .O(N__18952),
            .I(N__18941));
    CascadeMux I__2201 (
            .O(N__18951),
            .I(N__18938));
    InMux I__2200 (
            .O(N__18950),
            .I(N__18935));
    LocalMux I__2199 (
            .O(N__18947),
            .I(N__18932));
    Span4Mux_v I__2198 (
            .O(N__18944),
            .I(N__18929));
    InMux I__2197 (
            .O(N__18941),
            .I(N__18926));
    InMux I__2196 (
            .O(N__18938),
            .I(N__18923));
    LocalMux I__2195 (
            .O(N__18935),
            .I(data_out_frame2_9_2));
    Odrv12 I__2194 (
            .O(N__18932),
            .I(data_out_frame2_9_2));
    Odrv4 I__2193 (
            .O(N__18929),
            .I(data_out_frame2_9_2));
    LocalMux I__2192 (
            .O(N__18926),
            .I(data_out_frame2_9_2));
    LocalMux I__2191 (
            .O(N__18923),
            .I(data_out_frame2_9_2));
    InMux I__2190 (
            .O(N__18912),
            .I(N__18909));
    LocalMux I__2189 (
            .O(N__18909),
            .I(N__18906));
    Span4Mux_v I__2188 (
            .O(N__18906),
            .I(N__18903));
    Odrv4 I__2187 (
            .O(N__18903),
            .I(\c0.n18046 ));
    InMux I__2186 (
            .O(N__18900),
            .I(N__18897));
    LocalMux I__2185 (
            .O(N__18897),
            .I(N__18894));
    Span4Mux_h I__2184 (
            .O(N__18894),
            .I(N__18890));
    InMux I__2183 (
            .O(N__18893),
            .I(N__18887));
    Odrv4 I__2182 (
            .O(N__18890),
            .I(\c0.n17165 ));
    LocalMux I__2181 (
            .O(N__18887),
            .I(\c0.n17165 ));
    CascadeMux I__2180 (
            .O(N__18882),
            .I(N__18879));
    InMux I__2179 (
            .O(N__18879),
            .I(N__18876));
    LocalMux I__2178 (
            .O(N__18876),
            .I(\c0.n10334 ));
    InMux I__2177 (
            .O(N__18873),
            .I(N__18870));
    LocalMux I__2176 (
            .O(N__18870),
            .I(\c0.n10223 ));
    InMux I__2175 (
            .O(N__18867),
            .I(N__18864));
    LocalMux I__2174 (
            .O(N__18864),
            .I(N__18861));
    Span4Mux_v I__2173 (
            .O(N__18861),
            .I(N__18858));
    Odrv4 I__2172 (
            .O(N__18858),
            .I(\c0.n10_adj_2190 ));
    SRMux I__2171 (
            .O(N__18855),
            .I(N__18852));
    LocalMux I__2170 (
            .O(N__18852),
            .I(N__18849));
    Span4Mux_h I__2169 (
            .O(N__18849),
            .I(N__18846));
    Odrv4 I__2168 (
            .O(N__18846),
            .I(\c0.n3_adj_2282 ));
    SRMux I__2167 (
            .O(N__18843),
            .I(N__18840));
    LocalMux I__2166 (
            .O(N__18840),
            .I(\c0.n3_adj_2227 ));
    InMux I__2165 (
            .O(N__18837),
            .I(N__18832));
    InMux I__2164 (
            .O(N__18836),
            .I(N__18829));
    InMux I__2163 (
            .O(N__18835),
            .I(N__18825));
    LocalMux I__2162 (
            .O(N__18832),
            .I(N__18822));
    LocalMux I__2161 (
            .O(N__18829),
            .I(N__18819));
    InMux I__2160 (
            .O(N__18828),
            .I(N__18815));
    LocalMux I__2159 (
            .O(N__18825),
            .I(N__18812));
    Span4Mux_s3_h I__2158 (
            .O(N__18822),
            .I(N__18809));
    Span4Mux_s3_h I__2157 (
            .O(N__18819),
            .I(N__18806));
    InMux I__2156 (
            .O(N__18818),
            .I(N__18803));
    LocalMux I__2155 (
            .O(N__18815),
            .I(data_out_frame2_7_6));
    Odrv4 I__2154 (
            .O(N__18812),
            .I(data_out_frame2_7_6));
    Odrv4 I__2153 (
            .O(N__18809),
            .I(data_out_frame2_7_6));
    Odrv4 I__2152 (
            .O(N__18806),
            .I(data_out_frame2_7_6));
    LocalMux I__2151 (
            .O(N__18803),
            .I(data_out_frame2_7_6));
    InMux I__2150 (
            .O(N__18792),
            .I(N__18788));
    InMux I__2149 (
            .O(N__18791),
            .I(N__18784));
    LocalMux I__2148 (
            .O(N__18788),
            .I(N__18781));
    InMux I__2147 (
            .O(N__18787),
            .I(N__18777));
    LocalMux I__2146 (
            .O(N__18784),
            .I(N__18774));
    Span4Mux_h I__2145 (
            .O(N__18781),
            .I(N__18771));
    InMux I__2144 (
            .O(N__18780),
            .I(N__18768));
    LocalMux I__2143 (
            .O(N__18777),
            .I(data_out_frame2_6_4));
    Odrv12 I__2142 (
            .O(N__18774),
            .I(data_out_frame2_6_4));
    Odrv4 I__2141 (
            .O(N__18771),
            .I(data_out_frame2_6_4));
    LocalMux I__2140 (
            .O(N__18768),
            .I(data_out_frame2_6_4));
    InMux I__2139 (
            .O(N__18759),
            .I(N__18756));
    LocalMux I__2138 (
            .O(N__18756),
            .I(\c0.n6_adj_2339 ));
    InMux I__2137 (
            .O(N__18753),
            .I(N__18750));
    LocalMux I__2136 (
            .O(N__18750),
            .I(N__18747));
    Span4Mux_h I__2135 (
            .O(N__18747),
            .I(N__18744));
    Span4Mux_h I__2134 (
            .O(N__18744),
            .I(N__18740));
    InMux I__2133 (
            .O(N__18743),
            .I(N__18737));
    Odrv4 I__2132 (
            .O(N__18740),
            .I(\c0.n10507 ));
    LocalMux I__2131 (
            .O(N__18737),
            .I(\c0.n10507 ));
    InMux I__2130 (
            .O(N__18732),
            .I(N__18727));
    InMux I__2129 (
            .O(N__18731),
            .I(N__18723));
    CascadeMux I__2128 (
            .O(N__18730),
            .I(N__18719));
    LocalMux I__2127 (
            .O(N__18727),
            .I(N__18716));
    InMux I__2126 (
            .O(N__18726),
            .I(N__18713));
    LocalMux I__2125 (
            .O(N__18723),
            .I(N__18709));
    InMux I__2124 (
            .O(N__18722),
            .I(N__18706));
    InMux I__2123 (
            .O(N__18719),
            .I(N__18703));
    Span4Mux_s2_h I__2122 (
            .O(N__18716),
            .I(N__18700));
    LocalMux I__2121 (
            .O(N__18713),
            .I(N__18697));
    InMux I__2120 (
            .O(N__18712),
            .I(N__18694));
    Span4Mux_h I__2119 (
            .O(N__18709),
            .I(N__18691));
    LocalMux I__2118 (
            .O(N__18706),
            .I(N__18682));
    LocalMux I__2117 (
            .O(N__18703),
            .I(N__18682));
    Sp12to4 I__2116 (
            .O(N__18700),
            .I(N__18682));
    Sp12to4 I__2115 (
            .O(N__18697),
            .I(N__18682));
    LocalMux I__2114 (
            .O(N__18694),
            .I(data_out_frame2_15_0));
    Odrv4 I__2113 (
            .O(N__18691),
            .I(data_out_frame2_15_0));
    Odrv12 I__2112 (
            .O(N__18682),
            .I(data_out_frame2_15_0));
    InMux I__2111 (
            .O(N__18675),
            .I(N__18672));
    LocalMux I__2110 (
            .O(N__18672),
            .I(N__18669));
    Odrv12 I__2109 (
            .O(N__18669),
            .I(\c0.n17273 ));
    InMux I__2108 (
            .O(N__18666),
            .I(N__18661));
    InMux I__2107 (
            .O(N__18665),
            .I(N__18658));
    InMux I__2106 (
            .O(N__18664),
            .I(N__18655));
    LocalMux I__2105 (
            .O(N__18661),
            .I(N__18650));
    LocalMux I__2104 (
            .O(N__18658),
            .I(N__18650));
    LocalMux I__2103 (
            .O(N__18655),
            .I(N__18646));
    Sp12to4 I__2102 (
            .O(N__18650),
            .I(N__18643));
    InMux I__2101 (
            .O(N__18649),
            .I(N__18640));
    Span4Mux_h I__2100 (
            .O(N__18646),
            .I(N__18637));
    Span12Mux_v I__2099 (
            .O(N__18643),
            .I(N__18634));
    LocalMux I__2098 (
            .O(N__18640),
            .I(data_out_frame2_6_7));
    Odrv4 I__2097 (
            .O(N__18637),
            .I(data_out_frame2_6_7));
    Odrv12 I__2096 (
            .O(N__18634),
            .I(data_out_frame2_6_7));
    InMux I__2095 (
            .O(N__18627),
            .I(N__18623));
    InMux I__2094 (
            .O(N__18626),
            .I(N__18620));
    LocalMux I__2093 (
            .O(N__18623),
            .I(N__18614));
    LocalMux I__2092 (
            .O(N__18620),
            .I(N__18611));
    InMux I__2091 (
            .O(N__18619),
            .I(N__18606));
    InMux I__2090 (
            .O(N__18618),
            .I(N__18606));
    InMux I__2089 (
            .O(N__18617),
            .I(N__18603));
    Span4Mux_v I__2088 (
            .O(N__18614),
            .I(N__18598));
    Span4Mux_s3_h I__2087 (
            .O(N__18611),
            .I(N__18598));
    LocalMux I__2086 (
            .O(N__18606),
            .I(N__18595));
    LocalMux I__2085 (
            .O(N__18603),
            .I(data_out_frame2_16_1));
    Odrv4 I__2084 (
            .O(N__18598),
            .I(data_out_frame2_16_1));
    Odrv4 I__2083 (
            .O(N__18595),
            .I(data_out_frame2_16_1));
    InMux I__2082 (
            .O(N__18588),
            .I(N__18585));
    LocalMux I__2081 (
            .O(N__18585),
            .I(N__18582));
    Odrv12 I__2080 (
            .O(N__18582),
            .I(\c0.n17153 ));
    InMux I__2079 (
            .O(N__18579),
            .I(N__18576));
    LocalMux I__2078 (
            .O(N__18576),
            .I(\c0.n17168 ));
    CascadeMux I__2077 (
            .O(N__18573),
            .I(\c0.n17153_cascade_ ));
    InMux I__2076 (
            .O(N__18570),
            .I(N__18567));
    LocalMux I__2075 (
            .O(N__18567),
            .I(\c0.n26_adj_2203 ));
    CascadeMux I__2074 (
            .O(N__18564),
            .I(N__18561));
    InMux I__2073 (
            .O(N__18561),
            .I(N__18557));
    InMux I__2072 (
            .O(N__18560),
            .I(N__18553));
    LocalMux I__2071 (
            .O(N__18557),
            .I(N__18550));
    InMux I__2070 (
            .O(N__18556),
            .I(N__18547));
    LocalMux I__2069 (
            .O(N__18553),
            .I(N__18542));
    Span4Mux_v I__2068 (
            .O(N__18550),
            .I(N__18542));
    LocalMux I__2067 (
            .O(N__18547),
            .I(N__18539));
    Span4Mux_v I__2066 (
            .O(N__18542),
            .I(N__18534));
    Span4Mux_s3_h I__2065 (
            .O(N__18539),
            .I(N__18531));
    InMux I__2064 (
            .O(N__18538),
            .I(N__18526));
    InMux I__2063 (
            .O(N__18537),
            .I(N__18526));
    Odrv4 I__2062 (
            .O(N__18534),
            .I(data_out_frame2_5_7));
    Odrv4 I__2061 (
            .O(N__18531),
            .I(data_out_frame2_5_7));
    LocalMux I__2060 (
            .O(N__18526),
            .I(data_out_frame2_5_7));
    InMux I__2059 (
            .O(N__18519),
            .I(N__18513));
    InMux I__2058 (
            .O(N__18518),
            .I(N__18510));
    CascadeMux I__2057 (
            .O(N__18517),
            .I(N__18507));
    InMux I__2056 (
            .O(N__18516),
            .I(N__18504));
    LocalMux I__2055 (
            .O(N__18513),
            .I(N__18501));
    LocalMux I__2054 (
            .O(N__18510),
            .I(N__18498));
    InMux I__2053 (
            .O(N__18507),
            .I(N__18495));
    LocalMux I__2052 (
            .O(N__18504),
            .I(data_out_frame2_13_3));
    Odrv4 I__2051 (
            .O(N__18501),
            .I(data_out_frame2_13_3));
    Odrv12 I__2050 (
            .O(N__18498),
            .I(data_out_frame2_13_3));
    LocalMux I__2049 (
            .O(N__18495),
            .I(data_out_frame2_13_3));
    InMux I__2048 (
            .O(N__18486),
            .I(N__18483));
    LocalMux I__2047 (
            .O(N__18483),
            .I(N__18479));
    InMux I__2046 (
            .O(N__18482),
            .I(N__18476));
    Span12Mux_s3_h I__2045 (
            .O(N__18479),
            .I(N__18473));
    LocalMux I__2044 (
            .O(N__18476),
            .I(data_out_frame2_18_4));
    Odrv12 I__2043 (
            .O(N__18473),
            .I(data_out_frame2_18_4));
    InMux I__2042 (
            .O(N__18468),
            .I(N__18465));
    LocalMux I__2041 (
            .O(N__18465),
            .I(N__18460));
    InMux I__2040 (
            .O(N__18464),
            .I(N__18457));
    InMux I__2039 (
            .O(N__18463),
            .I(N__18454));
    Span4Mux_s2_h I__2038 (
            .O(N__18460),
            .I(N__18450));
    LocalMux I__2037 (
            .O(N__18457),
            .I(N__18447));
    LocalMux I__2036 (
            .O(N__18454),
            .I(N__18444));
    InMux I__2035 (
            .O(N__18453),
            .I(N__18441));
    Span4Mux_v I__2034 (
            .O(N__18450),
            .I(N__18436));
    Span4Mux_v I__2033 (
            .O(N__18447),
            .I(N__18436));
    Span4Mux_v I__2032 (
            .O(N__18444),
            .I(N__18433));
    LocalMux I__2031 (
            .O(N__18441),
            .I(data_out_frame2_5_5));
    Odrv4 I__2030 (
            .O(N__18436),
            .I(data_out_frame2_5_5));
    Odrv4 I__2029 (
            .O(N__18433),
            .I(data_out_frame2_5_5));
    CascadeMux I__2028 (
            .O(N__18426),
            .I(N__18422));
    InMux I__2027 (
            .O(N__18425),
            .I(N__18418));
    InMux I__2026 (
            .O(N__18422),
            .I(N__18415));
    InMux I__2025 (
            .O(N__18421),
            .I(N__18412));
    LocalMux I__2024 (
            .O(N__18418),
            .I(N__18408));
    LocalMux I__2023 (
            .O(N__18415),
            .I(N__18405));
    LocalMux I__2022 (
            .O(N__18412),
            .I(N__18402));
    InMux I__2021 (
            .O(N__18411),
            .I(N__18399));
    Span4Mux_s3_h I__2020 (
            .O(N__18408),
            .I(N__18396));
    Span4Mux_s3_h I__2019 (
            .O(N__18405),
            .I(N__18391));
    Span4Mux_s3_h I__2018 (
            .O(N__18402),
            .I(N__18391));
    LocalMux I__2017 (
            .O(N__18399),
            .I(data_out_frame2_7_3));
    Odrv4 I__2016 (
            .O(N__18396),
            .I(data_out_frame2_7_3));
    Odrv4 I__2015 (
            .O(N__18391),
            .I(data_out_frame2_7_3));
    InMux I__2014 (
            .O(N__18384),
            .I(N__18381));
    LocalMux I__2013 (
            .O(N__18381),
            .I(N__18378));
    Sp12to4 I__2012 (
            .O(N__18378),
            .I(N__18374));
    InMux I__2011 (
            .O(N__18377),
            .I(N__18371));
    Span12Mux_v I__2010 (
            .O(N__18374),
            .I(N__18368));
    LocalMux I__2009 (
            .O(N__18371),
            .I(data_out_frame2_17_4));
    Odrv12 I__2008 (
            .O(N__18368),
            .I(data_out_frame2_17_4));
    InMux I__2007 (
            .O(N__18363),
            .I(N__18360));
    LocalMux I__2006 (
            .O(N__18360),
            .I(N__18356));
    InMux I__2005 (
            .O(N__18359),
            .I(N__18353));
    Span4Mux_v I__2004 (
            .O(N__18356),
            .I(N__18350));
    LocalMux I__2003 (
            .O(N__18353),
            .I(data_out_frame2_17_7));
    Odrv4 I__2002 (
            .O(N__18350),
            .I(data_out_frame2_17_7));
    InMux I__2001 (
            .O(N__18345),
            .I(N__18342));
    LocalMux I__2000 (
            .O(N__18342),
            .I(N__18339));
    Span4Mux_h I__1999 (
            .O(N__18339),
            .I(N__18336));
    Odrv4 I__1998 (
            .O(N__18336),
            .I(\c0.n10356 ));
    CascadeMux I__1997 (
            .O(N__18333),
            .I(N__18330));
    InMux I__1996 (
            .O(N__18330),
            .I(N__18327));
    LocalMux I__1995 (
            .O(N__18327),
            .I(N__18324));
    Span4Mux_v I__1994 (
            .O(N__18324),
            .I(N__18320));
    InMux I__1993 (
            .O(N__18323),
            .I(N__18317));
    Odrv4 I__1992 (
            .O(N__18320),
            .I(\c0.n10572 ));
    LocalMux I__1991 (
            .O(N__18317),
            .I(\c0.n10572 ));
    InMux I__1990 (
            .O(N__18312),
            .I(N__18309));
    LocalMux I__1989 (
            .O(N__18309),
            .I(N__18306));
    Odrv4 I__1988 (
            .O(N__18306),
            .I(\c0.n16_adj_2170 ));
    InMux I__1987 (
            .O(N__18303),
            .I(N__18300));
    LocalMux I__1986 (
            .O(N__18300),
            .I(N__18296));
    InMux I__1985 (
            .O(N__18299),
            .I(N__18292));
    Span4Mux_v I__1984 (
            .O(N__18296),
            .I(N__18289));
    InMux I__1983 (
            .O(N__18295),
            .I(N__18285));
    LocalMux I__1982 (
            .O(N__18292),
            .I(N__18280));
    Span4Mux_v I__1981 (
            .O(N__18289),
            .I(N__18280));
    InMux I__1980 (
            .O(N__18288),
            .I(N__18277));
    LocalMux I__1979 (
            .O(N__18285),
            .I(data_out_frame2_6_5));
    Odrv4 I__1978 (
            .O(N__18280),
            .I(data_out_frame2_6_5));
    LocalMux I__1977 (
            .O(N__18277),
            .I(data_out_frame2_6_5));
    CascadeMux I__1976 (
            .O(N__18270),
            .I(\c0.n16_adj_2320_cascade_ ));
    InMux I__1975 (
            .O(N__18267),
            .I(N__18264));
    LocalMux I__1974 (
            .O(N__18264),
            .I(N__18261));
    Span4Mux_h I__1973 (
            .O(N__18261),
            .I(N__18257));
    InMux I__1972 (
            .O(N__18260),
            .I(N__18254));
    Odrv4 I__1971 (
            .O(N__18257),
            .I(\c0.n17216 ));
    LocalMux I__1970 (
            .O(N__18254),
            .I(\c0.n17216 ));
    InMux I__1969 (
            .O(N__18249),
            .I(N__18246));
    LocalMux I__1968 (
            .O(N__18246),
            .I(N__18243));
    Odrv4 I__1967 (
            .O(N__18243),
            .I(\c0.data_out_frame2_19_1 ));
    InMux I__1966 (
            .O(N__18240),
            .I(N__18237));
    LocalMux I__1965 (
            .O(N__18237),
            .I(\c0.n18058 ));
    CascadeMux I__1964 (
            .O(N__18234),
            .I(\c0.n6_adj_2175_cascade_ ));
    InMux I__1963 (
            .O(N__18231),
            .I(N__18227));
    InMux I__1962 (
            .O(N__18230),
            .I(N__18224));
    LocalMux I__1961 (
            .O(N__18227),
            .I(N__18221));
    LocalMux I__1960 (
            .O(N__18224),
            .I(N__18218));
    Span4Mux_s3_h I__1959 (
            .O(N__18221),
            .I(N__18215));
    Odrv4 I__1958 (
            .O(N__18218),
            .I(\c0.n17258 ));
    Odrv4 I__1957 (
            .O(N__18215),
            .I(\c0.n17258 ));
    InMux I__1956 (
            .O(N__18210),
            .I(N__18207));
    LocalMux I__1955 (
            .O(N__18207),
            .I(N__18203));
    CascadeMux I__1954 (
            .O(N__18206),
            .I(N__18198));
    Span4Mux_s3_h I__1953 (
            .O(N__18203),
            .I(N__18194));
    InMux I__1952 (
            .O(N__18202),
            .I(N__18189));
    InMux I__1951 (
            .O(N__18201),
            .I(N__18189));
    InMux I__1950 (
            .O(N__18198),
            .I(N__18184));
    InMux I__1949 (
            .O(N__18197),
            .I(N__18184));
    Odrv4 I__1948 (
            .O(N__18194),
            .I(data_out_frame2_11_2));
    LocalMux I__1947 (
            .O(N__18189),
            .I(data_out_frame2_11_2));
    LocalMux I__1946 (
            .O(N__18184),
            .I(data_out_frame2_11_2));
    InMux I__1945 (
            .O(N__18177),
            .I(N__18173));
    InMux I__1944 (
            .O(N__18176),
            .I(N__18170));
    LocalMux I__1943 (
            .O(N__18173),
            .I(N__18165));
    LocalMux I__1942 (
            .O(N__18170),
            .I(N__18165));
    Span4Mux_v I__1941 (
            .O(N__18165),
            .I(N__18162));
    Odrv4 I__1940 (
            .O(N__18162),
            .I(\c0.n17171 ));
    CascadeMux I__1939 (
            .O(N__18159),
            .I(N__18156));
    InMux I__1938 (
            .O(N__18156),
            .I(N__18153));
    LocalMux I__1937 (
            .O(N__18153),
            .I(N__18150));
    Span4Mux_h I__1936 (
            .O(N__18150),
            .I(N__18147));
    Odrv4 I__1935 (
            .O(N__18147),
            .I(\c0.n17132 ));
    InMux I__1934 (
            .O(N__18144),
            .I(N__18141));
    LocalMux I__1933 (
            .O(N__18141),
            .I(N__18137));
    InMux I__1932 (
            .O(N__18140),
            .I(N__18134));
    Span4Mux_h I__1931 (
            .O(N__18137),
            .I(N__18131));
    LocalMux I__1930 (
            .O(N__18134),
            .I(N__18128));
    Odrv4 I__1929 (
            .O(N__18131),
            .I(\c0.n17184 ));
    Odrv4 I__1928 (
            .O(N__18128),
            .I(\c0.n17184 ));
    InMux I__1927 (
            .O(N__18123),
            .I(N__18120));
    LocalMux I__1926 (
            .O(N__18120),
            .I(\c0.n32 ));
    InMux I__1925 (
            .O(N__18117),
            .I(N__18114));
    LocalMux I__1924 (
            .O(N__18114),
            .I(N__18111));
    Span4Mux_h I__1923 (
            .O(N__18111),
            .I(N__18108));
    Span4Mux_s1_h I__1922 (
            .O(N__18108),
            .I(N__18105));
    Odrv4 I__1921 (
            .O(N__18105),
            .I(\c0.n10437 ));
    CascadeMux I__1920 (
            .O(N__18102),
            .I(\c0.n17249_cascade_ ));
    InMux I__1919 (
            .O(N__18099),
            .I(N__18096));
    LocalMux I__1918 (
            .O(N__18096),
            .I(N__18093));
    Span4Mux_v I__1917 (
            .O(N__18093),
            .I(N__18090));
    Odrv4 I__1916 (
            .O(N__18090),
            .I(\c0.n12_adj_2298 ));
    InMux I__1915 (
            .O(N__18087),
            .I(N__18081));
    InMux I__1914 (
            .O(N__18086),
            .I(N__18077));
    CascadeMux I__1913 (
            .O(N__18085),
            .I(N__18074));
    CascadeMux I__1912 (
            .O(N__18084),
            .I(N__18071));
    LocalMux I__1911 (
            .O(N__18081),
            .I(N__18068));
    InMux I__1910 (
            .O(N__18080),
            .I(N__18065));
    LocalMux I__1909 (
            .O(N__18077),
            .I(N__18062));
    InMux I__1908 (
            .O(N__18074),
            .I(N__18058));
    InMux I__1907 (
            .O(N__18071),
            .I(N__18055));
    Span4Mux_h I__1906 (
            .O(N__18068),
            .I(N__18052));
    LocalMux I__1905 (
            .O(N__18065),
            .I(N__18049));
    Span4Mux_v I__1904 (
            .O(N__18062),
            .I(N__18046));
    InMux I__1903 (
            .O(N__18061),
            .I(N__18043));
    LocalMux I__1902 (
            .O(N__18058),
            .I(data_out_frame2_8_1));
    LocalMux I__1901 (
            .O(N__18055),
            .I(data_out_frame2_8_1));
    Odrv4 I__1900 (
            .O(N__18052),
            .I(data_out_frame2_8_1));
    Odrv4 I__1899 (
            .O(N__18049),
            .I(data_out_frame2_8_1));
    Odrv4 I__1898 (
            .O(N__18046),
            .I(data_out_frame2_8_1));
    LocalMux I__1897 (
            .O(N__18043),
            .I(data_out_frame2_8_1));
    InMux I__1896 (
            .O(N__18030),
            .I(N__18027));
    LocalMux I__1895 (
            .O(N__18027),
            .I(N__18024));
    Span4Mux_v I__1894 (
            .O(N__18024),
            .I(N__18021));
    Span4Mux_s0_h I__1893 (
            .O(N__18021),
            .I(N__18018));
    Odrv4 I__1892 (
            .O(N__18018),
            .I(\c0.n20 ));
    InMux I__1891 (
            .O(N__18015),
            .I(N__18012));
    LocalMux I__1890 (
            .O(N__18012),
            .I(N__18009));
    Span4Mux_v I__1889 (
            .O(N__18009),
            .I(N__18006));
    Span4Mux_h I__1888 (
            .O(N__18006),
            .I(N__18003));
    Odrv4 I__1887 (
            .O(N__18003),
            .I(\c0.n17678 ));
    InMux I__1886 (
            .O(N__18000),
            .I(N__17996));
    InMux I__1885 (
            .O(N__17999),
            .I(N__17993));
    LocalMux I__1884 (
            .O(N__17996),
            .I(N__17990));
    LocalMux I__1883 (
            .O(N__17993),
            .I(N__17987));
    Span4Mux_v I__1882 (
            .O(N__17990),
            .I(N__17984));
    Span4Mux_v I__1881 (
            .O(N__17987),
            .I(N__17981));
    Span4Mux_h I__1880 (
            .O(N__17984),
            .I(N__17978));
    Odrv4 I__1879 (
            .O(N__17981),
            .I(\c0.n17279 ));
    Odrv4 I__1878 (
            .O(N__17978),
            .I(\c0.n17279 ));
    InMux I__1877 (
            .O(N__17973),
            .I(N__17970));
    LocalMux I__1876 (
            .O(N__17970),
            .I(N__17967));
    Sp12to4 I__1875 (
            .O(N__17967),
            .I(N__17964));
    Odrv12 I__1874 (
            .O(N__17964),
            .I(\c0.data_out_frame2_20_1 ));
    InMux I__1873 (
            .O(N__17961),
            .I(N__17953));
    InMux I__1872 (
            .O(N__17960),
            .I(N__17953));
    CascadeMux I__1871 (
            .O(N__17959),
            .I(N__17950));
    InMux I__1870 (
            .O(N__17958),
            .I(N__17947));
    LocalMux I__1869 (
            .O(N__17953),
            .I(N__17944));
    InMux I__1868 (
            .O(N__17950),
            .I(N__17941));
    LocalMux I__1867 (
            .O(N__17947),
            .I(N__17935));
    Span4Mux_v I__1866 (
            .O(N__17944),
            .I(N__17935));
    LocalMux I__1865 (
            .O(N__17941),
            .I(N__17932));
    InMux I__1864 (
            .O(N__17940),
            .I(N__17929));
    Span4Mux_h I__1863 (
            .O(N__17935),
            .I(N__17926));
    Span4Mux_h I__1862 (
            .O(N__17932),
            .I(N__17923));
    LocalMux I__1861 (
            .O(N__17929),
            .I(data_out_frame2_13_0));
    Odrv4 I__1860 (
            .O(N__17926),
            .I(data_out_frame2_13_0));
    Odrv4 I__1859 (
            .O(N__17923),
            .I(data_out_frame2_13_0));
    InMux I__1858 (
            .O(N__17916),
            .I(N__17913));
    LocalMux I__1857 (
            .O(N__17913),
            .I(N__17910));
    Span4Mux_h I__1856 (
            .O(N__17910),
            .I(N__17906));
    InMux I__1855 (
            .O(N__17909),
            .I(N__17903));
    Odrv4 I__1854 (
            .O(N__17906),
            .I(\c0.n10424 ));
    LocalMux I__1853 (
            .O(N__17903),
            .I(\c0.n10424 ));
    InMux I__1852 (
            .O(N__17898),
            .I(N__17895));
    LocalMux I__1851 (
            .O(N__17895),
            .I(N__17892));
    Span4Mux_v I__1850 (
            .O(N__17892),
            .I(N__17889));
    Odrv4 I__1849 (
            .O(N__17889),
            .I(\c0.n14_adj_2346 ));
    CascadeMux I__1848 (
            .O(N__17886),
            .I(\c0.n15_adj_2341_cascade_ ));
    InMux I__1847 (
            .O(N__17883),
            .I(N__17879));
    InMux I__1846 (
            .O(N__17882),
            .I(N__17876));
    LocalMux I__1845 (
            .O(N__17879),
            .I(N__17870));
    LocalMux I__1844 (
            .O(N__17876),
            .I(N__17870));
    InMux I__1843 (
            .O(N__17875),
            .I(N__17866));
    Span4Mux_v I__1842 (
            .O(N__17870),
            .I(N__17863));
    InMux I__1841 (
            .O(N__17869),
            .I(N__17860));
    LocalMux I__1840 (
            .O(N__17866),
            .I(data_out_frame2_14_5));
    Odrv4 I__1839 (
            .O(N__17863),
            .I(data_out_frame2_14_5));
    LocalMux I__1838 (
            .O(N__17860),
            .I(data_out_frame2_14_5));
    CascadeMux I__1837 (
            .O(N__17853),
            .I(\c0.n18178_cascade_ ));
    InMux I__1836 (
            .O(N__17850),
            .I(N__17847));
    LocalMux I__1835 (
            .O(N__17847),
            .I(N__17844));
    Span4Mux_h I__1834 (
            .O(N__17844),
            .I(N__17841));
    Span4Mux_v I__1833 (
            .O(N__17841),
            .I(N__17838));
    Odrv4 I__1832 (
            .O(N__17838),
            .I(\c0.n6_adj_2161 ));
    InMux I__1831 (
            .O(N__17835),
            .I(N__17832));
    LocalMux I__1830 (
            .O(N__17832),
            .I(\c0.n18181 ));
    InMux I__1829 (
            .O(N__17829),
            .I(N__17825));
    InMux I__1828 (
            .O(N__17828),
            .I(N__17822));
    LocalMux I__1827 (
            .O(N__17825),
            .I(N__17819));
    LocalMux I__1826 (
            .O(N__17822),
            .I(N__17814));
    Span4Mux_h I__1825 (
            .O(N__17819),
            .I(N__17811));
    InMux I__1824 (
            .O(N__17818),
            .I(N__17806));
    InMux I__1823 (
            .O(N__17817),
            .I(N__17806));
    Odrv4 I__1822 (
            .O(N__17814),
            .I(data_out_frame2_16_6));
    Odrv4 I__1821 (
            .O(N__17811),
            .I(data_out_frame2_16_6));
    LocalMux I__1820 (
            .O(N__17806),
            .I(data_out_frame2_16_6));
    InMux I__1819 (
            .O(N__17799),
            .I(N__17796));
    LocalMux I__1818 (
            .O(N__17796),
            .I(\c0.n18112 ));
    CascadeMux I__1817 (
            .O(N__17793),
            .I(N__17789));
    InMux I__1816 (
            .O(N__17792),
            .I(N__17784));
    InMux I__1815 (
            .O(N__17789),
            .I(N__17784));
    LocalMux I__1814 (
            .O(N__17784),
            .I(data_out_frame2_17_6));
    InMux I__1813 (
            .O(N__17781),
            .I(N__17778));
    LocalMux I__1812 (
            .O(N__17778),
            .I(N__17775));
    Span4Mux_v I__1811 (
            .O(N__17775),
            .I(N__17772));
    Odrv4 I__1810 (
            .O(N__17772),
            .I(\c0.data_out_frame2_20_6 ));
    CascadeMux I__1809 (
            .O(N__17769),
            .I(\c0.n18115_cascade_ ));
    CascadeMux I__1808 (
            .O(N__17766),
            .I(N__17763));
    InMux I__1807 (
            .O(N__17763),
            .I(N__17760));
    LocalMux I__1806 (
            .O(N__17760),
            .I(\c0.n22_adj_2364 ));
    InMux I__1805 (
            .O(N__17757),
            .I(N__17753));
    InMux I__1804 (
            .O(N__17756),
            .I(N__17750));
    LocalMux I__1803 (
            .O(N__17753),
            .I(data_out_frame2_18_6));
    LocalMux I__1802 (
            .O(N__17750),
            .I(data_out_frame2_18_6));
    InMux I__1801 (
            .O(N__17745),
            .I(N__17742));
    LocalMux I__1800 (
            .O(N__17742),
            .I(\c0.n18031 ));
    CascadeMux I__1799 (
            .O(N__17739),
            .I(N__17736));
    InMux I__1798 (
            .O(N__17736),
            .I(N__17733));
    LocalMux I__1797 (
            .O(N__17733),
            .I(N__17730));
    Span4Mux_s3_h I__1796 (
            .O(N__17730),
            .I(N__17727));
    Odrv4 I__1795 (
            .O(N__17727),
            .I(\c0.n10548 ));
    SRMux I__1794 (
            .O(N__17724),
            .I(N__17721));
    LocalMux I__1793 (
            .O(N__17721),
            .I(\c0.n3_adj_2278 ));
    SRMux I__1792 (
            .O(N__17718),
            .I(N__17715));
    LocalMux I__1791 (
            .O(N__17715),
            .I(N__17712));
    Odrv4 I__1790 (
            .O(N__17712),
            .I(\c0.n3_adj_2266 ));
    CascadeMux I__1789 (
            .O(N__17709),
            .I(N__17706));
    InMux I__1788 (
            .O(N__17706),
            .I(N__17703));
    LocalMux I__1787 (
            .O(N__17703),
            .I(N__17700));
    Span4Mux_h I__1786 (
            .O(N__17700),
            .I(N__17697));
    Odrv4 I__1785 (
            .O(N__17697),
            .I(\c0.data_out_frame2_19_6 ));
    IoInMux I__1784 (
            .O(N__17694),
            .I(N__17691));
    LocalMux I__1783 (
            .O(N__17691),
            .I(N__17688));
    Span4Mux_s2_h I__1782 (
            .O(N__17688),
            .I(N__17685));
    Odrv4 I__1781 (
            .O(N__17685),
            .I(tx2_enable));
    SRMux I__1780 (
            .O(N__17682),
            .I(N__17679));
    LocalMux I__1779 (
            .O(N__17679),
            .I(N__17676));
    Odrv4 I__1778 (
            .O(N__17676),
            .I(\c0.n3_adj_2232 ));
    CascadeMux I__1777 (
            .O(N__17673),
            .I(N__17667));
    InMux I__1776 (
            .O(N__17672),
            .I(N__17664));
    InMux I__1775 (
            .O(N__17671),
            .I(N__17660));
    InMux I__1774 (
            .O(N__17670),
            .I(N__17657));
    InMux I__1773 (
            .O(N__17667),
            .I(N__17654));
    LocalMux I__1772 (
            .O(N__17664),
            .I(N__17651));
    InMux I__1771 (
            .O(N__17663),
            .I(N__17648));
    LocalMux I__1770 (
            .O(N__17660),
            .I(N__17645));
    LocalMux I__1769 (
            .O(N__17657),
            .I(N__17640));
    LocalMux I__1768 (
            .O(N__17654),
            .I(N__17640));
    Span4Mux_h I__1767 (
            .O(N__17651),
            .I(N__17637));
    LocalMux I__1766 (
            .O(N__17648),
            .I(data_out_frame2_9_1));
    Odrv4 I__1765 (
            .O(N__17645),
            .I(data_out_frame2_9_1));
    Odrv12 I__1764 (
            .O(N__17640),
            .I(data_out_frame2_9_1));
    Odrv4 I__1763 (
            .O(N__17637),
            .I(data_out_frame2_9_1));
    InMux I__1762 (
            .O(N__17628),
            .I(N__17625));
    LocalMux I__1761 (
            .O(N__17625),
            .I(N__17621));
    InMux I__1760 (
            .O(N__17624),
            .I(N__17618));
    Odrv4 I__1759 (
            .O(N__17621),
            .I(\c0.n10346 ));
    LocalMux I__1758 (
            .O(N__17618),
            .I(\c0.n10346 ));
    InMux I__1757 (
            .O(N__17613),
            .I(N__17610));
    LocalMux I__1756 (
            .O(N__17610),
            .I(N__17606));
    InMux I__1755 (
            .O(N__17609),
            .I(N__17603));
    Odrv12 I__1754 (
            .O(N__17606),
            .I(\c0.n17231 ));
    LocalMux I__1753 (
            .O(N__17603),
            .I(\c0.n17231 ));
    InMux I__1752 (
            .O(N__17598),
            .I(N__17595));
    LocalMux I__1751 (
            .O(N__17595),
            .I(N__17592));
    Odrv4 I__1750 (
            .O(N__17592),
            .I(\c0.n18076 ));
    InMux I__1749 (
            .O(N__17589),
            .I(N__17584));
    InMux I__1748 (
            .O(N__17588),
            .I(N__17581));
    InMux I__1747 (
            .O(N__17587),
            .I(N__17578));
    LocalMux I__1746 (
            .O(N__17584),
            .I(N__17571));
    LocalMux I__1745 (
            .O(N__17581),
            .I(N__17571));
    LocalMux I__1744 (
            .O(N__17578),
            .I(N__17568));
    InMux I__1743 (
            .O(N__17577),
            .I(N__17563));
    InMux I__1742 (
            .O(N__17576),
            .I(N__17563));
    Odrv4 I__1741 (
            .O(N__17571),
            .I(data_out_frame2_9_5));
    Odrv4 I__1740 (
            .O(N__17568),
            .I(data_out_frame2_9_5));
    LocalMux I__1739 (
            .O(N__17563),
            .I(data_out_frame2_9_5));
    InMux I__1738 (
            .O(N__17556),
            .I(N__17553));
    LocalMux I__1737 (
            .O(N__17553),
            .I(N__17550));
    Span4Mux_s2_h I__1736 (
            .O(N__17550),
            .I(N__17547));
    Span4Mux_v I__1735 (
            .O(N__17547),
            .I(N__17544));
    Odrv4 I__1734 (
            .O(N__17544),
            .I(\c0.n18109 ));
    InMux I__1733 (
            .O(N__17541),
            .I(N__17537));
    InMux I__1732 (
            .O(N__17540),
            .I(N__17534));
    LocalMux I__1731 (
            .O(N__17537),
            .I(N__17530));
    LocalMux I__1730 (
            .O(N__17534),
            .I(N__17526));
    InMux I__1729 (
            .O(N__17533),
            .I(N__17523));
    Span4Mux_v I__1728 (
            .O(N__17530),
            .I(N__17520));
    InMux I__1727 (
            .O(N__17529),
            .I(N__17517));
    Span4Mux_s1_h I__1726 (
            .O(N__17526),
            .I(N__17514));
    LocalMux I__1725 (
            .O(N__17523),
            .I(data_out_frame2_6_3));
    Odrv4 I__1724 (
            .O(N__17520),
            .I(data_out_frame2_6_3));
    LocalMux I__1723 (
            .O(N__17517),
            .I(data_out_frame2_6_3));
    Odrv4 I__1722 (
            .O(N__17514),
            .I(data_out_frame2_6_3));
    CascadeMux I__1721 (
            .O(N__17505),
            .I(\c0.n10334_cascade_ ));
    InMux I__1720 (
            .O(N__17502),
            .I(N__17498));
    InMux I__1719 (
            .O(N__17501),
            .I(N__17495));
    LocalMux I__1718 (
            .O(N__17498),
            .I(\c0.n10533 ));
    LocalMux I__1717 (
            .O(N__17495),
            .I(\c0.n10533 ));
    InMux I__1716 (
            .O(N__17490),
            .I(N__17487));
    LocalMux I__1715 (
            .O(N__17487),
            .I(\c0.n10_adj_2297 ));
    CascadeMux I__1714 (
            .O(N__17484),
            .I(\c0.n14_adj_2296_cascade_ ));
    InMux I__1713 (
            .O(N__17481),
            .I(N__17478));
    LocalMux I__1712 (
            .O(N__17478),
            .I(N__17474));
    InMux I__1711 (
            .O(N__17477),
            .I(N__17471));
    Sp12to4 I__1710 (
            .O(N__17474),
            .I(N__17468));
    LocalMux I__1709 (
            .O(N__17471),
            .I(N__17465));
    Odrv12 I__1708 (
            .O(N__17468),
            .I(\c0.n17267 ));
    Odrv12 I__1707 (
            .O(N__17465),
            .I(\c0.n17267 ));
    InMux I__1706 (
            .O(N__17460),
            .I(N__17457));
    LocalMux I__1705 (
            .O(N__17457),
            .I(N__17453));
    InMux I__1704 (
            .O(N__17456),
            .I(N__17450));
    Span4Mux_v I__1703 (
            .O(N__17453),
            .I(N__17447));
    LocalMux I__1702 (
            .O(N__17450),
            .I(N__17444));
    Span4Mux_v I__1701 (
            .O(N__17447),
            .I(N__17438));
    Span4Mux_v I__1700 (
            .O(N__17444),
            .I(N__17435));
    InMux I__1699 (
            .O(N__17443),
            .I(N__17428));
    InMux I__1698 (
            .O(N__17442),
            .I(N__17428));
    InMux I__1697 (
            .O(N__17441),
            .I(N__17428));
    Odrv4 I__1696 (
            .O(N__17438),
            .I(data_out_frame2_13_2));
    Odrv4 I__1695 (
            .O(N__17435),
            .I(data_out_frame2_13_2));
    LocalMux I__1694 (
            .O(N__17428),
            .I(data_out_frame2_13_2));
    InMux I__1693 (
            .O(N__17421),
            .I(N__17418));
    LocalMux I__1692 (
            .O(N__17418),
            .I(N__17415));
    Span4Mux_s2_h I__1691 (
            .O(N__17415),
            .I(N__17411));
    InMux I__1690 (
            .O(N__17414),
            .I(N__17408));
    Odrv4 I__1689 (
            .O(N__17411),
            .I(\c0.n17309 ));
    LocalMux I__1688 (
            .O(N__17408),
            .I(\c0.n17309 ));
    InMux I__1687 (
            .O(N__17403),
            .I(N__17399));
    InMux I__1686 (
            .O(N__17402),
            .I(N__17396));
    LocalMux I__1685 (
            .O(N__17399),
            .I(N__17393));
    LocalMux I__1684 (
            .O(N__17396),
            .I(\c0.n17291 ));
    Odrv4 I__1683 (
            .O(N__17393),
            .I(\c0.n17291 ));
    InMux I__1682 (
            .O(N__17388),
            .I(N__17385));
    LocalMux I__1681 (
            .O(N__17385),
            .I(N__17382));
    Span4Mux_v I__1680 (
            .O(N__17382),
            .I(N__17378));
    InMux I__1679 (
            .O(N__17381),
            .I(N__17375));
    Odrv4 I__1678 (
            .O(N__17378),
            .I(\c0.n17303 ));
    LocalMux I__1677 (
            .O(N__17375),
            .I(\c0.n17303 ));
    InMux I__1676 (
            .O(N__17370),
            .I(N__17367));
    LocalMux I__1675 (
            .O(N__17367),
            .I(\c0.n25 ));
    CascadeMux I__1674 (
            .O(N__17364),
            .I(\c0.n28_adj_2200_cascade_ ));
    InMux I__1673 (
            .O(N__17361),
            .I(N__17358));
    LocalMux I__1672 (
            .O(N__17358),
            .I(\c0.n27_adj_2204 ));
    CascadeMux I__1671 (
            .O(N__17355),
            .I(\c0.n10223_cascade_ ));
    InMux I__1670 (
            .O(N__17352),
            .I(N__17349));
    LocalMux I__1669 (
            .O(N__17349),
            .I(\c0.n6_adj_2318 ));
    CascadeMux I__1668 (
            .O(N__17346),
            .I(N__17343));
    InMux I__1667 (
            .O(N__17343),
            .I(N__17340));
    LocalMux I__1666 (
            .O(N__17340),
            .I(N__17337));
    Span4Mux_s2_h I__1665 (
            .O(N__17337),
            .I(N__17334));
    Odrv4 I__1664 (
            .O(N__17334),
            .I(\c0.n17569 ));
    InMux I__1663 (
            .O(N__17331),
            .I(N__17328));
    LocalMux I__1662 (
            .O(N__17328),
            .I(N__17324));
    InMux I__1661 (
            .O(N__17327),
            .I(N__17321));
    Span4Mux_v I__1660 (
            .O(N__17324),
            .I(N__17318));
    LocalMux I__1659 (
            .O(N__17321),
            .I(data_out_frame2_17_5));
    Odrv4 I__1658 (
            .O(N__17318),
            .I(data_out_frame2_17_5));
    CascadeMux I__1657 (
            .O(N__17313),
            .I(N__17309));
    InMux I__1656 (
            .O(N__17312),
            .I(N__17306));
    InMux I__1655 (
            .O(N__17309),
            .I(N__17303));
    LocalMux I__1654 (
            .O(N__17306),
            .I(N__17298));
    LocalMux I__1653 (
            .O(N__17303),
            .I(N__17298));
    Odrv4 I__1652 (
            .O(N__17298),
            .I(\c0.n17138 ));
    CascadeMux I__1651 (
            .O(N__17295),
            .I(\c0.n6_adj_2228_cascade_ ));
    InMux I__1650 (
            .O(N__17292),
            .I(N__17289));
    LocalMux I__1649 (
            .O(N__17289),
            .I(N__17286));
    Span4Mux_s3_h I__1648 (
            .O(N__17286),
            .I(N__17282));
    InMux I__1647 (
            .O(N__17285),
            .I(N__17279));
    Odrv4 I__1646 (
            .O(N__17282),
            .I(\c0.n17312 ));
    LocalMux I__1645 (
            .O(N__17279),
            .I(\c0.n17312 ));
    InMux I__1644 (
            .O(N__17274),
            .I(N__17266));
    InMux I__1643 (
            .O(N__17273),
            .I(N__17266));
    InMux I__1642 (
            .O(N__17272),
            .I(N__17262));
    InMux I__1641 (
            .O(N__17271),
            .I(N__17259));
    LocalMux I__1640 (
            .O(N__17266),
            .I(N__17256));
    InMux I__1639 (
            .O(N__17265),
            .I(N__17253));
    LocalMux I__1638 (
            .O(N__17262),
            .I(N__17250));
    LocalMux I__1637 (
            .O(N__17259),
            .I(data_out_frame2_14_3));
    Odrv4 I__1636 (
            .O(N__17256),
            .I(data_out_frame2_14_3));
    LocalMux I__1635 (
            .O(N__17253),
            .I(data_out_frame2_14_3));
    Odrv4 I__1634 (
            .O(N__17250),
            .I(data_out_frame2_14_3));
    CascadeMux I__1633 (
            .O(N__17241),
            .I(\c0.n33_cascade_ ));
    CascadeMux I__1632 (
            .O(N__17238),
            .I(N__17235));
    InMux I__1631 (
            .O(N__17235),
            .I(N__17232));
    LocalMux I__1630 (
            .O(N__17232),
            .I(N__17229));
    Odrv4 I__1629 (
            .O(N__17229),
            .I(\c0.data_out_frame2_19_7 ));
    InMux I__1628 (
            .O(N__17226),
            .I(N__17223));
    LocalMux I__1627 (
            .O(N__17223),
            .I(\c0.n30_adj_2218 ));
    CascadeMux I__1626 (
            .O(N__17220),
            .I(\c0.n17300_cascade_ ));
    InMux I__1625 (
            .O(N__17217),
            .I(N__17214));
    LocalMux I__1624 (
            .O(N__17214),
            .I(\c0.n34 ));
    CascadeMux I__1623 (
            .O(N__17211),
            .I(N__17208));
    InMux I__1622 (
            .O(N__17208),
            .I(N__17205));
    LocalMux I__1621 (
            .O(N__17205),
            .I(N__17202));
    Odrv12 I__1620 (
            .O(N__17202),
            .I(\c0.n17237 ));
    CascadeMux I__1619 (
            .O(N__17199),
            .I(N__17196));
    InMux I__1618 (
            .O(N__17196),
            .I(N__17193));
    LocalMux I__1617 (
            .O(N__17193),
            .I(N__17190));
    Span4Mux_v I__1616 (
            .O(N__17190),
            .I(N__17187));
    Odrv4 I__1615 (
            .O(N__17187),
            .I(\c0.n10440 ));
    InMux I__1614 (
            .O(N__17184),
            .I(N__17181));
    LocalMux I__1613 (
            .O(N__17181),
            .I(\c0.n6_adj_2215 ));
    InMux I__1612 (
            .O(N__17178),
            .I(N__17175));
    LocalMux I__1611 (
            .O(N__17175),
            .I(\c0.n17219 ));
    InMux I__1610 (
            .O(N__17172),
            .I(N__17169));
    LocalMux I__1609 (
            .O(N__17169),
            .I(N__17166));
    Odrv4 I__1608 (
            .O(N__17166),
            .I(\c0.n17141 ));
    CascadeMux I__1607 (
            .O(N__17163),
            .I(\c0.n17219_cascade_ ));
    CascadeMux I__1606 (
            .O(N__17160),
            .I(\c0.n17_cascade_ ));
    InMux I__1605 (
            .O(N__17157),
            .I(N__17153));
    InMux I__1604 (
            .O(N__17156),
            .I(N__17150));
    LocalMux I__1603 (
            .O(N__17153),
            .I(N__17147));
    LocalMux I__1602 (
            .O(N__17150),
            .I(N__17144));
    Odrv4 I__1601 (
            .O(N__17147),
            .I(\c0.n17228 ));
    Odrv4 I__1600 (
            .O(N__17144),
            .I(\c0.n17228 ));
    CascadeMux I__1599 (
            .O(N__17139),
            .I(\c0.n17246_cascade_ ));
    InMux I__1598 (
            .O(N__17136),
            .I(N__17133));
    LocalMux I__1597 (
            .O(N__17133),
            .I(N__17130));
    Span4Mux_h I__1596 (
            .O(N__17130),
            .I(N__17127));
    Odrv4 I__1595 (
            .O(N__17127),
            .I(\c0.n17187 ));
    CascadeMux I__1594 (
            .O(N__17124),
            .I(\c0.n18238_cascade_ ));
    InMux I__1593 (
            .O(N__17121),
            .I(N__17118));
    LocalMux I__1592 (
            .O(N__17118),
            .I(\c0.n18241 ));
    InMux I__1591 (
            .O(N__17115),
            .I(N__17112));
    LocalMux I__1590 (
            .O(N__17112),
            .I(N__17109));
    Span4Mux_h I__1589 (
            .O(N__17109),
            .I(N__17106));
    Span4Mux_v I__1588 (
            .O(N__17106),
            .I(N__17100));
    InMux I__1587 (
            .O(N__17105),
            .I(N__17097));
    InMux I__1586 (
            .O(N__17104),
            .I(N__17092));
    InMux I__1585 (
            .O(N__17103),
            .I(N__17092));
    Odrv4 I__1584 (
            .O(N__17100),
            .I(data_out_frame2_7_7));
    LocalMux I__1583 (
            .O(N__17097),
            .I(data_out_frame2_7_7));
    LocalMux I__1582 (
            .O(N__17092),
            .I(data_out_frame2_7_7));
    InMux I__1581 (
            .O(N__17085),
            .I(N__17082));
    LocalMux I__1580 (
            .O(N__17082),
            .I(N__17079));
    Odrv4 I__1579 (
            .O(N__17079),
            .I(\c0.n5_adj_2137 ));
    InMux I__1578 (
            .O(N__17076),
            .I(N__17073));
    LocalMux I__1577 (
            .O(N__17073),
            .I(\c0.n18154 ));
    CascadeMux I__1576 (
            .O(N__17070),
            .I(\c0.n18130_cascade_ ));
    InMux I__1575 (
            .O(N__17067),
            .I(N__17064));
    LocalMux I__1574 (
            .O(N__17064),
            .I(N__17061));
    Span4Mux_v I__1573 (
            .O(N__17061),
            .I(N__17058));
    Span4Mux_v I__1572 (
            .O(N__17058),
            .I(N__17055));
    Odrv4 I__1571 (
            .O(N__17055),
            .I(\c0.data_out_frame2_20_7 ));
    CascadeMux I__1570 (
            .O(N__17052),
            .I(\c0.n18133_cascade_ ));
    CascadeMux I__1569 (
            .O(N__17049),
            .I(N__17046));
    InMux I__1568 (
            .O(N__17046),
            .I(N__17043));
    LocalMux I__1567 (
            .O(N__17043),
            .I(N__17040));
    Odrv4 I__1566 (
            .O(N__17040),
            .I(\c0.n22_adj_2363 ));
    InMux I__1565 (
            .O(N__17037),
            .I(N__17034));
    LocalMux I__1564 (
            .O(N__17034),
            .I(N__17031));
    Span4Mux_h I__1563 (
            .O(N__17031),
            .I(N__17028));
    Span4Mux_s1_h I__1562 (
            .O(N__17028),
            .I(N__17025));
    Span4Mux_h I__1561 (
            .O(N__17025),
            .I(N__17022));
    Odrv4 I__1560 (
            .O(N__17022),
            .I(\c0.n18028 ));
    CascadeMux I__1559 (
            .O(N__17019),
            .I(\c0.n18040_cascade_ ));
    CascadeMux I__1558 (
            .O(N__17016),
            .I(\c0.n18010_cascade_ ));
    CascadeMux I__1557 (
            .O(N__17013),
            .I(\c0.n18013_cascade_ ));
    CascadeMux I__1556 (
            .O(N__17010),
            .I(N__17007));
    InMux I__1555 (
            .O(N__17007),
            .I(N__17004));
    LocalMux I__1554 (
            .O(N__17004),
            .I(\c0.n22_adj_2375 ));
    InMux I__1553 (
            .O(N__17001),
            .I(N__16998));
    LocalMux I__1552 (
            .O(N__16998),
            .I(N__16995));
    Odrv4 I__1551 (
            .O(N__16995),
            .I(\c0.n18025 ));
    InMux I__1550 (
            .O(N__16992),
            .I(N__16989));
    LocalMux I__1549 (
            .O(N__16989),
            .I(N__16986));
    Odrv12 I__1548 (
            .O(N__16986),
            .I(\c0.n10530 ));
    CascadeMux I__1547 (
            .O(N__16983),
            .I(\c0.n10530_cascade_ ));
    InMux I__1546 (
            .O(N__16980),
            .I(N__16976));
    InMux I__1545 (
            .O(N__16979),
            .I(N__16973));
    LocalMux I__1544 (
            .O(N__16976),
            .I(N__16970));
    LocalMux I__1543 (
            .O(N__16973),
            .I(N__16967));
    Odrv4 I__1542 (
            .O(N__16970),
            .I(\c0.n10371 ));
    Odrv4 I__1541 (
            .O(N__16967),
            .I(\c0.n10371 ));
    InMux I__1540 (
            .O(N__16962),
            .I(N__16956));
    InMux I__1539 (
            .O(N__16961),
            .I(N__16953));
    InMux I__1538 (
            .O(N__16960),
            .I(N__16948));
    InMux I__1537 (
            .O(N__16959),
            .I(N__16948));
    LocalMux I__1536 (
            .O(N__16956),
            .I(N__16945));
    LocalMux I__1535 (
            .O(N__16953),
            .I(data_out_frame2_7_0));
    LocalMux I__1534 (
            .O(N__16948),
            .I(data_out_frame2_7_0));
    Odrv4 I__1533 (
            .O(N__16945),
            .I(data_out_frame2_7_0));
    CascadeMux I__1532 (
            .O(N__16938),
            .I(N__16934));
    InMux I__1531 (
            .O(N__16937),
            .I(N__16927));
    InMux I__1530 (
            .O(N__16934),
            .I(N__16927));
    InMux I__1529 (
            .O(N__16933),
            .I(N__16922));
    InMux I__1528 (
            .O(N__16932),
            .I(N__16922));
    LocalMux I__1527 (
            .O(N__16927),
            .I(N__16919));
    LocalMux I__1526 (
            .O(N__16922),
            .I(data_out_frame2_6_0));
    Odrv4 I__1525 (
            .O(N__16919),
            .I(data_out_frame2_6_0));
    CascadeMux I__1524 (
            .O(N__16914),
            .I(N__16911));
    InMux I__1523 (
            .O(N__16911),
            .I(N__16908));
    LocalMux I__1522 (
            .O(N__16908),
            .I(N__16905));
    Span4Mux_s1_h I__1521 (
            .O(N__16905),
            .I(N__16902));
    Odrv4 I__1520 (
            .O(N__16902),
            .I(\c0.n5_adj_2343 ));
    CascadeMux I__1519 (
            .O(N__16899),
            .I(N__16895));
    InMux I__1518 (
            .O(N__16898),
            .I(N__16892));
    InMux I__1517 (
            .O(N__16895),
            .I(N__16887));
    LocalMux I__1516 (
            .O(N__16892),
            .I(N__16884));
    InMux I__1515 (
            .O(N__16891),
            .I(N__16881));
    InMux I__1514 (
            .O(N__16890),
            .I(N__16878));
    LocalMux I__1513 (
            .O(N__16887),
            .I(N__16871));
    Span4Mux_v I__1512 (
            .O(N__16884),
            .I(N__16871));
    LocalMux I__1511 (
            .O(N__16881),
            .I(N__16871));
    LocalMux I__1510 (
            .O(N__16878),
            .I(data_out_frame2_15_5));
    Odrv4 I__1509 (
            .O(N__16871),
            .I(data_out_frame2_15_5));
    CascadeMux I__1508 (
            .O(N__16866),
            .I(\c0.n18100_cascade_ ));
    CascadeMux I__1507 (
            .O(N__16863),
            .I(N__16860));
    InMux I__1506 (
            .O(N__16860),
            .I(N__16857));
    LocalMux I__1505 (
            .O(N__16857),
            .I(N__16854));
    Span12Mux_s1_h I__1504 (
            .O(N__16854),
            .I(N__16851));
    Odrv12 I__1503 (
            .O(N__16851),
            .I(\c0.n18103 ));
    CascadeMux I__1502 (
            .O(N__16848),
            .I(\c0.n10520_cascade_ ));
    InMux I__1501 (
            .O(N__16845),
            .I(N__16842));
    LocalMux I__1500 (
            .O(N__16842),
            .I(N__16838));
    InMux I__1499 (
            .O(N__16841),
            .I(N__16835));
    Odrv12 I__1498 (
            .O(N__16838),
            .I(\c0.n10349 ));
    LocalMux I__1497 (
            .O(N__16835),
            .I(\c0.n10349 ));
    InMux I__1496 (
            .O(N__16830),
            .I(N__16827));
    LocalMux I__1495 (
            .O(N__16827),
            .I(N__16824));
    Odrv12 I__1494 (
            .O(N__16824),
            .I(\c0.n10462 ));
    InMux I__1493 (
            .O(N__16821),
            .I(N__16818));
    LocalMux I__1492 (
            .O(N__16818),
            .I(N__16815));
    Odrv12 I__1491 (
            .O(N__16815),
            .I(\c0.n15_adj_2312 ));
    CascadeMux I__1490 (
            .O(N__16812),
            .I(N__16808));
    InMux I__1489 (
            .O(N__16811),
            .I(N__16805));
    InMux I__1488 (
            .O(N__16808),
            .I(N__16802));
    LocalMux I__1487 (
            .O(N__16805),
            .I(N__16799));
    LocalMux I__1486 (
            .O(N__16802),
            .I(N__16796));
    Odrv4 I__1485 (
            .O(N__16799),
            .I(\c0.n17285 ));
    Odrv4 I__1484 (
            .O(N__16796),
            .I(\c0.n17285 ));
    InMux I__1483 (
            .O(N__16791),
            .I(N__16788));
    LocalMux I__1482 (
            .O(N__16788),
            .I(\c0.n18136 ));
    CascadeMux I__1481 (
            .O(N__16785),
            .I(N__16782));
    InMux I__1480 (
            .O(N__16782),
            .I(N__16779));
    LocalMux I__1479 (
            .O(N__16779),
            .I(N__16776));
    Span4Mux_v I__1478 (
            .O(N__16776),
            .I(N__16773));
    Odrv4 I__1477 (
            .O(N__16773),
            .I(\c0.data_out_frame2_19_2 ));
    InMux I__1476 (
            .O(N__16770),
            .I(N__16767));
    LocalMux I__1475 (
            .O(N__16767),
            .I(\c0.n17135 ));
    CascadeMux I__1474 (
            .O(N__16764),
            .I(\c0.n17092_cascade_ ));
    CascadeMux I__1473 (
            .O(N__16761),
            .I(\c0.n17_adj_2294_cascade_ ));
    CascadeMux I__1472 (
            .O(N__16758),
            .I(N__16755));
    InMux I__1471 (
            .O(N__16755),
            .I(N__16752));
    LocalMux I__1470 (
            .O(N__16752),
            .I(N__16749));
    Odrv12 I__1469 (
            .O(N__16749),
            .I(\c0.data_out_frame2_19_4 ));
    InMux I__1468 (
            .O(N__16746),
            .I(N__16743));
    LocalMux I__1467 (
            .O(N__16743),
            .I(\c0.n12 ));
    InMux I__1466 (
            .O(N__16740),
            .I(N__16735));
    InMux I__1465 (
            .O(N__16739),
            .I(N__16730));
    InMux I__1464 (
            .O(N__16738),
            .I(N__16730));
    LocalMux I__1463 (
            .O(N__16735),
            .I(N__16727));
    LocalMux I__1462 (
            .O(N__16730),
            .I(data_out_frame2_14_0));
    Odrv12 I__1461 (
            .O(N__16727),
            .I(data_out_frame2_14_0));
    CascadeMux I__1460 (
            .O(N__16722),
            .I(\c0.n17237_cascade_ ));
    InMux I__1459 (
            .O(N__16719),
            .I(N__16716));
    LocalMux I__1458 (
            .O(N__16716),
            .I(\c0.n16_adj_2293 ));
    InMux I__1457 (
            .O(N__16713),
            .I(N__16710));
    LocalMux I__1456 (
            .O(N__16710),
            .I(N__16707));
    Span4Mux_h I__1455 (
            .O(N__16707),
            .I(N__16704));
    Odrv4 I__1454 (
            .O(N__16704),
            .I(\c0.data_out_frame2_20_4 ));
    CascadeMux I__1453 (
            .O(N__16701),
            .I(\c0.n18277_cascade_ ));
    InMux I__1452 (
            .O(N__16698),
            .I(N__16695));
    LocalMux I__1451 (
            .O(N__16695),
            .I(\c0.n22_adj_2367 ));
    InMux I__1450 (
            .O(N__16692),
            .I(N__16689));
    LocalMux I__1449 (
            .O(N__16689),
            .I(\c0.n18034 ));
    InMux I__1448 (
            .O(N__16686),
            .I(N__16683));
    LocalMux I__1447 (
            .O(N__16683),
            .I(N__16679));
    CascadeMux I__1446 (
            .O(N__16682),
            .I(N__16676));
    Span4Mux_h I__1445 (
            .O(N__16679),
            .I(N__16673));
    InMux I__1444 (
            .O(N__16676),
            .I(N__16670));
    Odrv4 I__1443 (
            .O(N__16673),
            .I(\c0.n17225 ));
    LocalMux I__1442 (
            .O(N__16670),
            .I(\c0.n17225 ));
    CascadeMux I__1441 (
            .O(N__16665),
            .I(\c0.n17135_cascade_ ));
    CascadeMux I__1440 (
            .O(N__16662),
            .I(\c0.n21_cascade_ ));
    InMux I__1439 (
            .O(N__16659),
            .I(N__16656));
    LocalMux I__1438 (
            .O(N__16656),
            .I(\c0.n20_adj_2223 ));
    InMux I__1437 (
            .O(N__16653),
            .I(N__16650));
    LocalMux I__1436 (
            .O(N__16650),
            .I(\c0.n19_adj_2224 ));
    CascadeMux I__1435 (
            .O(N__16647),
            .I(\c0.n14_adj_2308_cascade_ ));
    InMux I__1434 (
            .O(N__16644),
            .I(N__16641));
    LocalMux I__1433 (
            .O(N__16641),
            .I(\c0.n18022 ));
    CascadeMux I__1432 (
            .O(N__16638),
            .I(\c0.n5_adj_2353_cascade_ ));
    InMux I__1431 (
            .O(N__16635),
            .I(N__16632));
    LocalMux I__1430 (
            .O(N__16632),
            .I(N__16629));
    Odrv4 I__1429 (
            .O(N__16629),
            .I(\c0.n6 ));
    InMux I__1428 (
            .O(N__16626),
            .I(N__16623));
    LocalMux I__1427 (
            .O(N__16623),
            .I(N__16620));
    Odrv4 I__1426 (
            .O(N__16620),
            .I(\c0.n6_adj_2138 ));
    InMux I__1425 (
            .O(N__16617),
            .I(N__16614));
    LocalMux I__1424 (
            .O(N__16614),
            .I(N__16611));
    Span4Mux_h I__1423 (
            .O(N__16611),
            .I(N__16608));
    Span4Mux_v I__1422 (
            .O(N__16608),
            .I(N__16605));
    Odrv4 I__1421 (
            .O(N__16605),
            .I(\c0.n17440 ));
    CascadeMux I__1420 (
            .O(N__16602),
            .I(\c0.n18037_cascade_ ));
    CascadeMux I__1419 (
            .O(N__16599),
            .I(\c0.n18274_cascade_ ));
    CascadeMux I__1418 (
            .O(N__16596),
            .I(\c0.n5_adj_2315_cascade_ ));
    InMux I__1417 (
            .O(N__16593),
            .I(N__16586));
    InMux I__1416 (
            .O(N__16592),
            .I(N__16586));
    InMux I__1415 (
            .O(N__16591),
            .I(N__16583));
    LocalMux I__1414 (
            .O(N__16586),
            .I(data_out_frame2_13_7));
    LocalMux I__1413 (
            .O(N__16583),
            .I(data_out_frame2_13_7));
    InMux I__1412 (
            .O(N__16578),
            .I(N__16574));
    InMux I__1411 (
            .O(N__16577),
            .I(N__16571));
    LocalMux I__1410 (
            .O(N__16574),
            .I(N__16568));
    LocalMux I__1409 (
            .O(N__16571),
            .I(data_out_frame2_18_5));
    Odrv4 I__1408 (
            .O(N__16568),
            .I(data_out_frame2_18_5));
    CascadeMux I__1407 (
            .O(N__16563),
            .I(\c0.n24_cascade_ ));
    InMux I__1406 (
            .O(N__16560),
            .I(N__16557));
    LocalMux I__1405 (
            .O(N__16557),
            .I(\c0.n22 ));
    InMux I__1404 (
            .O(N__16554),
            .I(N__16551));
    LocalMux I__1403 (
            .O(N__16551),
            .I(\c0.n17174 ));
    CascadeMux I__1402 (
            .O(N__16548),
            .I(\c0.n17174_cascade_ ));
    CascadeMux I__1401 (
            .O(N__16545),
            .I(\c0.n10356_cascade_ ));
    CascadeMux I__1400 (
            .O(N__16542),
            .I(N__16539));
    InMux I__1399 (
            .O(N__16539),
            .I(N__16536));
    LocalMux I__1398 (
            .O(N__16536),
            .I(N__16533));
    Odrv12 I__1397 (
            .O(N__16533),
            .I(\c0.n18139 ));
    InMux I__1396 (
            .O(N__16530),
            .I(N__16527));
    LocalMux I__1395 (
            .O(N__16527),
            .I(N__16524));
    Odrv4 I__1394 (
            .O(N__16524),
            .I(\c0.n14 ));
    CascadeMux I__1393 (
            .O(N__16521),
            .I(\c0.n15_cascade_ ));
    InMux I__1392 (
            .O(N__16518),
            .I(N__16515));
    LocalMux I__1391 (
            .O(N__16515),
            .I(\c0.data_out_frame2_20_5 ));
    CascadeMux I__1390 (
            .O(N__16512),
            .I(\c0.n17306_cascade_ ));
    CascadeMux I__1389 (
            .O(N__16509),
            .I(\c0.n18094_cascade_ ));
    CascadeMux I__1388 (
            .O(N__16506),
            .I(\c0.n18097_cascade_ ));
    CascadeMux I__1387 (
            .O(N__16503),
            .I(\c0.n18262_cascade_ ));
    InMux I__1386 (
            .O(N__16500),
            .I(N__16497));
    LocalMux I__1385 (
            .O(N__16497),
            .I(\c0.n22_adj_2365 ));
    CascadeMux I__1384 (
            .O(N__16494),
            .I(\c0.n18265_cascade_ ));
    CascadeMux I__1383 (
            .O(N__16491),
            .I(\c0.n10468_cascade_ ));
    CascadeMux I__1382 (
            .O(N__16488),
            .I(\c0.n17610_cascade_ ));
    InMux I__1381 (
            .O(N__16485),
            .I(N__16482));
    LocalMux I__1380 (
            .O(N__16482),
            .I(\c0.n18214 ));
    InMux I__1379 (
            .O(N__16479),
            .I(N__16476));
    LocalMux I__1378 (
            .O(N__16476),
            .I(\c0.n18217 ));
    IoInMux I__1377 (
            .O(N__16473),
            .I(N__16470));
    LocalMux I__1376 (
            .O(N__16470),
            .I(N__16467));
    IoSpan4Mux I__1375 (
            .O(N__16467),
            .I(N__16464));
    IoSpan4Mux I__1374 (
            .O(N__16464),
            .I(N__16461));
    IoSpan4Mux I__1373 (
            .O(N__16461),
            .I(N__16458));
    Odrv4 I__1372 (
            .O(N__16458),
            .I(CLK_pad_gb_input));
    defparam IN_MUX_bfv_10_25_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_25_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_25_0_));
    defparam IN_MUX_bfv_10_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_26_0_ (
            .carryinitin(n16017),
            .carryinitout(bfn_10_26_0_));
    defparam IN_MUX_bfv_10_27_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_27_0_ (
            .carryinitin(n16025),
            .carryinitout(bfn_10_27_0_));
    defparam IN_MUX_bfv_10_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_28_0_ (
            .carryinitin(n16033),
            .carryinitout(bfn_10_28_0_));
    defparam IN_MUX_bfv_5_23_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_23_0_));
    defparam IN_MUX_bfv_5_24_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_24_0_ (
            .carryinitin(n15986),
            .carryinitout(bfn_5_24_0_));
    defparam IN_MUX_bfv_5_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_25_0_ (
            .carryinitin(n15994),
            .carryinitout(bfn_5_25_0_));
    defparam IN_MUX_bfv_5_26_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_26_0_ (
            .carryinitin(n16002),
            .carryinitout(bfn_5_26_0_));
    defparam IN_MUX_bfv_6_24_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_24_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_24_0_));
    defparam IN_MUX_bfv_6_25_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_25_0_ (
            .carryinitin(\c0.tx2.n16139 ),
            .carryinitout(bfn_6_25_0_));
    defparam IN_MUX_bfv_16_28_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_28_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_28_0_));
    defparam IN_MUX_bfv_16_29_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_29_0_ (
            .carryinitin(\c0.tx.n16124 ),
            .carryinitout(bfn_16_29_0_));
    defparam IN_MUX_bfv_4_32_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_32_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_32_0_));
    defparam IN_MUX_bfv_12_31_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_31_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_31_0_));
    defparam IN_MUX_bfv_12_32_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_32_0_ (
            .carryinitin(\c0.n16073 ),
            .carryinitout(bfn_12_32_0_));
    defparam IN_MUX_bfv_4_27_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_27_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_27_0_));
    defparam IN_MUX_bfv_4_28_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_28_0_ (
            .carryinitin(\c0.n16086 ),
            .carryinitout(bfn_4_28_0_));
    defparam IN_MUX_bfv_4_29_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_29_0_ (
            .carryinitin(\c0.n16094 ),
            .carryinitout(bfn_4_29_0_));
    defparam IN_MUX_bfv_4_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_30_0_ (
            .carryinitin(\c0.n16102 ),
            .carryinitout(bfn_4_30_0_));
    defparam IN_MUX_bfv_9_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_17_0_));
    defparam IN_MUX_bfv_14_30_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_30_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_30_0_));
    defparam IN_MUX_bfv_9_29_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_29_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_29_0_));
    defparam IN_MUX_bfv_9_30_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_30_0_ (
            .carryinitin(n16048),
            .carryinitout(bfn_9_30_0_));
    defparam IN_MUX_bfv_9_31_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_31_0_ (
            .carryinitin(n16056),
            .carryinitout(bfn_9_31_0_));
    defparam IN_MUX_bfv_9_32_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_32_0_ (
            .carryinitin(n16064),
            .carryinitout(bfn_9_32_0_));
    ICE_GB CLK_pad_gb (
            .USERSIGNALTOGLOBALBUFFER(N__16473),
            .GLOBALBUFFEROUTPUT(CLK_c));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_695_LC_1_17_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_695_LC_1_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_695_LC_1_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_695_LC_1_17_1  (
            .in0(N__24937),
            .in1(N__17460),
            .in2(_gnd_net_),
            .in3(N__18732),
            .lcout(\c0.n10440 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18022_bdd_4_lut_LC_1_17_5 .C_ON=1'b0;
    defparam \c0.n18022_bdd_4_lut_LC_1_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.n18022_bdd_4_lut_LC_1_17_5 .LUT_INIT=16'b1101100111001000;
    LogicCell40 \c0.n18022_bdd_4_lut_LC_1_17_5  (
            .in0(N__28699),
            .in1(N__16644),
            .in2(N__17673),
            .in3(N__18086),
            .lcout(\c0.n18025 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15153_3_lut_LC_1_17_6 .C_ON=1'b0;
    defparam \c0.i15153_3_lut_LC_1_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.i15153_3_lut_LC_1_17_6 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \c0.i15153_3_lut_LC_1_17_6  (
            .in0(N__34724),
            .in1(N__28969),
            .in2(_gnd_net_),
            .in3(N__28700),
            .lcout(),
            .ltout(\c0.n17610_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18214_bdd_4_lut_LC_1_17_7 .C_ON=1'b0;
    defparam \c0.n18214_bdd_4_lut_LC_1_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.n18214_bdd_4_lut_LC_1_17_7 .LUT_INIT=16'b1100110010111000;
    LogicCell40 \c0.n18214_bdd_4_lut_LC_1_17_7  (
            .in0(N__16626),
            .in1(N__16485),
            .in2(N__16488),
            .in3(N__32463),
            .lcout(\c0.n18217 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15410_LC_1_18_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15410_LC_1_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15410_LC_1_18_3 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_15410_LC_1_18_3  (
            .in0(N__23412),
            .in1(N__32458),
            .in2(N__16542),
            .in3(N__32171),
            .lcout(\c0.n18214 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i7_LC_1_18_5 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i7_LC_1_18_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i7_LC_1_18_5 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \c0.tx2.r_Tx_Data_i7_LC_1_18_5  (
            .in0(N__16479),
            .in1(N__32459),
            .in2(N__17049),
            .in3(N__32289),
            .lcout(\c0.tx2.r_Tx_Data_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49627),
            .ce(N__24272),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15306_LC_1_19_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15306_LC_1_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15306_LC_1_19_0 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15306_LC_1_19_0  (
            .in0(N__28652),
            .in1(N__16578),
            .in2(N__19677),
            .in3(N__29048),
            .lcout(),
            .ltout(\c0.n18094_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18094_bdd_4_lut_LC_1_19_1 .C_ON=1'b0;
    defparam \c0.n18094_bdd_4_lut_LC_1_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.n18094_bdd_4_lut_LC_1_19_1 .LUT_INIT=16'b1110001111100000;
    LogicCell40 \c0.n18094_bdd_4_lut_LC_1_19_1  (
            .in0(N__17331),
            .in1(N__28653),
            .in2(N__16509),
            .in3(N__20561),
            .lcout(),
            .ltout(\c0.n18097_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_5_i22_4_lut_LC_1_19_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_5_i22_4_lut_LC_1_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_5_i22_4_lut_LC_1_19_2 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_5_i22_4_lut_LC_1_19_2  (
            .in0(N__32172),
            .in1(N__16518),
            .in2(N__16506),
            .in3(N__21210),
            .lcout(\c0.n22_adj_2365 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_LC_1_19_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_LC_1_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_LC_1_19_3 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_LC_1_19_3  (
            .in0(N__17556),
            .in1(N__32460),
            .in2(N__16863),
            .in3(N__32173),
            .lcout(),
            .ltout(\c0.n18262_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18262_bdd_4_lut_LC_1_19_4 .C_ON=1'b0;
    defparam \c0.n18262_bdd_4_lut_LC_1_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.n18262_bdd_4_lut_LC_1_19_4 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n18262_bdd_4_lut_LC_1_19_4  (
            .in0(N__32461),
            .in1(N__18015),
            .in2(N__16503),
            .in3(N__16635),
            .lcout(),
            .ltout(\c0.n18265_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i5_LC_1_19_5 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i5_LC_1_19_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i5_LC_1_19_5 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \c0.tx2.r_Tx_Data_i5_LC_1_19_5  (
            .in0(N__16500),
            .in1(N__32462),
            .in2(N__16494),
            .in3(N__32287),
            .lcout(\c0.tx2.r_Tx_Data_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49628),
            .ce(N__24269),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_adj_747_LC_1_20_0 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_adj_747_LC_1_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_adj_747_LC_1_20_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_adj_747_LC_1_20_0  (
            .in0(N__37582),
            .in1(N__37637),
            .in2(N__18426),
            .in3(N__17274),
            .lcout(\c0.n14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_477_LC_1_20_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_477_LC_1_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_477_LC_1_20_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_477_LC_1_20_1  (
            .in0(_gnd_net_),
            .in1(N__17670),
            .in2(_gnd_net_),
            .in3(N__18626),
            .lcout(),
            .ltout(\c0.n10468_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_430_LC_1_20_2 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_430_LC_1_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_430_LC_1_20_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_430_LC_1_20_2  (
            .in0(N__24396),
            .in1(N__18140),
            .in2(N__16491),
            .in3(N__16845),
            .lcout(),
            .ltout(\c0.n15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i166_LC_1_20_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i166_LC_1_20_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i166_LC_1_20_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_frame2_0___i166_LC_1_20_3  (
            .in0(N__16530),
            .in1(N__24705),
            .in2(N__16521),
            .in3(N__20145),
            .lcout(\c0.data_out_frame2_20_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49631),
            .ce(N__26610),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_431_LC_1_20_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_431_LC_1_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_431_LC_1_20_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_431_LC_1_20_5  (
            .in0(N__17273),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37581),
            .lcout(),
            .ltout(\c0.n17306_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i165_LC_1_20_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i165_LC_1_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i165_LC_1_20_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_frame2_0___i165_LC_1_20_6  (
            .in0(N__24942),
            .in1(N__16746),
            .in2(N__16512),
            .in3(N__21870),
            .lcout(\c0.data_out_frame2_20_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49631),
            .ce(N__26610),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_599_LC_1_20_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_599_LC_1_20_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_599_LC_1_20_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_599_LC_1_20_7  (
            .in0(N__21869),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23150),
            .lcout(\c0.n10437 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15288_LC_1_21_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15288_LC_1_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15288_LC_1_21_0 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15288_LC_1_21_0  (
            .in0(N__28684),
            .in1(N__29006),
            .in2(N__20396),
            .in3(N__24032),
            .lcout(\c0.n18064 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_721_LC_1_21_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_721_LC_1_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_721_LC_1_21_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_721_LC_1_21_1  (
            .in0(N__26054),
            .in1(N__24528),
            .in2(N__20439),
            .in3(N__20562),
            .lcout(\c0.n17225 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_3_i5_3_lut_LC_1_21_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_3_i5_3_lut_LC_1_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_3_i5_3_lut_LC_1_21_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_3_i5_3_lut_LC_1_21_2  (
            .in0(N__18425),
            .in1(N__29007),
            .in2(_gnd_net_),
            .in3(N__17529),
            .lcout(\c0.n5_adj_2337 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i105_LC_1_21_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i105_LC_1_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i105_LC_1_21_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_out_frame2_0___i105_LC_1_21_3  (
            .in0(N__17940),
            .in1(N__30921),
            .in2(_gnd_net_),
            .in3(N__26589),
            .lcout(data_out_frame2_13_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49635),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i74_LC_1_21_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i74_LC_1_21_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i74_LC_1_21_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i74_LC_1_21_4  (
            .in0(N__26588),
            .in1(N__30843),
            .in2(_gnd_net_),
            .in3(N__17663),
            .lcout(data_out_frame2_9_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49635),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_586_LC_1_21_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_586_LC_1_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_586_LC_1_21_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_586_LC_1_21_5  (
            .in0(N__17589),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23303),
            .lcout(\c0.n17187 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i150_LC_1_21_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i150_LC_1_21_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i150_LC_1_21_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i150_LC_1_21_6  (
            .in0(N__26587),
            .in1(N__30054),
            .in2(_gnd_net_),
            .in3(N__16577),
            .lcout(data_out_frame2_18_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49635),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_6_i6_4_lut_LC_1_21_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_6_i6_4_lut_LC_1_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_6_i6_4_lut_LC_1_21_7 .LUT_INIT=16'b1111000010001000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_6_i6_4_lut_LC_1_21_7  (
            .in0(N__29008),
            .in1(N__19819),
            .in2(N__16914),
            .in3(N__28685),
            .lcout(\c0.n6_adj_2161 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_422_LC_1_22_0 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_422_LC_1_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_422_LC_1_22_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_adj_422_LC_1_22_0  (
            .in0(N__24653),
            .in1(N__37203),
            .in2(N__16899),
            .in3(N__16560),
            .lcout(),
            .ltout(\c0.n24_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i168_LC_1_22_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i168_LC_1_22_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i168_LC_1_22_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_frame2_0___i168_LC_1_22_1  (
            .in0(N__18030),
            .in1(N__19638),
            .in2(N__16563),
            .in3(N__16811),
            .lcout(\c0.data_out_frame2_20_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49641),
            .ce(N__26611),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_LC_1_22_2 .C_ON=1'b0;
    defparam \c0.i9_4_lut_LC_1_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_LC_1_22_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_LC_1_22_2  (
            .in0(N__17312),
            .in1(N__16554),
            .in2(N__16682),
            .in3(N__23453),
            .lcout(\c0.n22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_648_LC_1_22_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_648_LC_1_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_648_LC_1_22_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_648_LC_1_22_3  (
            .in0(N__20087),
            .in1(N__18210),
            .in2(_gnd_net_),
            .in3(N__21828),
            .lcout(\c0.n17174 ),
            .ltout(\c0.n17174_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_494_LC_1_22_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_494_LC_1_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_494_LC_1_22_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_494_LC_1_22_4  (
            .in0(N__19763),
            .in1(N__20525),
            .in2(N__16548),
            .in3(N__24327),
            .lcout(\c0.n10356 ),
            .ltout(\c0.n10356_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_496_LC_1_22_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_496_LC_1_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_496_LC_1_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i2_3_lut_adj_496_LC_1_22_5  (
            .in0(_gnd_net_),
            .in1(N__18463),
            .in2(N__16545),
            .in3(N__24652),
            .lcout(\c0.n17184 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18136_bdd_4_lut_LC_1_23_0 .C_ON=1'b0;
    defparam \c0.n18136_bdd_4_lut_LC_1_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.n18136_bdd_4_lut_LC_1_23_0 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \c0.n18136_bdd_4_lut_LC_1_23_0  (
            .in0(N__16592),
            .in1(N__28694),
            .in2(N__20438),
            .in3(N__16791),
            .lcout(\c0.n18139 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i126_LC_1_23_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i126_LC_1_23_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i126_LC_1_23_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i126_LC_1_23_1  (
            .in0(N__30599),
            .in1(N__16890),
            .in2(_gnd_net_),
            .in3(N__26597),
            .lcout(data_out_frame2_15_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49647),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i47_LC_1_23_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i47_LC_1_23_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i47_LC_1_23_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i47_LC_1_23_3  (
            .in0(N__31458),
            .in1(N__19817),
            .in2(_gnd_net_),
            .in3(N__26598),
            .lcout(data_out_frame2_5_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49647),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i5_3_lut_LC_1_23_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i5_3_lut_LC_1_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i5_3_lut_LC_1_23_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_4_i5_3_lut_LC_1_23_4  (
            .in0(N__19762),
            .in1(N__29058),
            .in2(_gnd_net_),
            .in3(N__18792),
            .lcout(),
            .ltout(\c0.n5_adj_2315_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14663_4_lut_LC_1_23_5 .C_ON=1'b0;
    defparam \c0.i14663_4_lut_LC_1_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i14663_4_lut_LC_1_23_5 .LUT_INIT=16'b1110001011000000;
    LogicCell40 \c0.i14663_4_lut_LC_1_23_5  (
            .in0(N__29059),
            .in1(N__28695),
            .in2(N__16596),
            .in3(N__21795),
            .lcout(\c0.n17440 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_564_LC_1_23_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_564_LC_1_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_564_LC_1_23_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_564_LC_1_23_6  (
            .in0(_gnd_net_),
            .in1(N__23820),
            .in2(_gnd_net_),
            .in3(N__18080),
            .lcout(\c0.n17132 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i112_LC_1_23_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i112_LC_1_23_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i112_LC_1_23_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i112_LC_1_23_7  (
            .in0(N__31400),
            .in1(N__16593),
            .in2(_gnd_net_),
            .in3(N__26596),
            .lcout(data_out_frame2_13_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49647),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i64_LC_1_24_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i64_LC_1_24_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i64_LC_1_24_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i64_LC_1_24_0  (
            .in0(N__30466),
            .in1(N__17104),
            .in2(_gnd_net_),
            .in3(N__26600),
            .lcout(data_out_frame2_7_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49653),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_478_LC_1_24_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_478_LC_1_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_478_LC_1_24_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_478_LC_1_24_1  (
            .in0(N__16591),
            .in1(N__17540),
            .in2(_gnd_net_),
            .in3(N__24482),
            .lcout(\c0.n17285 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i78_LC_1_24_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i78_LC_1_24_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i78_LC_1_24_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_out_frame2_0___i78_LC_1_24_4  (
            .in0(N__17577),
            .in1(N__31514),
            .in2(_gnd_net_),
            .in3(N__26601),
            .lcout(data_out_frame2_9_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49653),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_683_LC_1_24_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_683_LC_1_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_683_LC_1_24_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_683_LC_1_24_5  (
            .in0(N__17103),
            .in1(N__23296),
            .in2(N__23449),
            .in3(N__17576),
            .lcout(\c0.n10349 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i128_LC_1_24_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i128_LC_1_24_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i128_LC_1_24_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i128_LC_1_24_6  (
            .in0(N__30465),
            .in1(N__24582),
            .in2(_gnd_net_),
            .in3(N__26599),
            .lcout(data_out_frame2_15_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49653),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i15_LC_1_25_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i15_LC_1_25_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i15_LC_1_25_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i15_LC_1_25_0  (
            .in0(_gnd_net_),
            .in1(N__19275),
            .in2(_gnd_net_),
            .in3(N__33220),
            .lcout(\c0.FRAME_MATCHER_i_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49661),
            .ce(),
            .sr(N__20856));
    defparam \c0.FRAME_MATCHER_i_i20_LC_1_26_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i20_LC_1_26_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i20_LC_1_26_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i20_LC_1_26_0  (
            .in0(_gnd_net_),
            .in1(N__19236),
            .in2(_gnd_net_),
            .in3(N__33247),
            .lcout(\c0.FRAME_MATCHER_i_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49669),
            .ce(),
            .sr(N__20757));
    defparam \c0.FRAME_MATCHER_i_i8_LC_1_27_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i8_LC_1_27_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i8_LC_1_27_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i8_LC_1_27_0  (
            .in0(N__19188),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33148),
            .lcout(\c0.FRAME_MATCHER_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49681),
            .ce(),
            .sr(N__20907));
    defparam \c0.FRAME_MATCHER_i_i14_LC_1_28_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i14_LC_1_28_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i14_LC_1_28_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i14_LC_1_28_0  (
            .in0(_gnd_net_),
            .in1(N__19287),
            .in2(_gnd_net_),
            .in3(N__33149),
            .lcout(\c0.FRAME_MATCHER_i_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49692),
            .ce(),
            .sr(N__27957));
    defparam \c0.FRAME_MATCHER_i_i4_LC_1_29_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i4_LC_1_29_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i4_LC_1_29_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i4_LC_1_29_0  (
            .in0(_gnd_net_),
            .in1(N__19008),
            .in2(_gnd_net_),
            .in3(N__33150),
            .lcout(\c0.FRAME_MATCHER_i_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49703),
            .ce(),
            .sr(N__19131));
    defparam \c0.FRAME_MATCHER_i_i11_LC_1_30_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i11_LC_1_30_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i11_LC_1_30_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i11_LC_1_30_0  (
            .in0(_gnd_net_),
            .in1(N__19167),
            .in2(_gnd_net_),
            .in3(N__33151),
            .lcout(\c0.FRAME_MATCHER_i_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49717),
            .ce(),
            .sr(N__20841));
    defparam \c0.FRAME_MATCHER_i_i23_LC_1_31_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i23_LC_1_31_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i23_LC_1_31_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i23_LC_1_31_0  (
            .in0(_gnd_net_),
            .in1(N__19386),
            .in2(_gnd_net_),
            .in3(N__33152),
            .lcout(\c0.FRAME_MATCHER_i_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49728),
            .ce(),
            .sr(N__20967));
    defparam \c0.data_out_5__0__2216_LC_1_32_5 .C_ON=1'b0;
    defparam \c0.data_out_5__0__2216_LC_1_32_5 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_5__0__2216_LC_1_32_5 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \c0.data_out_5__0__2216_LC_1_32_5  (
            .in0(N__48166),
            .in1(N__30873),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.data_out_6__1__N_537 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49738),
            .ce(N__50589),
            .sr(N__42807));
    defparam \c0.data_out_5__7__2209_LC_1_32_6 .C_ON=1'b0;
    defparam \c0.data_out_5__7__2209_LC_1_32_6 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_5__7__2209_LC_1_32_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.data_out_5__7__2209_LC_1_32_6  (
            .in0(_gnd_net_),
            .in1(N__48165),
            .in2(_gnd_net_),
            .in3(N__31344),
            .lcout(\c0.data_out_7__3__N_441 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49738),
            .ce(N__50589),
            .sr(N__42807));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15356_LC_2_17_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15356_LC_2_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15356_LC_2_17_0 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15356_LC_2_17_0  (
            .in0(N__28961),
            .in1(N__18726),
            .in2(N__28675),
            .in3(N__16740),
            .lcout(\c0.n18154 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15250_LC_2_17_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15250_LC_2_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15250_LC_2_17_1 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15250_LC_2_17_1  (
            .in0(N__21572),
            .in1(N__28631),
            .in2(N__20088),
            .in3(N__28962),
            .lcout(\c0.n18022 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_5_i5_3_lut_LC_2_17_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_5_i5_3_lut_LC_2_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_5_i5_3_lut_LC_2_17_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_5_i5_3_lut_LC_2_17_3  (
            .in0(N__28967),
            .in1(N__18303),
            .in2(_gnd_net_),
            .in3(N__21958),
            .lcout(),
            .ltout(\c0.n5_adj_2353_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_5_i6_4_lut_LC_2_17_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_5_i6_4_lut_LC_2_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_5_i6_4_lut_LC_2_17_4 .LUT_INIT=16'b1110001011000000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_5_i6_4_lut_LC_2_17_4  (
            .in0(N__18468),
            .in1(N__28638),
            .in2(N__16638),
            .in3(N__28968),
            .lcout(\c0.n6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_7_i6_4_lut_LC_2_17_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_7_i6_4_lut_LC_2_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_7_i6_4_lut_LC_2_17_6 .LUT_INIT=16'b1011100010001000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_7_i6_4_lut_LC_2_17_6  (
            .in0(N__17085),
            .in1(N__28637),
            .in2(N__18564),
            .in3(N__28966),
            .lcout(\c0.n6_adj_2138 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18034_bdd_4_lut_LC_2_18_0 .C_ON=1'b0;
    defparam \c0.n18034_bdd_4_lut_LC_2_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.n18034_bdd_4_lut_LC_2_18_0 .LUT_INIT=16'b1110111001010000;
    LogicCell40 \c0.n18034_bdd_4_lut_LC_2_18_0  (
            .in0(N__32442),
            .in1(N__16617),
            .in2(N__19701),
            .in3(N__16692),
            .lcout(),
            .ltout(\c0.n18037_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i4_LC_2_18_1 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i4_LC_2_18_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i4_LC_2_18_1 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \c0.tx2.r_Tx_Data_i4_LC_2_18_1  (
            .in0(N__16698),
            .in1(N__32443),
            .in2(N__16602),
            .in3(N__32288),
            .lcout(\c0.tx2.r_Tx_Data_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49629),
            .ce(N__24270),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_LC_2_18_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_LC_2_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_LC_2_18_2 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_LC_2_18_2  (
            .in0(N__18486),
            .in1(N__28639),
            .in2(N__16758),
            .in3(N__29047),
            .lcout(),
            .ltout(\c0.n18274_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18274_bdd_4_lut_LC_2_18_3 .C_ON=1'b0;
    defparam \c0.n18274_bdd_4_lut_LC_2_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.n18274_bdd_4_lut_LC_2_18_3 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n18274_bdd_4_lut_LC_2_18_3  (
            .in0(N__28640),
            .in1(N__18384),
            .in2(N__16599),
            .in3(N__20123),
            .lcout(),
            .ltout(\c0.n18277_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i22_4_lut_LC_2_18_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i22_4_lut_LC_2_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_4_i22_4_lut_LC_2_18_4 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_4_i22_4_lut_LC_2_18_4  (
            .in0(N__32175),
            .in1(N__16713),
            .in2(N__16701),
            .in3(N__21212),
            .lcout(\c0.n22_adj_2367 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15371_LC_2_18_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15371_LC_2_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15371_LC_2_18_5 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_15371_LC_2_18_5  (
            .in0(N__19848),
            .in1(N__32441),
            .in2(N__17346),
            .in3(N__32174),
            .lcout(\c0.n18034 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_667_LC_2_19_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_667_LC_2_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_667_LC_2_19_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_667_LC_2_19_0  (
            .in0(N__23389),
            .in1(N__23190),
            .in2(N__20187),
            .in3(N__20030),
            .lcout(\c0.n17135 ),
            .ltout(\c0.n17135_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_521_LC_2_19_1 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_521_LC_2_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_521_LC_2_19_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_521_LC_2_19_1  (
            .in0(N__18000),
            .in1(N__16686),
            .in2(N__16665),
            .in3(N__17421),
            .lcout(),
            .ltout(\c0.n21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i159_LC_2_19_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i159_LC_2_19_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i159_LC_2_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_out_frame2_0___i159_LC_2_19_2  (
            .in0(_gnd_net_),
            .in1(N__16659),
            .in2(N__16662),
            .in3(N__16653),
            .lcout(\c0.data_out_frame2_19_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49632),
            .ce(N__26564),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_518_LC_2_19_3 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_518_LC_2_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_518_LC_2_19_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i8_4_lut_adj_518_LC_2_19_3  (
            .in0(N__24105),
            .in1(N__24381),
            .in2(N__19941),
            .in3(N__20208),
            .lcout(\c0.n20_adj_2223 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_520_LC_2_19_5 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_520_LC_2_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_520_LC_2_19_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_520_LC_2_19_5  (
            .in0(N__17671),
            .in1(N__16992),
            .in2(N__17739),
            .in3(N__23859),
            .lcout(\c0.n19_adj_2224 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_571_LC_2_20_2 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_571_LC_2_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_571_LC_2_20_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i5_3_lut_adj_571_LC_2_20_2  (
            .in0(N__23207),
            .in1(N__21665),
            .in2(_gnd_net_),
            .in3(N__16980),
            .lcout(),
            .ltout(\c0.n14_adj_2308_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i155_LC_2_20_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i155_LC_2_20_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i155_LC_2_20_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_frame2_0___i155_LC_2_20_3  (
            .in0(N__17481),
            .in1(N__21537),
            .in2(N__16647),
            .in3(N__16821),
            .lcout(\c0.data_out_frame2_19_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49636),
            .ce(N__26608),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_538_LC_2_20_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_538_LC_2_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_538_LC_2_20_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_538_LC_2_20_4  (
            .in0(_gnd_net_),
            .in1(N__21525),
            .in2(_gnd_net_),
            .in3(N__23917),
            .lcout(),
            .ltout(\c0.n17092_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_535_LC_2_20_5 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_535_LC_2_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_535_LC_2_20_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_535_LC_2_20_5  (
            .in0(N__17156),
            .in1(N__16770),
            .in2(N__16764),
            .in3(N__41156),
            .lcout(),
            .ltout(\c0.n17_adj_2294_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i157_LC_2_20_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i157_LC_2_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i157_LC_2_20_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_frame2_0___i157_LC_2_20_6  (
            .in0(N__23208),
            .in1(N__17292),
            .in2(N__16761),
            .in3(N__16719),
            .lcout(\c0.data_out_frame2_19_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49636),
            .ce(N__26608),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_LC_2_21_0 .C_ON=1'b0;
    defparam \c0.i5_4_lut_LC_2_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_LC_2_21_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_LC_2_21_0  (
            .in0(N__23694),
            .in1(N__17402),
            .in2(N__20026),
            .in3(N__18231),
            .lcout(\c0.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i113_LC_2_21_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i113_LC_2_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i113_LC_2_21_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i113_LC_2_21_1  (
            .in0(N__30413),
            .in1(N__16739),
            .in2(_gnd_net_),
            .in3(N__26555),
            .lcout(data_out_frame2_14_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49642),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i52_LC_2_21_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i52_LC_2_21_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i52_LC_2_21_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i52_LC_2_21_2  (
            .in0(N__26554),
            .in1(N__31209),
            .in2(_gnd_net_),
            .in3(N__17533),
            .lcout(data_out_frame2_6_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49642),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_608_LC_2_21_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_608_LC_2_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_608_LC_2_21_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_608_LC_2_21_3  (
            .in0(N__17817),
            .in1(N__23024),
            .in2(_gnd_net_),
            .in3(N__16738),
            .lcout(\c0.n17237 ),
            .ltout(\c0.n17237_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_456_LC_2_21_4 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_456_LC_2_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_456_LC_2_21_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_456_LC_2_21_4  (
            .in0(N__24098),
            .in1(N__16959),
            .in2(N__16722),
            .in3(N__18957),
            .lcout(\c0.n17165 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i135_LC_2_21_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i135_LC_2_21_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i135_LC_2_21_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_out_frame2_0___i135_LC_2_21_5  (
            .in0(N__17818),
            .in1(N__29993),
            .in2(_gnd_net_),
            .in3(N__26556),
            .lcout(data_out_frame2_16_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49642),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_534_LC_2_21_6 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_534_LC_2_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_534_LC_2_21_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_534_LC_2_21_6  (
            .in0(N__18753),
            .in1(N__24782),
            .in2(N__23151),
            .in3(N__16960),
            .lcout(\c0.n16_adj_2293 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i66_LC_2_21_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i66_LC_2_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i66_LC_2_21_7 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \c0.data_out_frame2_0___i66_LC_2_21_7  (
            .in0(N__30278),
            .in1(_gnd_net_),
            .in2(N__18085),
            .in3(N__26557),
            .lcout(data_out_frame2_8_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49642),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15341_LC_2_22_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15341_LC_2_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15341_LC_2_22_0 .LUT_INIT=16'b1010111111000000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15341_LC_2_22_0  (
            .in0(N__24583),
            .in1(N__22095),
            .in2(N__28683),
            .in3(N__29024),
            .lcout(\c0.n18136 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_650_LC_2_22_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_650_LC_2_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_650_LC_2_22_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_650_LC_2_22_1  (
            .in0(N__18791),
            .in1(N__24852),
            .in2(N__21369),
            .in3(N__20241),
            .lcout(\c0.n17228 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15259_LC_2_22_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15259_LC_2_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15259_LC_2_22_2 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15259_LC_2_22_2  (
            .in0(N__28655),
            .in1(N__20580),
            .in2(N__16785),
            .in3(N__29023),
            .lcout(\c0.n18028 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_685_LC_2_22_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_685_LC_2_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_685_LC_2_22_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_685_LC_2_22_4  (
            .in0(N__23815),
            .in1(N__18061),
            .in2(_gnd_net_),
            .in3(N__21467),
            .lcout(\c0.n10371 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_553_LC_2_22_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_553_LC_2_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_553_LC_2_22_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_553_LC_2_22_5  (
            .in0(N__21364),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20240),
            .lcout(\c0.n10462 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i57_LC_2_22_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i57_LC_2_22_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i57_LC_2_22_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i57_LC_2_22_6  (
            .in0(N__29874),
            .in1(N__16961),
            .in2(_gnd_net_),
            .in3(N__26538),
            .lcout(data_out_frame2_7_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49648),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_LC_2_22_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_LC_2_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_LC_2_22_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_LC_2_22_7  (
            .in0(N__18556),
            .in1(N__18835),
            .in2(_gnd_net_),
            .in3(N__17588),
            .lcout(\c0.n17138 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i116_LC_2_23_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i116_LC_2_23_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i116_LC_2_23_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i116_LC_2_23_0  (
            .in0(N__31208),
            .in1(N__17271),
            .in2(_gnd_net_),
            .in3(N__26561),
            .lcout(data_out_frame2_14_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49654),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_614_LC_2_23_1 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_614_LC_2_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_614_LC_2_23_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_614_LC_2_23_1  (
            .in0(N__19880),
            .in1(N__21457),
            .in2(N__16938),
            .in3(N__17105),
            .lcout(\c0.n10424 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_530_LC_2_23_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_530_LC_2_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_530_LC_2_23_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_530_LC_2_23_3  (
            .in0(_gnd_net_),
            .in1(N__23725),
            .in2(_gnd_net_),
            .in3(N__21753),
            .lcout(),
            .ltout(\c0.n10520_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_484_LC_2_23_4 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_484_LC_2_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_484_LC_2_23_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i9_4_lut_adj_484_LC_2_23_4  (
            .in0(N__18664),
            .in1(N__23396),
            .in2(N__16848),
            .in3(N__16937),
            .lcout(\c0.n25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_592_LC_2_23_5 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_592_LC_2_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_592_LC_2_23_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_592_LC_2_23_5  (
            .in0(N__17352),
            .in1(N__16841),
            .in2(N__20397),
            .in3(N__21824),
            .lcout(\c0.n17216 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_524_LC_2_23_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_524_LC_2_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_524_LC_2_23_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_524_LC_2_23_6  (
            .in0(N__22972),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20124),
            .lcout(\c0.n10572 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_578_LC_2_23_7 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_578_LC_2_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_578_LC_2_23_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_578_LC_2_23_7  (
            .in0(N__17502),
            .in1(N__24879),
            .in2(N__40842),
            .in3(N__16830),
            .lcout(\c0.n15_adj_2312 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_483_LC_2_24_0 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_483_LC_2_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_483_LC_2_24_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_adj_483_LC_2_24_0  (
            .in0(N__27595),
            .in1(N__17609),
            .in2(N__16812),
            .in3(N__18260),
            .lcout(\c0.n27_adj_2204 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_492_LC_2_24_1 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_492_LC_2_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_492_LC_2_24_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_492_LC_2_24_1  (
            .in0(N__17909),
            .in1(N__18421),
            .in2(N__18952),
            .in3(N__18837),
            .lcout(\c0.n10_adj_2207 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i80_LC_2_24_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i80_LC_2_24_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i80_LC_2_24_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i80_LC_2_24_3  (
            .in0(N__31392),
            .in1(N__23448),
            .in2(_gnd_net_),
            .in3(N__26562),
            .lcout(data_out_frame2_9_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49662),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_476_LC_2_24_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_476_LC_2_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_476_LC_2_24_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_476_LC_2_24_5  (
            .in0(_gnd_net_),
            .in1(N__23960),
            .in2(_gnd_net_),
            .in3(N__21956),
            .lcout(\c0.n10346 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_516_LC_2_24_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_516_LC_2_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_516_LC_2_24_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_516_LC_2_24_6  (
            .in0(_gnd_net_),
            .in1(N__16891),
            .in2(_gnd_net_),
            .in3(N__22921),
            .lcout(\c0.n10530 ),
            .ltout(\c0.n10530_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_692_LC_2_24_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_692_LC_2_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_692_LC_2_24_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_692_LC_2_24_7  (
            .in0(N__19818),
            .in1(N__19905),
            .in2(N__16983),
            .in3(N__16979),
            .lcout(\c0.n17303 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_0_i5_3_lut_LC_2_25_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_0_i5_3_lut_LC_2_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_0_i5_3_lut_LC_2_25_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_0_i5_3_lut_LC_2_25_1  (
            .in0(N__16962),
            .in1(N__16932),
            .in2(_gnd_net_),
            .in3(N__29050),
            .lcout(\c0.n5_adj_2217 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i49_LC_2_25_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i49_LC_2_25_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i49_LC_2_25_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_out_frame2_0___i49_LC_2_25_2  (
            .in0(N__16933),
            .in1(N__30405),
            .in2(_gnd_net_),
            .in3(N__26563),
            .lcout(data_out_frame2_6_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49670),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_6_i5_3_lut_LC_2_25_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_6_i5_3_lut_LC_2_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_6_i5_3_lut_LC_2_25_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_6_i5_3_lut_LC_2_25_4  (
            .in0(N__29049),
            .in1(N__40892),
            .in2(_gnd_net_),
            .in3(N__18836),
            .lcout(\c0.n5_adj_2343 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15311_LC_2_25_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15311_LC_2_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15311_LC_2_25_5 .LUT_INIT=16'b1101101011010000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15311_LC_2_25_5  (
            .in0(N__28659),
            .in1(N__16898),
            .in2(N__29073),
            .in3(N__17869),
            .lcout(),
            .ltout(\c0.n18100_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18100_bdd_4_lut_LC_2_25_6 .C_ON=1'b0;
    defparam \c0.n18100_bdd_4_lut_LC_2_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.n18100_bdd_4_lut_LC_2_25_6 .LUT_INIT=16'b1111000011001010;
    LogicCell40 \c0.n18100_bdd_4_lut_LC_2_25_6  (
            .in0(N__20166),
            .in1(N__23723),
            .in2(N__16866),
            .in3(N__28660),
            .lcout(\c0.n18103 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i28_LC_2_26_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i28_LC_2_26_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i28_LC_2_26_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i28_LC_2_26_0  (
            .in0(_gnd_net_),
            .in1(N__41556),
            .in2(_gnd_net_),
            .in3(N__35200),
            .lcout(\c0.FRAME_MATCHER_state_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49682),
            .ce(),
            .sr(N__33600));
    defparam \c0.FRAME_MATCHER_i_i19_LC_2_27_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i19_LC_2_27_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i19_LC_2_27_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i19_LC_2_27_0  (
            .in0(_gnd_net_),
            .in1(N__19251),
            .in2(_gnd_net_),
            .in3(N__33221),
            .lcout(\c0.FRAME_MATCHER_i_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49693),
            .ce(),
            .sr(N__20826));
    defparam \c0.FRAME_MATCHER_i_i13_LC_2_28_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i13_LC_2_28_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i13_LC_2_28_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i13_LC_2_28_0  (
            .in0(N__33223),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19143),
            .lcout(\c0.FRAME_MATCHER_i_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49704),
            .ce(),
            .sr(N__17718));
    defparam \c0.FRAME_MATCHER_i_i1_LC_2_29_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i1_LC_2_29_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i1_LC_2_29_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i1_LC_2_29_0  (
            .in0(_gnd_net_),
            .in1(N__19107),
            .in2(_gnd_net_),
            .in3(N__33225),
            .lcout(\c0.FRAME_MATCHER_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49718),
            .ce(),
            .sr(N__25392));
    defparam \c0.FRAME_MATCHER_i_i28_LC_2_30_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i28_LC_2_30_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i28_LC_2_30_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i28_LC_2_30_0  (
            .in0(_gnd_net_),
            .in1(N__19359),
            .in2(_gnd_net_),
            .in3(N__33252),
            .lcout(\c0.FRAME_MATCHER_i_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49729),
            .ce(),
            .sr(N__22464));
    defparam \c0.FRAME_MATCHER_state_i16_LC_2_31_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i16_LC_2_31_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i16_LC_2_31_0 .LUT_INIT=16'b1110000011000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i16_LC_2_31_0  (
            .in0(N__45036),
            .in1(N__44817),
            .in2(N__37793),
            .in3(N__44611),
            .lcout(\c0.FRAME_MATCHER_state_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49739),
            .ce(),
            .sr(N__33582));
    defparam \c0.data_out_7__3__2197_LC_2_32_0 .C_ON=1'b0;
    defparam \c0.data_out_7__3__2197_LC_2_32_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__3__2197_LC_2_32_0 .LUT_INIT=16'b1100000011100010;
    LogicCell40 \c0.data_out_7__3__2197_LC_2_32_0  (
            .in0(N__48426),
            .in1(N__50337),
            .in2(N__31995),
            .in3(N__46476),
            .lcout(\c0.data_out_7_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49750),
            .ce(N__46935),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i1_LC_3_16_7 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i1_LC_3_16_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i1_LC_3_16_7 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \c0.tx2.r_Tx_Data_i1_LC_3_16_7  (
            .in0(N__17121),
            .in1(N__32424),
            .in2(N__17010),
            .in3(N__32275),
            .lcout(\c0.tx2.r_Tx_Data_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49633),
            .ce(N__24273),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15240_LC_3_17_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15240_LC_3_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15240_LC_3_17_0 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15240_LC_3_17_0  (
            .in0(N__29057),
            .in1(N__18249),
            .in2(N__28676),
            .in3(N__19587),
            .lcout(),
            .ltout(\c0.n18010_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18010_bdd_4_lut_LC_3_17_1 .C_ON=1'b0;
    defparam \c0.n18010_bdd_4_lut_LC_3_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.n18010_bdd_4_lut_LC_3_17_1 .LUT_INIT=16'b1111000010101100;
    LogicCell40 \c0.n18010_bdd_4_lut_LC_3_17_1  (
            .in0(N__19926),
            .in1(N__18627),
            .in2(N__17016),
            .in3(N__28636),
            .lcout(),
            .ltout(\c0.n18013_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_1_i22_4_lut_LC_3_17_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_1_i22_4_lut_LC_3_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_1_i22_4_lut_LC_3_17_2 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_1_i22_4_lut_LC_3_17_2  (
            .in0(N__21199),
            .in1(N__32153),
            .in2(N__17013),
            .in3(N__17973),
            .lcout(\c0.n22_adj_2375 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15425_LC_3_17_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15425_LC_3_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15425_LC_3_17_3 .LUT_INIT=16'b1111100000111000;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_15425_LC_3_17_3  (
            .in0(N__17001),
            .in1(N__32446),
            .in2(N__32170),
            .in3(N__23577),
            .lcout(),
            .ltout(\c0.n18238_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18238_bdd_4_lut_LC_3_17_4 .C_ON=1'b0;
    defparam \c0.n18238_bdd_4_lut_LC_3_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.n18238_bdd_4_lut_LC_3_17_4 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n18238_bdd_4_lut_LC_3_17_4  (
            .in0(N__32447),
            .in1(N__23061),
            .in2(N__17124),
            .in3(N__23349),
            .lcout(\c0.n18241 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_7_i5_3_lut_LC_3_17_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_7_i5_3_lut_LC_3_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_7_i5_3_lut_LC_3_17_5 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_7_i5_3_lut_LC_3_17_5  (
            .in0(N__18665),
            .in1(_gnd_net_),
            .in2(N__29022),
            .in3(N__17115),
            .lcout(\c0.n5_adj_2137 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18154_bdd_4_lut_LC_3_17_7 .C_ON=1'b0;
    defparam \c0.n18154_bdd_4_lut_LC_3_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.n18154_bdd_4_lut_LC_3_17_7 .LUT_INIT=16'b1010101011100100;
    LogicCell40 \c0.n18154_bdd_4_lut_LC_3_17_7  (
            .in0(N__17076),
            .in1(N__26053),
            .in2(N__17959),
            .in3(N__28632),
            .lcout(\c0.n18157 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15336_LC_3_18_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15336_LC_3_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15336_LC_3_18_0 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15336_LC_3_18_0  (
            .in0(N__28549),
            .in1(N__22005),
            .in2(N__17238),
            .in3(N__29056),
            .lcout(),
            .ltout(\c0.n18130_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18130_bdd_4_lut_LC_3_18_1 .C_ON=1'b0;
    defparam \c0.n18130_bdd_4_lut_LC_3_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.n18130_bdd_4_lut_LC_3_18_1 .LUT_INIT=16'b1111000010101100;
    LogicCell40 \c0.n18130_bdd_4_lut_LC_3_18_1  (
            .in0(N__18363),
            .in1(N__27655),
            .in2(N__17070),
            .in3(N__28550),
            .lcout(),
            .ltout(\c0.n18133_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_7_i22_4_lut_LC_3_18_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_7_i22_4_lut_LC_3_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_7_i22_4_lut_LC_3_18_2 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_7_i22_4_lut_LC_3_18_2  (
            .in0(N__17067),
            .in1(N__21203),
            .in2(N__17052),
            .in3(N__32169),
            .lcout(\c0.n22_adj_2363 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18028_bdd_4_lut_LC_3_18_4 .C_ON=1'b0;
    defparam \c0.n18028_bdd_4_lut_LC_3_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.n18028_bdd_4_lut_LC_3_18_4 .LUT_INIT=16'b1101100111001000;
    LogicCell40 \c0.n18028_bdd_4_lut_LC_3_18_4  (
            .in0(N__28548),
            .in1(N__17037),
            .in2(N__21984),
            .in3(N__20339),
            .lcout(\c0.n18031 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15264_LC_3_18_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15264_LC_3_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15264_LC_3_18_6 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15264_LC_3_18_6  (
            .in0(N__28546),
            .in1(N__21666),
            .in2(N__20625),
            .in3(N__29055),
            .lcout(),
            .ltout(\c0.n18040_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18040_bdd_4_lut_LC_3_18_7 .C_ON=1'b0;
    defparam \c0.n18040_bdd_4_lut_LC_3_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.n18040_bdd_4_lut_LC_3_18_7 .LUT_INIT=16'b1111000010101100;
    LogicCell40 \c0.n18040_bdd_4_lut_LC_3_18_7  (
            .in0(N__17456),
            .in1(N__23916),
            .in2(N__17019),
            .in3(N__28547),
            .lcout(\c0.n18043 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_502_LC_3_19_0 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_502_LC_3_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_502_LC_3_19_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_502_LC_3_19_0  (
            .in0(N__17184),
            .in1(N__40273),
            .in2(N__23046),
            .in3(N__17178),
            .lcout(\c0.n10263 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_500_LC_3_19_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_500_LC_3_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_500_LC_3_19_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_500_LC_3_19_1  (
            .in0(_gnd_net_),
            .in1(N__37587),
            .in2(_gnd_net_),
            .in3(N__40103),
            .lcout(\c0.n6_adj_2215 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_525_LC_3_19_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_525_LC_3_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_525_LC_3_19_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_525_LC_3_19_2  (
            .in0(_gnd_net_),
            .in1(N__17882),
            .in2(_gnd_net_),
            .in3(N__23259),
            .lcout(\c0.n17141 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_499_LC_3_19_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_499_LC_3_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_499_LC_3_19_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_499_LC_3_19_4  (
            .in0(N__37638),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34326),
            .lcout(\c0.n17219 ),
            .ltout(\c0.n17219_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_LC_3_19_5 .C_ON=1'b0;
    defparam \c0.i7_4_lut_LC_3_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_LC_3_19_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_LC_3_19_5  (
            .in0(N__18956),
            .in1(N__17172),
            .in2(N__17163),
            .in3(N__20340),
            .lcout(),
            .ltout(\c0.n17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i167_LC_3_19_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i167_LC_3_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i167_LC_3_19_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_frame2_0___i167_LC_3_19_6  (
            .in0(N__18312),
            .in1(N__24698),
            .in2(N__17160),
            .in3(N__17388),
            .lcout(\c0.data_out_frame2_20_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49637),
            .ce(N__26609),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_505_LC_3_20_0 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_505_LC_3_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_505_LC_3_20_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i11_4_lut_adj_505_LC_3_20_0  (
            .in0(N__18560),
            .in1(N__23654),
            .in2(N__40680),
            .in3(N__22937),
            .lcout(\c0.n30_adj_2218 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_503_LC_3_20_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_503_LC_3_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_503_LC_3_20_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_503_LC_3_20_1  (
            .in0(_gnd_net_),
            .in1(N__20284),
            .in2(_gnd_net_),
            .in3(N__17958),
            .lcout(),
            .ltout(\c0.n17246_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_adj_508_LC_3_20_2 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_508_LC_3_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_508_LC_3_20_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i14_4_lut_adj_508_LC_3_20_2  (
            .in0(N__17157),
            .in1(N__17477),
            .in2(N__17139),
            .in3(N__17136),
            .lcout(),
            .ltout(\c0.n33_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i160_LC_3_20_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i160_LC_3_20_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i160_LC_3_20_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_frame2_0___i160_LC_3_20_3  (
            .in0(N__17217),
            .in1(N__23676),
            .in2(N__17241),
            .in3(N__18123),
            .lcout(\c0.data_out_frame2_19_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49643),
            .ce(N__26607),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_504_LC_3_20_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_504_LC_3_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_504_LC_3_20_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_504_LC_3_20_4  (
            .in0(_gnd_net_),
            .in1(N__23019),
            .in2(_gnd_net_),
            .in3(N__21957),
            .lcout(),
            .ltout(\c0.n17300_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_adj_507_LC_3_20_5 .C_ON=1'b0;
    defparam \c0.i15_4_lut_adj_507_LC_3_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_adj_507_LC_3_20_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i15_4_lut_adj_507_LC_3_20_5  (
            .in0(N__17226),
            .in1(N__19829),
            .in2(N__17220),
            .in3(N__23186),
            .lcout(\c0.n34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_664_LC_3_21_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_664_LC_3_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_664_LC_3_21_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_664_LC_3_21_0  (
            .in0(N__20332),
            .in1(N__24426),
            .in2(_gnd_net_),
            .in3(N__20619),
            .lcout(\c0.n17291 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15269_LC_3_21_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15269_LC_3_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15269_LC_3_21_1 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15269_LC_3_21_1  (
            .in0(N__29004),
            .in1(N__20230),
            .in2(N__28654),
            .in3(N__18201),
            .lcout(\c0.n18046 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_LC_3_21_2 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_LC_3_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_LC_3_21_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_LC_3_21_2  (
            .in0(N__18202),
            .in1(N__24498),
            .in2(N__17211),
            .in3(N__21820),
            .lcout(\c0.n14_adj_2346 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15279_LC_3_21_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15279_LC_3_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15279_LC_3_21_3 .LUT_INIT=16'b1110010010101010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15279_LC_3_21_3  (
            .in0(N__29005),
            .in1(N__17272),
            .in2(N__24433),
            .in3(N__28596),
            .lcout(\c0.n18058 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_450_LC_3_21_4 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_450_LC_3_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_450_LC_3_21_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_450_LC_3_21_4  (
            .in0(N__18893),
            .in1(N__20460),
            .in2(N__17199),
            .in3(N__17628),
            .lcout(\c0.n15_adj_2185 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i101_LC_3_21_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i101_LC_3_21_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i101_LC_3_21_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i101_LC_3_21_5  (
            .in0(N__30110),
            .in1(N__20012),
            .in2(_gnd_net_),
            .in3(N__26459),
            .lcout(data_out_frame2_12_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49649),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18076_bdd_4_lut_LC_3_21_6 .C_ON=1'b0;
    defparam \c0.n18076_bdd_4_lut_LC_3_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.n18076_bdd_4_lut_LC_3_21_6 .LUT_INIT=16'b1111110000100010;
    LogicCell40 \c0.n18076_bdd_4_lut_LC_3_21_6  (
            .in0(N__20011),
            .in1(N__28589),
            .in2(N__41157),
            .in3(N__17598),
            .lcout(\c0.n17569 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i142_LC_3_21_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i142_LC_3_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i142_LC_3_21_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i142_LC_3_21_7  (
            .in0(N__30598),
            .in1(N__17327),
            .in2(_gnd_net_),
            .in3(N__26460),
            .lcout(data_out_frame2_17_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49649),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_438_LC_3_22_0 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_438_LC_3_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_438_LC_3_22_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_438_LC_3_22_0  (
            .in0(N__18230),
            .in1(N__24551),
            .in2(N__17313),
            .in3(N__17613),
            .lcout(\c0.n12_adj_2178 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_706_LC_3_22_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_706_LC_3_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_706_LC_3_22_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_706_LC_3_22_1  (
            .in0(N__23484),
            .in1(N__24483),
            .in2(_gnd_net_),
            .in3(N__24434),
            .lcout(\c0.n17312 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_527_LC_3_22_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_527_LC_3_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_527_LC_3_22_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_527_LC_3_22_3  (
            .in0(_gnd_net_),
            .in1(N__24367),
            .in2(_gnd_net_),
            .in3(N__18299),
            .lcout(),
            .ltout(\c0.n6_adj_2228_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_528_LC_3_22_4 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_528_LC_3_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_528_LC_3_22_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_528_LC_3_22_4  (
            .in0(N__24176),
            .in1(N__18323),
            .in2(N__17295),
            .in3(N__17285),
            .lcout(\c0.n17116 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_513_LC_3_22_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_513_LC_3_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_513_LC_3_22_5 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \c0.i1_2_lut_adj_513_LC_3_22_5  (
            .in0(N__24748),
            .in1(N__22973),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.n17279 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_722_LC_3_22_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_722_LC_3_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_722_LC_3_22_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_722_LC_3_22_6  (
            .in0(N__40863),
            .in1(N__21300),
            .in2(N__40934),
            .in3(N__20517),
            .lcout(\c0.n17309 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_545_LC_3_22_7 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_545_LC_3_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_545_LC_3_22_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_545_LC_3_22_7  (
            .in0(N__18177),
            .in1(N__17265),
            .in2(N__18084),
            .in3(N__40929),
            .lcout(\c0.n12_adj_2298 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_682_LC_3_23_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_682_LC_3_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_682_LC_3_23_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_682_LC_3_23_0  (
            .in0(N__26052),
            .in1(N__23239),
            .in2(_gnd_net_),
            .in3(N__21573),
            .lcout(\c0.n17194 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_684_LC_3_23_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_684_LC_3_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_684_LC_3_23_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_684_LC_3_23_1  (
            .in0(N__17442),
            .in1(N__24905),
            .in2(N__18730),
            .in3(N__17828),
            .lcout(\c0.n17267 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_549_LC_3_23_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_549_LC_3_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_549_LC_3_23_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_549_LC_3_23_2  (
            .in0(N__24904),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17441),
            .lcout(\c0.n17168 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i107_LC_3_23_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i107_LC_3_23_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i107_LC_3_23_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_out_frame2_0___i107_LC_3_23_3  (
            .in0(N__17443),
            .in1(N__31675),
            .in2(_gnd_net_),
            .in3(N__26583),
            .lcout(data_out_frame2_13_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49663),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_481_LC_3_23_4 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_481_LC_3_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_481_LC_3_23_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_4_lut_adj_481_LC_3_23_4  (
            .in0(N__17414),
            .in1(N__17403),
            .in2(N__41055),
            .in3(N__17381),
            .lcout(),
            .ltout(\c0.n28_adj_2200_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_LC_3_23_5 .C_ON=1'b0;
    defparam \c0.i15_4_lut_LC_3_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_LC_3_23_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i15_4_lut_LC_3_23_5  (
            .in0(N__17370),
            .in1(N__18570),
            .in2(N__17364),
            .in3(N__17361),
            .lcout(\c0.n10223 ),
            .ltout(\c0.n10223_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_adj_729_LC_3_23_6 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_adj_729_LC_3_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_adj_729_LC_3_23_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_adj_729_LC_3_23_6  (
            .in0(N__18722),
            .in1(N__18464),
            .in2(N__17355),
            .in3(N__23666),
            .lcout(\c0.n14_adj_2206 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_591_LC_3_23_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_591_LC_3_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_591_LC_3_23_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_591_LC_3_23_7  (
            .in0(_gnd_net_),
            .in1(N__18288),
            .in2(_gnd_net_),
            .in3(N__20557),
            .lcout(\c0.n6_adj_2318 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i75_LC_3_24_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i75_LC_3_24_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i75_LC_3_24_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i75_LC_3_24_0  (
            .in0(N__26580),
            .in1(N__31676),
            .in2(_gnd_net_),
            .in3(N__18950),
            .lcout(data_out_frame2_9_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49671),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i111_LC_3_24_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i111_LC_3_24_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i111_LC_3_24_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i111_LC_3_24_1  (
            .in0(N__31453),
            .in1(N__22927),
            .in2(_gnd_net_),
            .in3(N__26581),
            .lcout(data_out_frame2_13_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49671),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_556_LC_3_24_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_556_LC_3_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_556_LC_3_24_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_556_LC_3_24_2  (
            .in0(_gnd_net_),
            .in1(N__18619),
            .in2(_gnd_net_),
            .in3(N__23958),
            .lcout(\c0.n10533 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_734_LC_3_24_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_734_LC_3_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_734_LC_3_24_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_734_LC_3_24_3  (
            .in0(N__18618),
            .in1(N__17672),
            .in2(N__18517),
            .in3(N__17624),
            .lcout(\c0.n17231 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15301_LC_3_24_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15301_LC_3_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15301_LC_3_24_4 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15301_LC_3_24_4  (
            .in0(N__24783),
            .in1(N__28662),
            .in2(N__20526),
            .in3(N__29054),
            .lcout(\c0.n18076 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18106_bdd_4_lut_LC_3_24_5 .C_ON=1'b0;
    defparam \c0.n18106_bdd_4_lut_LC_3_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.n18106_bdd_4_lut_LC_3_24_5 .LUT_INIT=16'b1101110010011000;
    LogicCell40 \c0.n18106_bdd_4_lut_LC_3_24_5  (
            .in0(N__28663),
            .in1(N__20352),
            .in2(N__40938),
            .in3(N__17587),
            .lcout(\c0.n18109 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_2_lut_3_lut_LC_3_24_6 .C_ON=1'b0;
    defparam \c0.i2_2_lut_3_lut_LC_3_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_2_lut_3_lut_LC_3_24_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_2_lut_3_lut_LC_3_24_6  (
            .in0(N__27648),
            .in1(N__24079),
            .in2(_gnd_net_),
            .in3(N__27596),
            .lcout(\c0.n10_adj_2297 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i118_LC_3_24_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i118_LC_3_24_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i118_LC_3_24_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i118_LC_3_24_7  (
            .in0(N__31089),
            .in1(N__17875),
            .in2(_gnd_net_),
            .in3(N__26582),
            .lcout(data_out_frame2_14_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49671),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_699_LC_3_25_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_699_LC_3_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_699_LC_3_25_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_699_LC_3_25_0  (
            .in0(N__21522),
            .in1(N__23903),
            .in2(_gnd_net_),
            .in3(N__20019),
            .lcout(\c0.n10334 ),
            .ltout(\c0.n10334_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_542_LC_3_25_1 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_542_LC_3_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_542_LC_3_25_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_542_LC_3_25_1  (
            .in0(N__18743),
            .in1(N__17541),
            .in2(N__17505),
            .in3(N__17501),
            .lcout(),
            .ltout(\c0.n14_adj_2296_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_544_LC_3_25_2 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_544_LC_3_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_544_LC_3_25_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_544_LC_3_25_2  (
            .in0(N__18519),
            .in1(N__17490),
            .in2(N__17484),
            .in3(N__23447),
            .lcout(\c0.n17171 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i121_LC_3_25_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i121_LC_3_25_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i121_LC_3_25_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i121_LC_3_25_3  (
            .in0(N__26559),
            .in1(N__29872),
            .in2(_gnd_net_),
            .in3(N__18712),
            .lcout(data_out_frame2_15_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49683),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i102_LC_3_25_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i102_LC_3_25_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i102_LC_3_25_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i102_LC_3_25_4  (
            .in0(N__30049),
            .in1(N__20167),
            .in2(_gnd_net_),
            .in3(N__26560),
            .lcout(data_out_frame2_12_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49683),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i110_LC_3_25_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i110_LC_3_25_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i110_LC_3_25_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i110_LC_3_25_5  (
            .in0(N__26558),
            .in1(N__31506),
            .in2(_gnd_net_),
            .in3(N__23724),
            .lcout(data_out_frame2_13_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49683),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.o_Tx_Serial_I_0_1_lut_LC_3_25_6 .C_ON=1'b0;
    defparam \c0.tx2.o_Tx_Serial_I_0_1_lut_LC_3_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.o_Tx_Serial_I_0_1_lut_LC_3_25_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \c0.tx2.o_Tx_Serial_I_0_1_lut_LC_3_25_6  (
            .in0(N__22121),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(tx2_enable),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i3_LC_3_26_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i3_LC_3_26_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i3_LC_3_26_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i3_LC_3_26_0  (
            .in0(_gnd_net_),
            .in1(N__19056),
            .in2(_gnd_net_),
            .in3(N__33246),
            .lcout(\c0.FRAME_MATCHER_i_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49694),
            .ce(),
            .sr(N__18843));
    defparam \c0.FRAME_MATCHER_i_i7_LC_3_27_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i7_LC_3_27_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i7_LC_3_27_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i7_LC_3_27_0  (
            .in0(_gnd_net_),
            .in1(N__19197),
            .in2(_gnd_net_),
            .in3(N__33219),
            .lcout(\c0.FRAME_MATCHER_i_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49705),
            .ce(),
            .sr(N__17724));
    defparam \c0.i18_4_lut_adj_674_LC_3_28_0 .C_ON=1'b0;
    defparam \c0.i18_4_lut_adj_674_LC_3_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.i18_4_lut_adj_674_LC_3_28_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i18_4_lut_adj_674_LC_3_28_0  (
            .in0(N__27081),
            .in1(N__25867),
            .in2(N__27206),
            .in3(N__19326),
            .lcout(\c0.n43_adj_2380 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i29_LC_3_28_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i29_LC_3_28_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i29_LC_3_28_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i29_LC_3_28_1  (
            .in0(_gnd_net_),
            .in1(N__19311),
            .in2(_gnd_net_),
            .in3(N__33222),
            .lcout(\c0.FRAME_MATCHER_i_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49719),
            .ce(),
            .sr(N__17682));
    defparam \c0.select_219_Select_29_i3_2_lut_3_lut_LC_3_28_2 .C_ON=1'b0;
    defparam \c0.select_219_Select_29_i3_2_lut_3_lut_LC_3_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.select_219_Select_29_i3_2_lut_3_lut_LC_3_28_2 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \c0.select_219_Select_29_i3_2_lut_3_lut_LC_3_28_2  (
            .in0(N__41906),
            .in1(N__27840),
            .in2(_gnd_net_),
            .in3(N__19328),
            .lcout(\c0.n3_adj_2232 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10659_2_lut_LC_3_28_3 .C_ON=1'b0;
    defparam \c0.i10659_2_lut_LC_3_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.i10659_2_lut_LC_3_28_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i10659_2_lut_LC_3_28_3  (
            .in0(N__19327),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41903),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_219_Select_7_i3_2_lut_3_lut_LC_3_28_5 .C_ON=1'b0;
    defparam \c0.select_219_Select_7_i3_2_lut_3_lut_LC_3_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.select_219_Select_7_i3_2_lut_3_lut_LC_3_28_5 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \c0.select_219_Select_7_i3_2_lut_3_lut_LC_3_28_5  (
            .in0(N__27842),
            .in1(N__27082),
            .in2(_gnd_net_),
            .in3(N__41907),
            .lcout(\c0.n3_adj_2278 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_219_Select_13_i3_2_lut_3_lut_LC_3_28_6 .C_ON=1'b0;
    defparam \c0.select_219_Select_13_i3_2_lut_3_lut_LC_3_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.select_219_Select_13_i3_2_lut_3_lut_LC_3_28_6 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \c0.select_219_Select_13_i3_2_lut_3_lut_LC_3_28_6  (
            .in0(N__41905),
            .in1(N__27198),
            .in2(_gnd_net_),
            .in3(N__27841),
            .lcout(\c0.n3_adj_2266 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10676_2_lut_LC_3_28_7 .C_ON=1'b0;
    defparam \c0.i10676_2_lut_LC_3_28_7 .SEQ_MODE=4'b0000;
    defparam \c0.i10676_2_lut_LC_3_28_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i10676_2_lut_LC_3_28_7  (
            .in0(N__25868),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41904),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i22_LC_3_29_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i22_LC_3_29_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i22_LC_3_29_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i22_LC_3_29_0  (
            .in0(_gnd_net_),
            .in1(N__19209),
            .in2(_gnd_net_),
            .in3(N__33224),
            .lcout(\c0.FRAME_MATCHER_i_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49730),
            .ce(),
            .sr(N__25362));
    defparam \c0.FRAME_MATCHER_i_i31_LC_3_30_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i31_LC_3_30_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i31_LC_3_30_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i31_LC_3_30_0  (
            .in0(_gnd_net_),
            .in1(N__19569),
            .in2(_gnd_net_),
            .in3(N__33251),
            .lcout(\c0.FRAME_MATCHER_i_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49740),
            .ce(),
            .sr(N__22344));
    defparam \c0.FRAME_MATCHER_i_i30_LC_3_31_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i30_LC_3_31_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i30_LC_3_31_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i30_LC_3_31_0  (
            .in0(_gnd_net_),
            .in1(N__19299),
            .in2(_gnd_net_),
            .in3(N__33248),
            .lcout(\c0.FRAME_MATCHER_i_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49751),
            .ce(),
            .sr(N__22452));
    defparam \c0.FRAME_MATCHER_i_i21_LC_3_32_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i21_LC_3_32_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i21_LC_3_32_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i21_LC_3_32_0  (
            .in0(N__19221),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33249),
            .lcout(\c0.FRAME_MATCHER_i_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49763),
            .ce(),
            .sr(N__20769));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15321_LC_4_16_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15321_LC_4_16_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15321_LC_4_16_2 .LUT_INIT=16'b1110010010101010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15321_LC_4_16_2  (
            .in0(N__28970),
            .in1(N__17756),
            .in2(N__17709),
            .in3(N__28598),
            .lcout(\c0.n18112 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i6_LC_4_16_5 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i6_LC_4_16_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i6_LC_4_16_5 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \c0.tx2.r_Tx_Data_i6_LC_4_16_5  (
            .in0(N__17835),
            .in1(N__32423),
            .in2(N__17766),
            .in3(N__32261),
            .lcout(\c0.tx2.r_Tx_Data_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49638),
            .ce(N__24271),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i143_LC_4_17_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i143_LC_4_17_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i143_LC_4_17_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i143_LC_4_17_0  (
            .in0(N__30533),
            .in1(N__17792),
            .in2(_gnd_net_),
            .in3(N__26545),
            .lcout(data_out_frame2_17_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49630),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15400_LC_4_17_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15400_LC_4_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15400_LC_4_17_1 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_15400_LC_4_17_1  (
            .in0(N__21429),
            .in1(N__32444),
            .in2(N__22905),
            .in3(N__32147),
            .lcout(),
            .ltout(\c0.n18178_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18178_bdd_4_lut_LC_4_17_2 .C_ON=1'b0;
    defparam \c0.n18178_bdd_4_lut_LC_4_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.n18178_bdd_4_lut_LC_4_17_2 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n18178_bdd_4_lut_LC_4_17_2  (
            .in0(N__32445),
            .in1(N__22806),
            .in2(N__17853),
            .in3(N__17850),
            .lcout(\c0.n18181 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18112_bdd_4_lut_LC_4_17_3 .C_ON=1'b0;
    defparam \c0.n18112_bdd_4_lut_LC_4_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.n18112_bdd_4_lut_LC_4_17_3 .LUT_INIT=16'b1100110011100010;
    LogicCell40 \c0.n18112_bdd_4_lut_LC_4_17_3  (
            .in0(N__17829),
            .in1(N__17799),
            .in2(N__17793),
            .in3(N__28651),
            .lcout(),
            .ltout(\c0.n18115_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_6_i22_4_lut_LC_4_17_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_6_i22_4_lut_LC_4_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_6_i22_4_lut_LC_4_17_4 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_6_i22_4_lut_LC_4_17_4  (
            .in0(N__32148),
            .in1(N__17781),
            .in2(N__17769),
            .in3(N__21213),
            .lcout(\c0.n22_adj_2364 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i151_LC_4_17_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i151_LC_4_17_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i151_LC_4_17_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i151_LC_4_17_6  (
            .in0(N__29992),
            .in1(N__17757),
            .in2(_gnd_net_),
            .in3(N__26546),
            .lcout(data_out_frame2_18_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49630),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_2_i22_4_lut_LC_4_17_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_2_i22_4_lut_LC_4_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_2_i22_4_lut_LC_4_17_7 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_2_i22_4_lut_LC_4_17_7  (
            .in0(N__17745),
            .in1(N__21195),
            .in2(N__19773),
            .in3(N__32146),
            .lcout(\c0.n22_adj_2372 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_515_LC_4_18_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_515_LC_4_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_515_LC_4_18_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_515_LC_4_18_0  (
            .in0(_gnd_net_),
            .in1(N__23564),
            .in2(_gnd_net_),
            .in3(N__23523),
            .lcout(\c0.n10548 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_655_LC_4_18_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_655_LC_4_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_655_LC_4_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_655_LC_4_18_1  (
            .in0(N__23565),
            .in1(N__20395),
            .in2(_gnd_net_),
            .in3(N__23622),
            .lcout(\c0.n17249 ),
            .ltout(\c0.n17249_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i156_LC_4_18_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i156_LC_4_18_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i156_LC_4_18_2 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_frame2_0___i156_LC_4_18_2  (
            .in0(N__18117),
            .in1(N__18666),
            .in2(N__18102),
            .in3(N__18099),
            .lcout(\c0.data_out_frame2_19_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49639),
            .ce(N__26543),
            .sr(_gnd_net_));
    defparam \c0.i7_3_lut_4_lut_LC_4_18_3 .C_ON=1'b0;
    defparam \c0.i7_3_lut_4_lut_LC_4_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i7_3_lut_4_lut_LC_4_18_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_3_lut_4_lut_LC_4_18_3  (
            .in0(N__23025),
            .in1(N__18087),
            .in2(N__34325),
            .in3(N__21963),
            .lcout(\c0.n20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15151_3_lut_LC_4_18_4 .C_ON=1'b0;
    defparam \c0.i15151_3_lut_LC_4_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i15151_3_lut_LC_4_18_4 .LUT_INIT=16'b0000111100001010;
    LogicCell40 \c0.i15151_3_lut_LC_4_18_4  (
            .in0(N__29052),
            .in1(_gnd_net_),
            .in2(N__28597),
            .in3(N__34318),
            .lcout(\c0.n17678 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15004_2_lut_3_lut_LC_4_18_5 .C_ON=1'b0;
    defparam \c0.i15004_2_lut_3_lut_LC_4_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.i15004_2_lut_3_lut_LC_4_18_5 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \c0.i15004_2_lut_3_lut_LC_4_18_5  (
            .in0(N__40104),
            .in1(N__28483),
            .in2(_gnd_net_),
            .in3(N__29051),
            .lcout(\c0.n17586 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i162_LC_4_19_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i162_LC_4_19_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i162_LC_4_19_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_frame2_0___i162_LC_4_19_0  (
            .in0(N__17999),
            .in1(N__17961),
            .in2(N__20292),
            .in3(N__18867),
            .lcout(\c0.data_out_frame2_20_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49644),
            .ce(N__26518),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_615_LC_4_19_1 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_615_LC_4_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_615_LC_4_19_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_615_LC_4_19_1  (
            .in0(N__17960),
            .in1(N__17916),
            .in2(N__23772),
            .in3(N__23261),
            .lcout(),
            .ltout(\c0.n15_adj_2341_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i153_LC_4_19_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i153_LC_4_19_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i153_LC_4_19_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_frame2_0___i153_LC_4_19_2  (
            .in0(N__17898),
            .in1(N__18588),
            .in2(N__17886),
            .in3(N__23045),
            .lcout(\c0.data_out_frame2_19_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49644),
            .ce(N__26518),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_717_LC_4_19_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_717_LC_4_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_717_LC_4_19_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_717_LC_4_19_3  (
            .in0(N__17883),
            .in1(N__21571),
            .in2(_gnd_net_),
            .in3(N__23260),
            .lcout(\c0.n17234 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_596_LC_4_19_4 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_596_LC_4_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_596_LC_4_19_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_596_LC_4_19_4  (
            .in0(N__34725),
            .in1(N__23612),
            .in2(N__24003),
            .in3(N__23771),
            .lcout(),
            .ltout(\c0.n16_adj_2320_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i154_LC_4_19_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i154_LC_4_19_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i154_LC_4_19_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_frame2_0___i154_LC_4_19_5  (
            .in0(N__18675),
            .in1(N__24798),
            .in2(N__18270),
            .in3(N__18267),
            .lcout(\c0.data_out_frame2_19_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49644),
            .ce(N__26518),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i83_LC_4_20_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i83_LC_4_20_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i83_LC_4_20_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i83_LC_4_20_0  (
            .in0(N__31272),
            .in1(N__20234),
            .in2(_gnd_net_),
            .in3(N__26386),
            .lcout(data_out_frame2_10_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49650),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18058_bdd_4_lut_LC_4_20_1 .C_ON=1'b0;
    defparam \c0.n18058_bdd_4_lut_LC_4_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.n18058_bdd_4_lut_LC_4_20_1 .LUT_INIT=16'b1010101011011000;
    LogicCell40 \c0.n18058_bdd_4_lut_LC_4_20_1  (
            .in0(N__18240),
            .in1(N__18518),
            .in2(N__23563),
            .in3(N__28590),
            .lcout(\c0.n18061 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_433_LC_4_20_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_433_LC_4_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_433_LC_4_20_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_433_LC_4_20_2  (
            .in0(_gnd_net_),
            .in1(N__40093),
            .in2(_gnd_net_),
            .in3(N__20453),
            .lcout(),
            .ltout(\c0.n6_adj_2175_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_434_LC_4_20_3 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_434_LC_4_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_434_LC_4_20_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_434_LC_4_20_3  (
            .in0(N__23851),
            .in1(N__21664),
            .in2(N__18234),
            .in3(N__21896),
            .lcout(\c0.n17258 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_472_LC_4_20_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_472_LC_4_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_472_LC_4_20_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_472_LC_4_20_4  (
            .in0(_gnd_net_),
            .in1(N__18197),
            .in2(_gnd_net_),
            .in3(N__23185),
            .lcout(\c0.n17156 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i91_LC_4_20_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i91_LC_4_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i91_LC_4_20_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \c0.data_out_frame2_0___i91_LC_4_20_5  (
            .in0(N__26385),
            .in1(_gnd_net_),
            .in2(N__18206),
            .in3(N__30783),
            .lcout(data_out_frame2_11_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49650),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_LC_4_20_6 .C_ON=1'b0;
    defparam \c0.i13_4_lut_LC_4_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_LC_4_20_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i13_4_lut_LC_4_20_6  (
            .in0(N__19662),
            .in1(N__18176),
            .in2(N__18159),
            .in3(N__18144),
            .lcout(\c0.n32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i61_LC_4_21_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i61_LC_4_21_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i61_LC_4_21_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i61_LC_4_21_0  (
            .in0(N__26349),
            .in1(N__30657),
            .in2(_gnd_net_),
            .in3(N__19752),
            .lcout(data_out_frame2_7_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49655),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i149_LC_4_21_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i149_LC_4_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i149_LC_4_21_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i149_LC_4_21_1  (
            .in0(N__30109),
            .in1(N__18482),
            .in2(_gnd_net_),
            .in3(N__26351),
            .lcout(data_out_frame2_18_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49655),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i46_LC_4_21_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i46_LC_4_21_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i46_LC_4_21_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i46_LC_4_21_2  (
            .in0(N__26347),
            .in1(N__31515),
            .in2(_gnd_net_),
            .in3(N__18453),
            .lcout(data_out_frame2_5_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49655),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i60_LC_4_21_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i60_LC_4_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i60_LC_4_21_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_out_frame2_0___i60_LC_4_21_3  (
            .in0(N__18411),
            .in1(N__30709),
            .in2(_gnd_net_),
            .in3(N__26352),
            .lcout(data_out_frame2_7_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49655),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i55_LC_4_21_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i55_LC_4_21_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i55_LC_4_21_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i55_LC_4_21_4  (
            .in0(N__26348),
            .in1(N__31030),
            .in2(_gnd_net_),
            .in3(N__40864),
            .lcout(data_out_frame2_6_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49655),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i141_LC_4_21_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i141_LC_4_21_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i141_LC_4_21_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i141_LC_4_21_5  (
            .in0(N__30656),
            .in1(N__18377),
            .in2(_gnd_net_),
            .in3(N__26350),
            .lcout(data_out_frame2_17_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49655),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i144_LC_4_21_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i144_LC_4_21_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i144_LC_4_21_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i144_LC_4_21_6  (
            .in0(N__26346),
            .in1(N__30467),
            .in2(_gnd_net_),
            .in3(N__18359),
            .lcout(data_out_frame2_17_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49655),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_LC_4_21_7 .C_ON=1'b0;
    defparam \c0.i6_4_lut_LC_4_21_7 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_LC_4_21_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_LC_4_21_7  (
            .in0(N__18345),
            .in1(N__21359),
            .in2(N__18333),
            .in3(N__21962),
            .lcout(\c0.n16_adj_2170 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i54_LC_4_22_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i54_LC_4_22_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i54_LC_4_22_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i54_LC_4_22_0  (
            .in0(N__26378),
            .in1(N__31090),
            .in2(_gnd_net_),
            .in3(N__18295),
            .lcout(data_out_frame2_6_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49664),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i53_LC_4_22_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i53_LC_4_22_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i53_LC_4_22_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i53_LC_4_22_1  (
            .in0(N__31150),
            .in1(N__18787),
            .in2(_gnd_net_),
            .in3(N__26382),
            .lcout(data_out_frame2_6_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49664),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i56_LC_4_22_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i56_LC_4_22_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i56_LC_4_22_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i56_LC_4_22_2  (
            .in0(N__26379),
            .in1(N__30970),
            .in2(_gnd_net_),
            .in3(N__18649),
            .lcout(data_out_frame2_6_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49664),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i67_LC_4_22_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i67_LC_4_22_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i67_LC_4_22_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i67_LC_4_22_3  (
            .in0(N__30210),
            .in1(N__37238),
            .in2(_gnd_net_),
            .in3(N__26384),
            .lcout(data_out_frame2_8_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49664),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i51_LC_4_22_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i51_LC_4_22_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i51_LC_4_22_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i51_LC_4_22_4  (
            .in0(N__26377),
            .in1(N__31263),
            .in2(_gnd_net_),
            .in3(N__23814),
            .lcout(data_out_frame2_6_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49664),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i130_LC_4_22_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i130_LC_4_22_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i130_LC_4_22_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i130_LC_4_22_5  (
            .in0(N__30257),
            .in1(N__18617),
            .in2(_gnd_net_),
            .in3(N__26381),
            .lcout(data_out_frame2_16_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49664),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i99_LC_4_22_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i99_LC_4_22_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i99_LC_4_22_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i99_LC_4_22_6  (
            .in0(N__26380),
            .in1(N__30211),
            .in2(_gnd_net_),
            .in3(N__23902),
            .lcout(data_out_frame2_12_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49664),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i63_LC_4_22_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i63_LC_4_22_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i63_LC_4_22_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i63_LC_4_22_7  (
            .in0(N__30534),
            .in1(N__18828),
            .in2(_gnd_net_),
            .in3(N__26383),
            .lcout(data_out_frame2_7_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49664),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_610_LC_4_23_0 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_610_LC_4_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_610_LC_4_23_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_610_LC_4_23_0  (
            .in0(N__21353),
            .in1(N__18759),
            .in2(N__37252),
            .in3(N__20207),
            .lcout(\c0.n17153 ),
            .ltout(\c0.n17153_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_LC_4_23_1 .C_ON=1'b0;
    defparam \c0.i10_4_lut_LC_4_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_LC_4_23_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i10_4_lut_LC_4_23_1  (
            .in0(N__18537),
            .in1(N__18579),
            .in2(N__18573),
            .in3(N__24282),
            .lcout(\c0.n26_adj_2203 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i48_LC_4_23_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i48_LC_4_23_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i48_LC_4_23_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i48_LC_4_23_2  (
            .in0(N__26571),
            .in1(N__31399),
            .in2(_gnd_net_),
            .in3(N__18538),
            .lcout(data_out_frame2_5_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49672),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i108_LC_4_23_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i108_LC_4_23_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i108_LC_4_23_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i108_LC_4_23_3  (
            .in0(N__31618),
            .in1(N__18516),
            .in2(_gnd_net_),
            .in3(N__26573),
            .lcout(data_out_frame2_13_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49672),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_621_LC_4_23_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_621_LC_4_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_621_LC_4_23_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_621_LC_4_23_4  (
            .in0(N__18818),
            .in1(N__18780),
            .in2(_gnd_net_),
            .in3(N__24846),
            .lcout(\c0.n6_adj_2339 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i79_LC_4_23_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i79_LC_4_23_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i79_LC_4_23_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i79_LC_4_23_5  (
            .in0(N__31449),
            .in1(N__21456),
            .in2(_gnd_net_),
            .in3(N__26575),
            .lcout(data_out_frame2_9_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49672),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i96_LC_4_23_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i96_LC_4_23_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i96_LC_4_23_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i96_LC_4_23_6  (
            .in0(N__26572),
            .in1(N__30447),
            .in2(_gnd_net_),
            .in3(N__23240),
            .lcout(data_out_frame2_11_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49672),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i77_LC_4_23_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i77_LC_4_23_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i77_LC_4_23_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_out_frame2_0___i77_LC_4_23_7  (
            .in0(N__19884),
            .in1(N__31565),
            .in2(_gnd_net_),
            .in3(N__26574),
            .lcout(data_out_frame2_9_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49672),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i41_LC_4_24_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i41_LC_4_24_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i41_LC_4_24_0 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \c0.data_out_frame2_0___i41_LC_4_24_0  (
            .in0(N__26577),
            .in1(_gnd_net_),
            .in2(N__21304),
            .in3(N__30915),
            .lcout(data_out_frame2_5_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49684),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i122_LC_4_24_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i122_LC_4_24_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i122_LC_4_24_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i122_LC_4_24_1  (
            .in0(N__29810),
            .in1(N__23959),
            .in2(_gnd_net_),
            .in3(N__26579),
            .lcout(data_out_frame2_15_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49684),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i50_LC_4_24_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i50_LC_4_24_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i50_LC_4_24_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \c0.data_out_frame2_0___i50_LC_4_24_2  (
            .in0(N__26578),
            .in1(_gnd_net_),
            .in2(N__30351),
            .in3(N__23295),
            .lcout(data_out_frame2_6_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49684),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_665_LC_4_24_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_665_LC_4_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_665_LC_4_24_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_665_LC_4_24_3  (
            .in0(N__20620),
            .in1(N__21293),
            .in2(N__37254),
            .in3(N__20323),
            .lcout(\c0.n10507 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_590_LC_4_24_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_590_LC_4_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_590_LC_4_24_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_590_LC_4_24_4  (
            .in0(_gnd_net_),
            .in1(N__23667),
            .in2(_gnd_net_),
            .in3(N__18731),
            .lcout(\c0.n17273 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18046_bdd_4_lut_LC_4_24_5 .C_ON=1'b0;
    defparam \c0.n18046_bdd_4_lut_LC_4_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.n18046_bdd_4_lut_LC_4_24_5 .LUT_INIT=16'b1111101001000100;
    LogicCell40 \c0.n18046_bdd_4_lut_LC_4_24_5  (
            .in0(N__28701),
            .in1(N__37245),
            .in2(N__18951),
            .in3(N__18912),
            .lcout(\c0.n18049 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i129_LC_4_24_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i129_LC_4_24_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i129_LC_4_24_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i129_LC_4_24_6  (
            .in0(N__26576),
            .in1(N__29459),
            .in2(_gnd_net_),
            .in3(N__24915),
            .lcout(data_out_frame2_16_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49684),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_459_LC_4_24_7 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_459_LC_4_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_459_LC_4_24_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_459_LC_4_24_7  (
            .in0(N__21794),
            .in1(N__18900),
            .in2(N__18882),
            .in3(N__18873),
            .lcout(\c0.n10_adj_2190 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i0_LC_4_25_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i0_LC_4_25_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i0_LC_4_25_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i0_LC_4_25_0  (
            .in0(_gnd_net_),
            .in1(N__19119),
            .in2(_gnd_net_),
            .in3(N__33160),
            .lcout(\c0.FRAME_MATCHER_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49695),
            .ce(),
            .sr(N__22437));
    defparam \c0.i1_2_lut_3_lut_adj_663_LC_4_26_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_663_LC_4_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_663_LC_4_26_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_663_LC_4_26_0  (
            .in0(N__18983),
            .in1(N__27835),
            .in2(_gnd_net_),
            .in3(N__41863),
            .lcout(\c0.n3_adj_2282 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i5_LC_4_26_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i5_LC_4_26_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i5_LC_4_26_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i5_LC_4_26_1  (
            .in0(_gnd_net_),
            .in1(N__18966),
            .in2(_gnd_net_),
            .in3(N__33197),
            .lcout(\c0.FRAME_MATCHER_i_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49706),
            .ce(),
            .sr(N__18855));
    defparam \c0.i2_3_lut_adj_656_LC_4_26_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_656_LC_4_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_656_LC_4_26_2 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.i2_3_lut_adj_656_LC_4_26_2  (
            .in0(N__18981),
            .in1(N__19038),
            .in2(_gnd_net_),
            .in3(N__19074),
            .lcout(\c0.n15164 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_552_LC_4_26_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_552_LC_4_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_552_LC_4_26_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i1_2_lut_adj_552_LC_4_26_3  (
            .in0(N__41861),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18982),
            .lcout(\c0.n43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_219_Select_3_i3_2_lut_3_lut_LC_4_26_4 .C_ON=1'b0;
    defparam \c0.select_219_Select_3_i3_2_lut_3_lut_LC_4_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.select_219_Select_3_i3_2_lut_3_lut_LC_4_26_4 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \c0.select_219_Select_3_i3_2_lut_3_lut_LC_4_26_4  (
            .in0(N__27839),
            .in1(N__19075),
            .in2(_gnd_net_),
            .in3(N__41864),
            .lcout(\c0.n3_adj_2227 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_219_Select_4_i3_2_lut_3_lut_LC_4_26_5 .C_ON=1'b0;
    defparam \c0.select_219_Select_4_i3_2_lut_3_lut_LC_4_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.select_219_Select_4_i3_2_lut_3_lut_LC_4_26_5 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \c0.select_219_Select_4_i3_2_lut_3_lut_LC_4_26_5  (
            .in0(N__41865),
            .in1(_gnd_net_),
            .in2(N__27843),
            .in3(N__19040),
            .lcout(\c0.n3_adj_2179 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_407_LC_4_26_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_407_LC_4_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_407_LC_4_26_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_407_LC_4_26_6  (
            .in0(_gnd_net_),
            .in1(N__19039),
            .in2(_gnd_net_),
            .in3(N__41860),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_750_LC_4_26_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_750_LC_4_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_750_LC_4_26_7 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \c0.i1_2_lut_adj_750_LC_4_26_7  (
            .in0(N__41862),
            .in1(N__19079),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_2_lut_LC_4_27_0 .C_ON=1'b1;
    defparam \c0.add_977_2_lut_LC_4_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_2_lut_LC_4_27_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_977_2_lut_LC_4_27_0  (
            .in0(N__27048),
            .in1(N__37155),
            .in2(N__19545),
            .in3(N__19110),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_0 ),
            .ltout(),
            .carryin(bfn_4_27_0_),
            .carryout(\c0.n16079 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_3_lut_LC_4_27_1 .C_ON=1'b1;
    defparam \c0.add_977_3_lut_LC_4_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_3_lut_LC_4_27_1 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \c0.add_977_3_lut_LC_4_27_1  (
            .in0(N__25377),
            .in1(N__19494),
            .in2(N__32872),
            .in3(N__19095),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_1 ),
            .ltout(),
            .carryin(\c0.n16079 ),
            .carryout(\c0.n16080 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_4_lut_LC_4_27_2 .C_ON=1'b1;
    defparam \c0.add_977_4_lut_LC_4_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_4_lut_LC_4_27_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_977_4_lut_LC_4_27_2  (
            .in0(N__22332),
            .in1(N__37088),
            .in2(N__19546),
            .in3(N__19092),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_2 ),
            .ltout(),
            .carryin(\c0.n16080 ),
            .carryout(\c0.n16081 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_5_lut_LC_4_27_3 .C_ON=1'b1;
    defparam \c0.add_977_5_lut_LC_4_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_5_lut_LC_4_27_3 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \c0.add_977_5_lut_LC_4_27_3  (
            .in0(N__19089),
            .in1(N__19498),
            .in2(N__19083),
            .in3(N__19050),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_3 ),
            .ltout(),
            .carryin(\c0.n16081 ),
            .carryout(\c0.n16082 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_6_lut_LC_4_27_4 .C_ON=1'b1;
    defparam \c0.add_977_6_lut_LC_4_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_6_lut_LC_4_27_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_977_6_lut_LC_4_27_4  (
            .in0(N__19047),
            .in1(N__19041),
            .in2(N__19547),
            .in3(N__18996),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_4 ),
            .ltout(),
            .carryin(\c0.n16082 ),
            .carryout(\c0.n16083 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_7_lut_LC_4_27_5 .C_ON=1'b1;
    defparam \c0.add_977_7_lut_LC_4_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_7_lut_LC_4_27_5 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \c0.add_977_7_lut_LC_4_27_5  (
            .in0(N__18993),
            .in1(N__19502),
            .in2(N__18987),
            .in3(N__18960),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_5 ),
            .ltout(),
            .carryin(\c0.n16083 ),
            .carryout(\c0.n16084 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_8_lut_LC_4_27_6 .C_ON=1'b1;
    defparam \c0.add_977_8_lut_LC_4_27_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_8_lut_LC_4_27_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_977_8_lut_LC_4_27_6  (
            .in0(N__20862),
            .in1(N__20880),
            .in2(N__19548),
            .in3(N__19200),
            .lcout(\c0.n3 ),
            .ltout(),
            .carryin(\c0.n16084 ),
            .carryout(\c0.n16085 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_9_lut_LC_4_27_7 .C_ON=1'b1;
    defparam \c0.add_977_9_lut_LC_4_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_9_lut_LC_4_27_7 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \c0.add_977_9_lut_LC_4_27_7  (
            .in0(N__27063),
            .in1(N__19506),
            .in2(N__27095),
            .in3(N__19191),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_7 ),
            .ltout(),
            .carryin(\c0.n16085 ),
            .carryout(\c0.n16086 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_10_lut_LC_4_28_0 .C_ON=1'b1;
    defparam \c0.add_977_10_lut_LC_4_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_10_lut_LC_4_28_0 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \c0.add_977_10_lut_LC_4_28_0  (
            .in0(N__20892),
            .in1(N__19507),
            .in2(N__22192),
            .in3(N__19176),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_8 ),
            .ltout(),
            .carryin(bfn_4_28_0_),
            .carryout(\c0.n16087 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_11_lut_LC_4_28_1 .C_ON=1'b1;
    defparam \c0.add_977_11_lut_LC_4_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_11_lut_LC_4_28_1 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_977_11_lut_LC_4_28_1  (
            .in0(N__20886),
            .in1(N__22632),
            .in2(N__19549),
            .in3(N__19173),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_9 ),
            .ltout(),
            .carryin(\c0.n16087 ),
            .carryout(\c0.n16088 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_12_lut_LC_4_28_2 .C_ON=1'b1;
    defparam \c0.add_977_12_lut_LC_4_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_12_lut_LC_4_28_2 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \c0.add_977_12_lut_LC_4_28_2  (
            .in0(N__27969),
            .in1(N__19511),
            .in2(N__28005),
            .in3(N__19170),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_10 ),
            .ltout(),
            .carryin(\c0.n16088 ),
            .carryout(\c0.n16089 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_13_lut_LC_4_28_3 .C_ON=1'b1;
    defparam \c0.add_977_13_lut_LC_4_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_13_lut_LC_4_28_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_977_13_lut_LC_4_28_3  (
            .in0(N__27114),
            .in1(N__27158),
            .in2(N__19550),
            .in3(N__19155),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_11 ),
            .ltout(),
            .carryin(\c0.n16089 ),
            .carryout(\c0.n16090 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_14_lut_LC_4_28_4 .C_ON=1'b1;
    defparam \c0.add_977_14_lut_LC_4_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_14_lut_LC_4_28_4 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \c0.add_977_14_lut_LC_4_28_4  (
            .in0(N__19152),
            .in1(N__19515),
            .in2(N__25872),
            .in3(N__19146),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_12 ),
            .ltout(),
            .carryin(\c0.n16090 ),
            .carryout(\c0.n16091 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_15_lut_LC_4_28_5 .C_ON=1'b1;
    defparam \c0.add_977_15_lut_LC_4_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_15_lut_LC_4_28_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_977_15_lut_LC_4_28_5  (
            .in0(N__27174),
            .in1(N__27202),
            .in2(N__19551),
            .in3(N__19134),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_13 ),
            .ltout(),
            .carryin(\c0.n16091 ),
            .carryout(\c0.n16092 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_16_lut_LC_4_28_6 .C_ON=1'b1;
    defparam \c0.add_977_16_lut_LC_4_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_16_lut_LC_4_28_6 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \c0.add_977_16_lut_LC_4_28_6  (
            .in0(N__27900),
            .in1(N__19519),
            .in2(N__27941),
            .in3(N__19278),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_14 ),
            .ltout(),
            .carryin(\c0.n16092 ),
            .carryout(\c0.n16093 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_17_lut_LC_4_28_7 .C_ON=1'b1;
    defparam \c0.add_977_17_lut_LC_4_28_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_17_lut_LC_4_28_7 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_977_17_lut_LC_4_28_7  (
            .in0(N__27222),
            .in1(N__27263),
            .in2(N__19552),
            .in3(N__19263),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_15 ),
            .ltout(),
            .carryin(\c0.n16093 ),
            .carryout(\c0.n16094 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_18_lut_LC_4_29_0 .C_ON=1'b1;
    defparam \c0.add_977_18_lut_LC_4_29_0 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_18_lut_LC_4_29_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_977_18_lut_LC_4_29_0  (
            .in0(N__24954),
            .in1(N__27891),
            .in2(N__19553),
            .in3(N__19260),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_16 ),
            .ltout(),
            .carryin(bfn_4_29_0_),
            .carryout(\c0.n16095 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_19_lut_LC_4_29_1 .C_ON=1'b1;
    defparam \c0.add_977_19_lut_LC_4_29_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_19_lut_LC_4_29_1 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_977_19_lut_LC_4_29_1  (
            .in0(N__20781),
            .in1(N__20799),
            .in2(N__19557),
            .in3(N__19257),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_17 ),
            .ltout(),
            .carryin(\c0.n16095 ),
            .carryout(\c0.n16096 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_20_lut_LC_4_29_2 .C_ON=1'b1;
    defparam \c0.add_977_20_lut_LC_4_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_20_lut_LC_4_29_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_977_20_lut_LC_4_29_2  (
            .in0(N__25404),
            .in1(N__25432),
            .in2(N__19554),
            .in3(N__19254),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_18 ),
            .ltout(),
            .carryin(\c0.n16096 ),
            .carryout(\c0.n16097 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_21_lut_LC_4_29_3 .C_ON=1'b1;
    defparam \c0.add_977_21_lut_LC_4_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_21_lut_LC_4_29_3 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \c0.add_977_21_lut_LC_4_29_3  (
            .in0(N__24969),
            .in1(N__19529),
            .in2(N__25008),
            .in3(N__19239),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_19 ),
            .ltout(),
            .carryin(\c0.n16097 ),
            .carryout(\c0.n16098 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_22_lut_LC_4_29_4 .C_ON=1'b1;
    defparam \c0.add_977_22_lut_LC_4_29_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_22_lut_LC_4_29_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_977_22_lut_LC_4_29_4  (
            .in0(N__25020),
            .in1(N__25059),
            .in2(N__19555),
            .in3(N__19224),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_20 ),
            .ltout(),
            .carryin(\c0.n16098 ),
            .carryout(\c0.n16099 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_23_lut_LC_4_29_5 .C_ON=1'b1;
    defparam \c0.add_977_23_lut_LC_4_29_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_23_lut_LC_4_29_5 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \c0.add_977_23_lut_LC_4_29_5  (
            .in0(N__20919),
            .in1(N__19533),
            .in2(N__20952),
            .in3(N__19212),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_21 ),
            .ltout(),
            .carryin(\c0.n16099 ),
            .carryout(\c0.n16100 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_24_lut_LC_4_29_6 .C_ON=1'b1;
    defparam \c0.add_977_24_lut_LC_4_29_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_24_lut_LC_4_29_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_977_24_lut_LC_4_29_6  (
            .in0(N__25311),
            .in1(N__25327),
            .in2(N__19556),
            .in3(N__19203),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_22 ),
            .ltout(),
            .carryin(\c0.n16100 ),
            .carryout(\c0.n16101 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_25_lut_LC_4_29_7 .C_ON=1'b1;
    defparam \c0.add_977_25_lut_LC_4_29_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_25_lut_LC_4_29_7 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \c0.add_977_25_lut_LC_4_29_7  (
            .in0(N__25074),
            .in1(N__19537),
            .in2(N__25124),
            .in3(N__19374),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_23 ),
            .ltout(),
            .carryin(\c0.n16101 ),
            .carryout(\c0.n16102 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_26_lut_LC_4_30_0 .C_ON=1'b1;
    defparam \c0.add_977_26_lut_LC_4_30_0 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_26_lut_LC_4_30_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_977_26_lut_LC_4_30_0  (
            .in0(N__25140),
            .in1(N__25170),
            .in2(N__19541),
            .in3(N__19371),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_24 ),
            .ltout(),
            .carryin(bfn_4_30_0_),
            .carryout(\c0.n16103 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_27_lut_LC_4_30_1 .C_ON=1'b1;
    defparam \c0.add_977_27_lut_LC_4_30_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_27_lut_LC_4_30_1 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \c0.add_977_27_lut_LC_4_30_1  (
            .in0(N__25182),
            .in1(N__19478),
            .in2(N__25221),
            .in3(N__19368),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_25 ),
            .ltout(),
            .carryin(\c0.n16103 ),
            .carryout(\c0.n16104 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_28_lut_LC_4_30_2 .C_ON=1'b1;
    defparam \c0.add_977_28_lut_LC_4_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_28_lut_LC_4_30_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_977_28_lut_LC_4_30_2  (
            .in0(N__25233),
            .in1(N__25281),
            .in2(N__19542),
            .in3(N__19365),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_26 ),
            .ltout(),
            .carryin(\c0.n16104 ),
            .carryout(\c0.n16105 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_29_lut_LC_4_30_3 .C_ON=1'b1;
    defparam \c0.add_977_29_lut_LC_4_30_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_29_lut_LC_4_30_3 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \c0.add_977_29_lut_LC_4_30_3  (
            .in0(N__20913),
            .in1(N__19482),
            .in2(N__22698),
            .in3(N__19362),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_27 ),
            .ltout(),
            .carryin(\c0.n16105 ),
            .carryout(\c0.n16106 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_30_lut_LC_4_30_4 .C_ON=1'b1;
    defparam \c0.add_977_30_lut_LC_4_30_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_30_lut_LC_4_30_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_977_30_lut_LC_4_30_4  (
            .in0(N__26997),
            .in1(N__27024),
            .in2(N__19543),
            .in3(N__19350),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_28 ),
            .ltout(),
            .carryin(\c0.n16106 ),
            .carryout(\c0.n16107 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_31_lut_LC_4_30_5 .C_ON=1'b1;
    defparam \c0.add_977_31_lut_LC_4_30_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_31_lut_LC_4_30_5 .LUT_INIT=16'b1000101110111000;
    LogicCell40 \c0.add_977_31_lut_LC_4_30_5  (
            .in0(N__19347),
            .in1(N__19486),
            .in2(N__19335),
            .in3(N__19302),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_29 ),
            .ltout(),
            .carryin(\c0.n16107 ),
            .carryout(\c0.n16108 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_32_lut_LC_4_30_6 .C_ON=1'b1;
    defparam \c0.add_977_32_lut_LC_4_30_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_32_lut_LC_4_30_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.add_977_32_lut_LC_4_30_6  (
            .in0(N__33618),
            .in1(N__33651),
            .in2(N__19544),
            .in3(N__19293),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_30 ),
            .ltout(),
            .carryin(\c0.n16108 ),
            .carryout(\c0.n16109 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_977_33_lut_LC_4_30_7 .C_ON=1'b0;
    defparam \c0.add_977_33_lut_LC_4_30_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_977_33_lut_LC_4_30_7 .LUT_INIT=16'b1101000111100010;
    LogicCell40 \c0.add_977_33_lut_LC_4_30_7  (
            .in0(N__29542),
            .in1(N__19490),
            .in2(N__21039),
            .in3(N__19290),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1278_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Bit_Index_i0_LC_4_31_0 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_i0_LC_4_31_0 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Bit_Index_i0_LC_4_31_0 .LUT_INIT=16'b1001100100000000;
    LogicCell40 \c0.rx.r_Bit_Index_i0_LC_4_31_0  (
            .in0(N__37852),
            .in1(N__25624),
            .in2(_gnd_net_),
            .in3(N__21119),
            .lcout(r_Bit_Index_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49764),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2593_2_lut_LC_4_31_1 .C_ON=1'b0;
    defparam \c0.rx.i2593_2_lut_LC_4_31_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2593_2_lut_LC_4_31_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.rx.i2593_2_lut_LC_4_31_1  (
            .in0(_gnd_net_),
            .in1(N__37851),
            .in2(_gnd_net_),
            .in3(N__37933),
            .lcout(n5244),
            .ltout(n5244_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i14631_3_lut_4_lut_LC_4_31_2 .C_ON=1'b0;
    defparam \c0.rx.i14631_3_lut_4_lut_LC_4_31_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i14631_3_lut_4_lut_LC_4_31_2 .LUT_INIT=16'b1111111100101010;
    LogicCell40 \c0.rx.i14631_3_lut_4_lut_LC_4_31_2  (
            .in0(N__25544),
            .in1(N__37902),
            .in2(N__19563),
            .in3(N__25623),
            .lcout(n11018),
            .ltout(n11018_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Bit_Index_i1_LC_4_31_3 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_i1_LC_4_31_3 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Bit_Index_i1_LC_4_31_3 .LUT_INIT=16'b1011000001000000;
    LogicCell40 \c0.rx.r_Bit_Index_i1_LC_4_31_3  (
            .in0(N__25625),
            .in1(N__37853),
            .in2(N__19560),
            .in3(N__37934),
            .lcout(r_Bit_Index_1_adj_2436),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49764),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i15231_1_lut_LC_4_31_4 .C_ON=1'b0;
    defparam \c0.rx.i15231_1_lut_LC_4_31_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i15231_1_lut_LC_4_31_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \c0.rx.i15231_1_lut_LC_4_31_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39016),
            .lcout(\c0.n18008 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i15224_2_lut_3_lut_LC_4_31_5 .C_ON=1'b0;
    defparam \c0.rx.i15224_2_lut_3_lut_LC_4_31_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i15224_2_lut_3_lut_LC_4_31_5 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \c0.rx.i15224_2_lut_3_lut_LC_4_31_5  (
            .in0(N__25484),
            .in1(N__25545),
            .in2(_gnd_net_),
            .in3(N__31851),
            .lcout(\c0.rx.n17058 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_2__I_0_56_Mux_0_i2_3_lut_4_lut_LC_4_31_6 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_2__I_0_56_Mux_0_i2_3_lut_4_lut_LC_4_31_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_SM_Main_2__I_0_56_Mux_0_i2_3_lut_4_lut_LC_4_31_6 .LUT_INIT=16'b1111000001111111;
    LogicCell40 \c0.rx.r_SM_Main_2__I_0_56_Mux_0_i2_3_lut_4_lut_LC_4_31_6  (
            .in0(N__21131),
            .in1(N__37903),
            .in2(N__25602),
            .in3(N__25485),
            .lcout(),
            .ltout(n13692_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_i0_LC_4_31_7 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_i0_LC_4_31_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_SM_Main_i0_LC_4_31_7 .LUT_INIT=16'b0001010100000100;
    LogicCell40 \c0.rx.r_SM_Main_i0_LC_4_31_7  (
            .in0(N__31852),
            .in1(N__25546),
            .in2(N__19392),
            .in3(N__21009),
            .lcout(\c0.rx.r_SM_Main_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49764),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Clock_Count__i0_LC_4_32_0 .C_ON=1'b1;
    defparam \c0.rx.r_Clock_Count__i0_LC_4_32_0 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i0_LC_4_32_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.r_Clock_Count__i0_LC_4_32_0  (
            .in0(_gnd_net_),
            .in1(N__22559),
            .in2(_gnd_net_),
            .in3(N__19389),
            .lcout(\c0.rx.r_Clock_Count_0 ),
            .ltout(),
            .carryin(bfn_4_32_0_),
            .carryout(\c0.rx.n16125 ),
            .clk(N__49776),
            .ce(N__20979),
            .sr(N__21018));
    defparam \c0.rx.r_Clock_Count__i1_LC_4_32_1 .C_ON=1'b1;
    defparam \c0.rx.r_Clock_Count__i1_LC_4_32_1 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i1_LC_4_32_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.r_Clock_Count__i1_LC_4_32_1  (
            .in0(_gnd_net_),
            .in1(N__20991),
            .in2(_gnd_net_),
            .in3(N__19608),
            .lcout(\c0.rx.r_Clock_Count_1 ),
            .ltout(),
            .carryin(\c0.rx.n16125 ),
            .carryout(\c0.rx.n16126 ),
            .clk(N__49776),
            .ce(N__20979),
            .sr(N__21018));
    defparam \c0.rx.r_Clock_Count__i2_LC_4_32_2 .C_ON=1'b1;
    defparam \c0.rx.r_Clock_Count__i2_LC_4_32_2 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i2_LC_4_32_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.r_Clock_Count__i2_LC_4_32_2  (
            .in0(_gnd_net_),
            .in1(N__22574),
            .in2(_gnd_net_),
            .in3(N__19605),
            .lcout(\c0.rx.r_Clock_Count_2 ),
            .ltout(),
            .carryin(\c0.rx.n16126 ),
            .carryout(\c0.rx.n16127 ),
            .clk(N__49776),
            .ce(N__20979),
            .sr(N__21018));
    defparam \c0.rx.r_Clock_Count__i3_LC_4_32_3 .C_ON=1'b1;
    defparam \c0.rx.r_Clock_Count__i3_LC_4_32_3 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i3_LC_4_32_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.r_Clock_Count__i3_LC_4_32_3  (
            .in0(_gnd_net_),
            .in1(N__22541),
            .in2(_gnd_net_),
            .in3(N__19602),
            .lcout(\c0.rx.r_Clock_Count_3 ),
            .ltout(),
            .carryin(\c0.rx.n16127 ),
            .carryout(\c0.rx.n16128 ),
            .clk(N__49776),
            .ce(N__20979),
            .sr(N__21018));
    defparam \c0.rx.r_Clock_Count__i4_LC_4_32_4 .C_ON=1'b1;
    defparam \c0.rx.r_Clock_Count__i4_LC_4_32_4 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i4_LC_4_32_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.r_Clock_Count__i4_LC_4_32_4  (
            .in0(_gnd_net_),
            .in1(N__21003),
            .in2(_gnd_net_),
            .in3(N__19599),
            .lcout(\c0.rx.r_Clock_Count_4 ),
            .ltout(),
            .carryin(\c0.rx.n16128 ),
            .carryout(\c0.rx.n16129 ),
            .clk(N__49776),
            .ce(N__20979),
            .sr(N__21018));
    defparam \c0.rx.r_Clock_Count__i5_LC_4_32_5 .C_ON=1'b1;
    defparam \c0.rx.r_Clock_Count__i5_LC_4_32_5 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i5_LC_4_32_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.r_Clock_Count__i5_LC_4_32_5  (
            .in0(_gnd_net_),
            .in1(N__31933),
            .in2(_gnd_net_),
            .in3(N__19596),
            .lcout(\c0.rx.r_Clock_Count_5 ),
            .ltout(),
            .carryin(\c0.rx.n16129 ),
            .carryout(\c0.rx.n16130 ),
            .clk(N__49776),
            .ce(N__20979),
            .sr(N__21018));
    defparam \c0.rx.r_Clock_Count__i6_LC_4_32_6 .C_ON=1'b1;
    defparam \c0.rx.r_Clock_Count__i6_LC_4_32_6 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i6_LC_4_32_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.r_Clock_Count__i6_LC_4_32_6  (
            .in0(_gnd_net_),
            .in1(N__31726),
            .in2(_gnd_net_),
            .in3(N__19593),
            .lcout(\c0.rx.r_Clock_Count_6 ),
            .ltout(),
            .carryin(\c0.rx.n16130 ),
            .carryout(\c0.rx.n16131 ),
            .clk(N__49776),
            .ce(N__20979),
            .sr(N__21018));
    defparam \c0.rx.r_Clock_Count__i7_LC_4_32_7 .C_ON=1'b0;
    defparam \c0.rx.r_Clock_Count__i7_LC_4_32_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Clock_Count__i7_LC_4_32_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.rx.r_Clock_Count__i7_LC_4_32_7  (
            .in0(_gnd_net_),
            .in1(N__31767),
            .in2(_gnd_net_),
            .in3(N__19590),
            .lcout(\c0.rx.r_Clock_Count_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49776),
            .ce(N__20979),
            .sr(N__21018));
    defparam \c0.data_out_frame2_0___i146_LC_5_14_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i146_LC_5_14_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i146_LC_5_14_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i146_LC_5_14_0  (
            .in0(N__30264),
            .in1(N__19586),
            .in2(_gnd_net_),
            .in3(N__26517),
            .lcout(data_out_frame2_18_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49656),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_i7_LC_5_16_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_i7_LC_5_16_0 .SEQ_MODE=4'b1001;
    defparam \c0.byte_transmit_counter2_i7_LC_5_16_0 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \c0.byte_transmit_counter2_i7_LC_5_16_0  (
            .in0(N__26664),
            .in1(N__39702),
            .in2(N__34477),
            .in3(N__42095),
            .lcout(\c0.byte_transmit_counter2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49645),
            .ce(),
            .sr(N__32043));
    defparam \c0.i5_3_lut_4_lut_adj_690_LC_5_17_0 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_adj_690_LC_5_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_adj_690_LC_5_17_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_adj_690_LC_5_17_0  (
            .in0(N__19830),
            .in1(N__21524),
            .in2(N__19971),
            .in3(N__19904),
            .lcout(),
            .ltout(\c0.n14_adj_2188_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i163_LC_5_17_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i163_LC_5_17_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i163_LC_5_17_1 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_frame2_0___i163_LC_5_17_1  (
            .in0(N__20043),
            .in1(N__19722),
            .in2(N__19791),
            .in3(N__19788),
            .lcout(\c0.data_out_frame2_20_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49634),
            .ce(N__26544),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_447_LC_5_17_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_447_LC_5_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_447_LC_5_17_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_447_LC_5_17_2  (
            .in0(_gnd_net_),
            .in1(N__40290),
            .in2(_gnd_net_),
            .in3(N__23999),
            .lcout(\c0.n17294 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_470_LC_5_17_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_470_LC_5_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_470_LC_5_17_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_470_LC_5_17_3  (
            .in0(N__40673),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19764),
            .lcout(\c0.n17240 ),
            .ltout(\c0.n17240_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i161_LC_5_17_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i161_LC_5_17_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i161_LC_5_17_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_frame2_0___i161_LC_5_17_4  (
            .in0(N__20478),
            .in1(N__20265),
            .in2(N__19716),
            .in3(N__19713),
            .lcout(\c0.data_out_frame2_20_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49634),
            .ce(N__26544),
            .sr(_gnd_net_));
    defparam \c0.i15015_3_lut_LC_5_17_6 .C_ON=1'b0;
    defparam \c0.i15015_3_lut_LC_5_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.i15015_3_lut_LC_5_17_6 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \c0.i15015_3_lut_LC_5_17_6  (
            .in0(N__28648),
            .in1(N__40672),
            .in2(_gnd_net_),
            .in3(N__28972),
            .lcout(\c0.n17603 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14662_3_lut_LC_5_17_7 .C_ON=1'b0;
    defparam \c0.i14662_3_lut_LC_5_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.i14662_3_lut_LC_5_17_7 .LUT_INIT=16'b1010101001000100;
    LogicCell40 \c0.i14662_3_lut_LC_5_17_7  (
            .in0(N__28971),
            .in1(N__37636),
            .in2(_gnd_net_),
            .in3(N__28647),
            .lcout(\c0.n17439 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i158_LC_5_18_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i158_LC_5_18_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i158_LC_5_18_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_frame2_0___i158_LC_5_18_0  (
            .in0(N__19977),
            .in1(N__19614),
            .in2(N__19686),
            .in3(N__20138),
            .lcout(\c0.data_out_frame2_19_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49646),
            .ce(N__26542),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_531_LC_5_18_1 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_531_LC_5_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_531_LC_5_18_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_531_LC_5_18_1  (
            .in0(N__19836),
            .in1(N__19661),
            .in2(N__19631),
            .in3(N__24845),
            .lcout(\c0.n15_adj_2291 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_710_LC_5_18_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_710_LC_5_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_710_LC_5_18_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_710_LC_5_18_2  (
            .in0(N__24080),
            .in1(N__26645),
            .in2(N__23922),
            .in3(N__41107),
            .lcout(\c0.n17288 ),
            .ltout(\c0.n17288_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_adj_671_LC_5_18_3 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_adj_671_LC_5_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_adj_671_LC_5_18_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_adj_671_LC_5_18_3  (
            .in0(N__23381),
            .in1(N__20034),
            .in2(N__19980),
            .in3(N__26055),
            .lcout(\c0.n14_adj_2292 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_523_LC_5_18_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_523_LC_5_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_523_LC_5_18_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_523_LC_5_18_5  (
            .in0(N__26646),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24081),
            .lcout(),
            .ltout(\c0.n10428_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i164_LC_5_18_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i164_LC_5_18_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i164_LC_5_18_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_frame2_0___i164_LC_5_18_6  (
            .in0(N__19970),
            .in1(N__20624),
            .in2(N__19956),
            .in3(N__19953),
            .lcout(\c0.data_out_frame2_20_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49646),
            .ce(N__26542),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_522_LC_5_18_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_522_LC_5_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_522_LC_5_18_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_522_LC_5_18_7  (
            .in0(N__41106),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23918),
            .lcout(\c0.n10504 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i90_LC_5_19_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i90_LC_5_19_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i90_LC_5_19_0 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \c0.data_out_frame2_0___i90_LC_5_19_0  (
            .in0(_gnd_net_),
            .in1(N__26415),
            .in2(N__20080),
            .in3(N__29812),
            .lcout(data_out_frame2_11_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49651),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i138_LC_5_19_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i138_LC_5_19_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i138_LC_5_19_1 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \c0.data_out_frame2_0___i138_LC_5_19_1  (
            .in0(N__29811),
            .in1(N__19922),
            .in2(N__26547),
            .in3(_gnd_net_),
            .lcout(data_out_frame2_17_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49651),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18208_bdd_4_lut_LC_5_19_2 .C_ON=1'b0;
    defparam \c0.n18208_bdd_4_lut_LC_5_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.n18208_bdd_4_lut_LC_5_19_2 .LUT_INIT=16'b1111101001000100;
    LogicCell40 \c0.n18208_bdd_4_lut_LC_5_19_2  (
            .in0(N__28649),
            .in1(N__24380),
            .in2(N__19903),
            .in3(N__21687),
            .lcout(\c0.n17568 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_529_LC_5_19_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_529_LC_5_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_529_LC_5_19_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_529_LC_5_19_3  (
            .in0(_gnd_net_),
            .in1(N__21311),
            .in2(_gnd_net_),
            .in3(N__20521),
            .lcout(\c0.n10554 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_486_LC_5_19_4 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_486_LC_5_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_486_LC_5_19_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_486_LC_5_19_4  (
            .in0(N__20288),
            .in1(N__20183),
            .in2(N__24555),
            .in3(N__20431),
            .lcout(\c0.n15_adj_2205 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_3_i6_4_lut_LC_5_19_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_3_i6_4_lut_LC_5_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_3_i6_4_lut_LC_5_19_5 .LUT_INIT=16'b1011100010001000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_3_i6_4_lut_LC_5_19_5  (
            .in0(N__20256),
            .in1(N__28650),
            .in2(N__23522),
            .in3(N__29053),
            .lcout(\c0.n6_adj_2139 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_609_LC_5_19_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_609_LC_5_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_609_LC_5_19_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_609_LC_5_19_6  (
            .in0(N__23602),
            .in1(N__20106),
            .in2(_gnd_net_),
            .in3(N__20229),
            .lcout(\c0.n10492 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_714_LC_5_19_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_714_LC_5_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_714_LC_5_19_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_714_LC_5_19_7  (
            .in0(N__20182),
            .in1(N__23744),
            .in2(_gnd_net_),
            .in3(N__21752),
            .lcout(\c0.n17255 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i133_LC_5_20_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i133_LC_5_20_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i133_LC_5_20_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_out_frame2_0___i133_LC_5_20_0  (
            .in0(N__30105),
            .in1(N__26363),
            .in2(_gnd_net_),
            .in3(N__20113),
            .lcout(data_out_frame2_16_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49657),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i98_LC_5_20_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i98_LC_5_20_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i98_LC_5_20_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \c0.data_out_frame2_0___i98_LC_5_20_1  (
            .in0(N__26361),
            .in1(_gnd_net_),
            .in2(N__30274),
            .in3(N__23613),
            .lcout(data_out_frame2_12_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49657),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i94_LC_5_20_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i94_LC_5_20_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i94_LC_5_20_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_out_frame2_0___i94_LC_5_20_2  (
            .in0(N__30594),
            .in1(N__26364),
            .in2(_gnd_net_),
            .in3(N__21866),
            .lcout(data_out_frame2_11_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49657),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i93_LC_5_20_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i93_LC_5_20_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i93_LC_5_20_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i93_LC_5_20_3  (
            .in0(N__26360),
            .in1(N__30646),
            .in2(_gnd_net_),
            .in3(N__21897),
            .lcout(data_out_frame2_11_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49657),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_445_LC_5_20_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_445_LC_5_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_445_LC_5_20_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_445_LC_5_20_4  (
            .in0(N__20064),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24744),
            .lcout(),
            .ltout(\c0.n6_adj_2182_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_446_LC_5_20_5 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_446_LC_5_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_446_LC_5_20_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_446_LC_5_20_5  (
            .in0(N__21745),
            .in1(N__20474),
            .in2(N__20463),
            .in3(N__24036),
            .lcout(\c0.n10229 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i103_LC_5_20_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i103_LC_5_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i103_LC_5_20_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_out_frame2_0___i103_LC_5_20_6  (
            .in0(N__29991),
            .in1(N__26362),
            .in2(_gnd_net_),
            .in3(N__22962),
            .lcout(data_out_frame2_12_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49657),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i68_LC_5_20_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i68_LC_5_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i68_LC_5_20_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i68_LC_5_20_7  (
            .in0(N__26359),
            .in1(N__30158),
            .in2(_gnd_net_),
            .in3(N__24832),
            .lcout(data_out_frame2_8_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49657),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i76_LC_5_21_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i76_LC_5_21_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i76_LC_5_21_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_out_frame2_0___i76_LC_5_21_0  (
            .in0(N__24636),
            .in1(N__31623),
            .in2(_gnd_net_),
            .in3(N__26337),
            .lcout(data_out_frame2_9_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49665),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_4_lut_LC_5_21_1 .C_ON=1'b0;
    defparam \c0.i3_4_lut_4_lut_LC_5_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_4_lut_LC_5_21_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \c0.i3_4_lut_4_lut_LC_5_21_1  (
            .in0(N__40248),
            .in1(N__36092),
            .in2(N__33687),
            .in3(N__39758),
            .lcout(n10725),
            .ltout(n10725_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i104_LC_5_21_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i104_LC_5_21_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i104_LC_5_21_2 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \c0.data_out_frame2_0___i104_LC_5_21_2  (
            .in0(_gnd_net_),
            .in1(N__29916),
            .in2(N__20442),
            .in3(N__20424),
            .lcout(data_out_frame2_12_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49665),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i84_LC_5_21_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i84_LC_5_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i84_LC_5_21_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i84_LC_5_21_3  (
            .in0(N__26335),
            .in1(N__31194),
            .in2(_gnd_net_),
            .in3(N__20379),
            .lcout(data_out_frame2_10_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49665),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15316_LC_5_21_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15316_LC_5_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15316_LC_5_21_4 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15316_LC_5_21_4  (
            .in0(N__28641),
            .in1(N__28959),
            .in2(N__24073),
            .in3(N__21868),
            .lcout(\c0.n18106 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i131_LC_5_21_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i131_LC_5_21_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i131_LC_5_21_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i131_LC_5_21_5  (
            .in0(N__26334),
            .in1(N__30215),
            .in2(_gnd_net_),
            .in3(N__20322),
            .lcout(data_out_frame2_16_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49665),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i123_LC_5_21_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i123_LC_5_21_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i123_LC_5_21_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i123_LC_5_21_6  (
            .in0(N__30780),
            .in1(N__20612),
            .in2(_gnd_net_),
            .in3(N__26336),
            .lcout(data_out_frame2_15_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49665),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i124_LC_5_21_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i124_LC_5_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i124_LC_5_21_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i124_LC_5_21_7  (
            .in0(N__26333),
            .in1(N__30708),
            .in2(_gnd_net_),
            .in3(N__24422),
            .lcout(data_out_frame2_15_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49665),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i137_LC_5_22_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i137_LC_5_22_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i137_LC_5_22_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_out_frame2_0___i137_LC_5_22_0  (
            .in0(N__29861),
            .in1(N__26343),
            .in2(_gnd_net_),
            .in3(N__21713),
            .lcout(data_out_frame2_17_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49673),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i147_LC_5_22_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i147_LC_5_22_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i147_LC_5_22_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i147_LC_5_22_1  (
            .in0(N__26340),
            .in1(N__30209),
            .in2(_gnd_net_),
            .in3(N__20576),
            .lcout(data_out_frame2_18_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49673),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i89_LC_5_22_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i89_LC_5_22_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i89_LC_5_22_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_out_frame2_0___i89_LC_5_22_2  (
            .in0(N__29862),
            .in1(N__26345),
            .in2(_gnd_net_),
            .in3(N__24743),
            .lcout(data_out_frame2_11_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49673),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i134_LC_5_22_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i134_LC_5_22_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i134_LC_5_22_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i134_LC_5_22_3  (
            .in0(N__26339),
            .in1(N__30039),
            .in2(_gnd_net_),
            .in3(N__20547),
            .lcout(data_out_frame2_16_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49673),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i81_LC_5_22_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i81_LC_5_22_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i81_LC_5_22_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_out_frame2_0___i81_LC_5_22_4  (
            .in0(N__30406),
            .in1(N__26344),
            .in2(_gnd_net_),
            .in3(N__21360),
            .lcout(data_out_frame2_10_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49673),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i125_LC_5_22_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i125_LC_5_22_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i125_LC_5_22_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i125_LC_5_22_5  (
            .in0(N__26338),
            .in1(N__30645),
            .in2(_gnd_net_),
            .in3(N__20513),
            .lcout(data_out_frame2_15_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49673),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i120_LC_5_22_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i120_LC_5_22_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i120_LC_5_22_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_out_frame2_0___i120_LC_5_22_6  (
            .in0(N__30960),
            .in1(N__26342),
            .in2(_gnd_net_),
            .in3(N__22094),
            .lcout(data_out_frame2_14_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49673),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i71_LC_5_22_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i71_LC_5_22_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i71_LC_5_22_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i71_LC_5_22_7  (
            .in0(N__26341),
            .in1(N__29966),
            .in2(_gnd_net_),
            .in3(N__21509),
            .lcout(data_out_frame2_8_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49673),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2358__i0_LC_5_23_0.C_ON=1'b1;
    defparam rand_data_2358__i0_LC_5_23_0.SEQ_MODE=4'b1000;
    defparam rand_data_2358__i0_LC_5_23_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2358__i0_LC_5_23_0 (
            .in0(_gnd_net_),
            .in1(N__29431),
            .in2(_gnd_net_),
            .in3(N__20652),
            .lcout(rand_data_0),
            .ltout(),
            .carryin(bfn_5_23_0_),
            .carryout(n15979),
            .clk(N__49685),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2358__i1_LC_5_23_1.C_ON=1'b1;
    defparam rand_data_2358__i1_LC_5_23_1.SEQ_MODE=4'b1000;
    defparam rand_data_2358__i1_LC_5_23_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2358__i1_LC_5_23_1 (
            .in0(_gnd_net_),
            .in1(N__30250),
            .in2(_gnd_net_),
            .in3(N__20649),
            .lcout(rand_data_1),
            .ltout(),
            .carryin(n15979),
            .carryout(n15980),
            .clk(N__49685),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2358__i2_LC_5_23_2.C_ON=1'b1;
    defparam rand_data_2358__i2_LC_5_23_2.SEQ_MODE=4'b1000;
    defparam rand_data_2358__i2_LC_5_23_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2358__i2_LC_5_23_2 (
            .in0(_gnd_net_),
            .in1(N__30205),
            .in2(_gnd_net_),
            .in3(N__20646),
            .lcout(rand_data_2),
            .ltout(),
            .carryin(n15980),
            .carryout(n15981),
            .clk(N__49685),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2358__i3_LC_5_23_3.C_ON=1'b1;
    defparam rand_data_2358__i3_LC_5_23_3.SEQ_MODE=4'b1000;
    defparam rand_data_2358__i3_LC_5_23_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2358__i3_LC_5_23_3 (
            .in0(_gnd_net_),
            .in1(N__30143),
            .in2(_gnd_net_),
            .in3(N__20643),
            .lcout(rand_data_3),
            .ltout(),
            .carryin(n15981),
            .carryout(n15982),
            .clk(N__49685),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2358__i4_LC_5_23_4.C_ON=1'b1;
    defparam rand_data_2358__i4_LC_5_23_4.SEQ_MODE=4'b1000;
    defparam rand_data_2358__i4_LC_5_23_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2358__i4_LC_5_23_4 (
            .in0(_gnd_net_),
            .in1(N__30088),
            .in2(_gnd_net_),
            .in3(N__20640),
            .lcout(rand_data_4),
            .ltout(),
            .carryin(n15982),
            .carryout(n15983),
            .clk(N__49685),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2358__i5_LC_5_23_5.C_ON=1'b1;
    defparam rand_data_2358__i5_LC_5_23_5.SEQ_MODE=4'b1000;
    defparam rand_data_2358__i5_LC_5_23_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2358__i5_LC_5_23_5 (
            .in0(_gnd_net_),
            .in1(N__30031),
            .in2(_gnd_net_),
            .in3(N__20637),
            .lcout(rand_data_5),
            .ltout(),
            .carryin(n15983),
            .carryout(n15984),
            .clk(N__49685),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2358__i6_LC_5_23_6.C_ON=1'b1;
    defparam rand_data_2358__i6_LC_5_23_6.SEQ_MODE=4'b1000;
    defparam rand_data_2358__i6_LC_5_23_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2358__i6_LC_5_23_6 (
            .in0(_gnd_net_),
            .in1(N__29965),
            .in2(_gnd_net_),
            .in3(N__20634),
            .lcout(rand_data_6),
            .ltout(),
            .carryin(n15984),
            .carryout(n15985),
            .clk(N__49685),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2358__i7_LC_5_23_7.C_ON=1'b1;
    defparam rand_data_2358__i7_LC_5_23_7.SEQ_MODE=4'b1000;
    defparam rand_data_2358__i7_LC_5_23_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2358__i7_LC_5_23_7 (
            .in0(_gnd_net_),
            .in1(N__29903),
            .in2(_gnd_net_),
            .in3(N__20631),
            .lcout(rand_data_7),
            .ltout(),
            .carryin(n15985),
            .carryout(n15986),
            .clk(N__49685),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2358__i8_LC_5_24_0.C_ON=1'b1;
    defparam rand_data_2358__i8_LC_5_24_0.SEQ_MODE=4'b1000;
    defparam rand_data_2358__i8_LC_5_24_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2358__i8_LC_5_24_0 (
            .in0(_gnd_net_),
            .in1(N__29846),
            .in2(_gnd_net_),
            .in3(N__20628),
            .lcout(rand_data_8),
            .ltout(),
            .carryin(bfn_5_24_0_),
            .carryout(n15987),
            .clk(N__49696),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2358__i9_LC_5_24_1.C_ON=1'b1;
    defparam rand_data_2358__i9_LC_5_24_1.SEQ_MODE=4'b1000;
    defparam rand_data_2358__i9_LC_5_24_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2358__i9_LC_5_24_1 (
            .in0(_gnd_net_),
            .in1(N__29783),
            .in2(_gnd_net_),
            .in3(N__20679),
            .lcout(rand_data_9),
            .ltout(),
            .carryin(n15987),
            .carryout(n15988),
            .clk(N__49696),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2358__i10_LC_5_24_2.C_ON=1'b1;
    defparam rand_data_2358__i10_LC_5_24_2.SEQ_MODE=4'b1000;
    defparam rand_data_2358__i10_LC_5_24_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2358__i10_LC_5_24_2 (
            .in0(_gnd_net_),
            .in1(N__30751),
            .in2(_gnd_net_),
            .in3(N__20676),
            .lcout(rand_data_10),
            .ltout(),
            .carryin(n15988),
            .carryout(n15989),
            .clk(N__49696),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2358__i11_LC_5_24_3.C_ON=1'b1;
    defparam rand_data_2358__i11_LC_5_24_3.SEQ_MODE=4'b1000;
    defparam rand_data_2358__i11_LC_5_24_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2358__i11_LC_5_24_3 (
            .in0(_gnd_net_),
            .in1(N__30681),
            .in2(_gnd_net_),
            .in3(N__20673),
            .lcout(rand_data_11),
            .ltout(),
            .carryin(n15989),
            .carryout(n15990),
            .clk(N__49696),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2358__i12_LC_5_24_4.C_ON=1'b1;
    defparam rand_data_2358__i12_LC_5_24_4.SEQ_MODE=4'b1000;
    defparam rand_data_2358__i12_LC_5_24_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2358__i12_LC_5_24_4 (
            .in0(_gnd_net_),
            .in1(N__30629),
            .in2(_gnd_net_),
            .in3(N__20670),
            .lcout(rand_data_12),
            .ltout(),
            .carryin(n15990),
            .carryout(n15991),
            .clk(N__49696),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2358__i13_LC_5_24_5.C_ON=1'b1;
    defparam rand_data_2358__i13_LC_5_24_5.SEQ_MODE=4'b1000;
    defparam rand_data_2358__i13_LC_5_24_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2358__i13_LC_5_24_5 (
            .in0(_gnd_net_),
            .in1(N__30574),
            .in2(_gnd_net_),
            .in3(N__20667),
            .lcout(rand_data_13),
            .ltout(),
            .carryin(n15991),
            .carryout(n15992),
            .clk(N__49696),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2358__i14_LC_5_24_6.C_ON=1'b1;
    defparam rand_data_2358__i14_LC_5_24_6.SEQ_MODE=4'b1000;
    defparam rand_data_2358__i14_LC_5_24_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2358__i14_LC_5_24_6 (
            .in0(_gnd_net_),
            .in1(N__30502),
            .in2(_gnd_net_),
            .in3(N__20664),
            .lcout(rand_data_14),
            .ltout(),
            .carryin(n15992),
            .carryout(n15993),
            .clk(N__49696),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2358__i15_LC_5_24_7.C_ON=1'b1;
    defparam rand_data_2358__i15_LC_5_24_7.SEQ_MODE=4'b1000;
    defparam rand_data_2358__i15_LC_5_24_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2358__i15_LC_5_24_7 (
            .in0(_gnd_net_),
            .in1(N__30446),
            .in2(_gnd_net_),
            .in3(N__20661),
            .lcout(rand_data_15),
            .ltout(),
            .carryin(n15993),
            .carryout(n15994),
            .clk(N__49696),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2358__i16_LC_5_25_0.C_ON=1'b1;
    defparam rand_data_2358__i16_LC_5_25_0.SEQ_MODE=4'b1000;
    defparam rand_data_2358__i16_LC_5_25_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2358__i16_LC_5_25_0 (
            .in0(_gnd_net_),
            .in1(N__30392),
            .in2(_gnd_net_),
            .in3(N__20658),
            .lcout(rand_data_16),
            .ltout(),
            .carryin(bfn_5_25_0_),
            .carryout(n15995),
            .clk(N__49707),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2358__i17_LC_5_25_1.C_ON=1'b1;
    defparam rand_data_2358__i17_LC_5_25_1.SEQ_MODE=4'b1000;
    defparam rand_data_2358__i17_LC_5_25_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2358__i17_LC_5_25_1 (
            .in0(_gnd_net_),
            .in1(N__30329),
            .in2(_gnd_net_),
            .in3(N__20655),
            .lcout(rand_data_17),
            .ltout(),
            .carryin(n15995),
            .carryout(n15996),
            .clk(N__49707),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2358__i18_LC_5_25_2.C_ON=1'b1;
    defparam rand_data_2358__i18_LC_5_25_2.SEQ_MODE=4'b1000;
    defparam rand_data_2358__i18_LC_5_25_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2358__i18_LC_5_25_2 (
            .in0(_gnd_net_),
            .in1(N__31238),
            .in2(_gnd_net_),
            .in3(N__20706),
            .lcout(rand_data_18),
            .ltout(),
            .carryin(n15996),
            .carryout(n15997),
            .clk(N__49707),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2358__i19_LC_5_25_3.C_ON=1'b1;
    defparam rand_data_2358__i19_LC_5_25_3.SEQ_MODE=4'b1000;
    defparam rand_data_2358__i19_LC_5_25_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2358__i19_LC_5_25_3 (
            .in0(_gnd_net_),
            .in1(N__31181),
            .in2(_gnd_net_),
            .in3(N__20703),
            .lcout(rand_data_19),
            .ltout(),
            .carryin(n15997),
            .carryout(n15998),
            .clk(N__49707),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2358__i20_LC_5_25_4.C_ON=1'b1;
    defparam rand_data_2358__i20_LC_5_25_4.SEQ_MODE=4'b1000;
    defparam rand_data_2358__i20_LC_5_25_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2358__i20_LC_5_25_4 (
            .in0(_gnd_net_),
            .in1(N__31127),
            .in2(_gnd_net_),
            .in3(N__20700),
            .lcout(rand_data_20),
            .ltout(),
            .carryin(n15998),
            .carryout(n15999),
            .clk(N__49707),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2358__i21_LC_5_25_5.C_ON=1'b1;
    defparam rand_data_2358__i21_LC_5_25_5.SEQ_MODE=4'b1000;
    defparam rand_data_2358__i21_LC_5_25_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2358__i21_LC_5_25_5 (
            .in0(_gnd_net_),
            .in1(N__31064),
            .in2(_gnd_net_),
            .in3(N__20697),
            .lcout(rand_data_21),
            .ltout(),
            .carryin(n15999),
            .carryout(n16000),
            .clk(N__49707),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2358__i22_LC_5_25_6.C_ON=1'b1;
    defparam rand_data_2358__i22_LC_5_25_6.SEQ_MODE=4'b1000;
    defparam rand_data_2358__i22_LC_5_25_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2358__i22_LC_5_25_6 (
            .in0(_gnd_net_),
            .in1(N__31002),
            .in2(_gnd_net_),
            .in3(N__20694),
            .lcout(rand_data_22),
            .ltout(),
            .carryin(n16000),
            .carryout(n16001),
            .clk(N__49707),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2358__i23_LC_5_25_7.C_ON=1'b1;
    defparam rand_data_2358__i23_LC_5_25_7.SEQ_MODE=4'b1000;
    defparam rand_data_2358__i23_LC_5_25_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2358__i23_LC_5_25_7 (
            .in0(_gnd_net_),
            .in1(N__30948),
            .in2(_gnd_net_),
            .in3(N__20691),
            .lcout(rand_data_23),
            .ltout(),
            .carryin(n16001),
            .carryout(n16002),
            .clk(N__49707),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2358__i24_LC_5_26_0.C_ON=1'b1;
    defparam rand_data_2358__i24_LC_5_26_0.SEQ_MODE=4'b1000;
    defparam rand_data_2358__i24_LC_5_26_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2358__i24_LC_5_26_0 (
            .in0(_gnd_net_),
            .in1(N__30899),
            .in2(_gnd_net_),
            .in3(N__20688),
            .lcout(rand_data_24),
            .ltout(),
            .carryin(bfn_5_26_0_),
            .carryout(n16003),
            .clk(N__49720),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2358__i25_LC_5_26_1.C_ON=1'b1;
    defparam rand_data_2358__i25_LC_5_26_1.SEQ_MODE=4'b1000;
    defparam rand_data_2358__i25_LC_5_26_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2358__i25_LC_5_26_1 (
            .in0(_gnd_net_),
            .in1(N__30810),
            .in2(_gnd_net_),
            .in3(N__20685),
            .lcout(rand_data_25),
            .ltout(),
            .carryin(n16003),
            .carryout(n16004),
            .clk(N__49720),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2358__i26_LC_5_26_2.C_ON=1'b1;
    defparam rand_data_2358__i26_LC_5_26_2.SEQ_MODE=4'b1000;
    defparam rand_data_2358__i26_LC_5_26_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2358__i26_LC_5_26_2 (
            .in0(_gnd_net_),
            .in1(N__31655),
            .in2(_gnd_net_),
            .in3(N__20682),
            .lcout(rand_data_26),
            .ltout(),
            .carryin(n16004),
            .carryout(n16005),
            .clk(N__49720),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2358__i27_LC_5_26_3.C_ON=1'b1;
    defparam rand_data_2358__i27_LC_5_26_3.SEQ_MODE=4'b1000;
    defparam rand_data_2358__i27_LC_5_26_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2358__i27_LC_5_26_3 (
            .in0(_gnd_net_),
            .in1(N__31596),
            .in2(_gnd_net_),
            .in3(N__20742),
            .lcout(rand_data_27),
            .ltout(),
            .carryin(n16005),
            .carryout(n16006),
            .clk(N__49720),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2358__i28_LC_5_26_4.C_ON=1'b1;
    defparam rand_data_2358__i28_LC_5_26_4.SEQ_MODE=4'b1000;
    defparam rand_data_2358__i28_LC_5_26_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2358__i28_LC_5_26_4 (
            .in0(_gnd_net_),
            .in1(N__31544),
            .in2(_gnd_net_),
            .in3(N__20739),
            .lcout(rand_data_28),
            .ltout(),
            .carryin(n16006),
            .carryout(n16007),
            .clk(N__49720),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2358__i29_LC_5_26_5.C_ON=1'b1;
    defparam rand_data_2358__i29_LC_5_26_5.SEQ_MODE=4'b1000;
    defparam rand_data_2358__i29_LC_5_26_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2358__i29_LC_5_26_5 (
            .in0(_gnd_net_),
            .in1(N__31482),
            .in2(_gnd_net_),
            .in3(N__20736),
            .lcout(rand_data_29),
            .ltout(),
            .carryin(n16007),
            .carryout(n16008),
            .clk(N__49720),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2358__i30_LC_5_26_6.C_ON=1'b1;
    defparam rand_data_2358__i30_LC_5_26_6.SEQ_MODE=4'b1000;
    defparam rand_data_2358__i30_LC_5_26_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2358__i30_LC_5_26_6 (
            .in0(_gnd_net_),
            .in1(N__31430),
            .in2(_gnd_net_),
            .in3(N__20733),
            .lcout(rand_data_30),
            .ltout(),
            .carryin(n16008),
            .carryout(n16009),
            .clk(N__49720),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_data_2358__i31_LC_5_26_7.C_ON=1'b0;
    defparam rand_data_2358__i31_LC_5_26_7.SEQ_MODE=4'b1000;
    defparam rand_data_2358__i31_LC_5_26_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_data_2358__i31_LC_5_26_7 (
            .in0(_gnd_net_),
            .in1(N__31376),
            .in2(_gnd_net_),
            .in3(N__20730),
            .lcout(rand_data_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49720),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i6_LC_5_27_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i6_LC_5_27_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i6_LC_5_27_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i6_LC_5_27_0  (
            .in0(_gnd_net_),
            .in1(N__20727),
            .in2(_gnd_net_),
            .in3(N__33218),
            .lcout(\c0.FRAME_MATCHER_i_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49731),
            .ce(),
            .sr(N__20718));
    defparam \c0.i1_2_lut_adj_659_LC_5_27_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_659_LC_5_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_659_LC_5_27_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i1_2_lut_adj_659_LC_5_27_1  (
            .in0(_gnd_net_),
            .in1(N__25288),
            .in2(_gnd_net_),
            .in3(N__20877),
            .lcout(),
            .ltout(\c0.n26_adj_2373_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i19_4_lut_adj_669_LC_5_27_2 .C_ON=1'b0;
    defparam \c0.i19_4_lut_adj_669_LC_5_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.i19_4_lut_adj_669_LC_5_27_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i19_4_lut_adj_669_LC_5_27_2  (
            .in0(N__24993),
            .in1(N__27147),
            .in2(N__20721),
            .in3(N__27258),
            .lcout(\c0.n44_adj_2378 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_652_LC_5_27_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_652_LC_5_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_652_LC_5_27_3 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_652_LC_5_27_3  (
            .in0(N__41883),
            .in1(_gnd_net_),
            .in2(N__27830),
            .in3(N__20879),
            .lcout(\c0.n3_adj_2280 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_579_LC_5_27_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_579_LC_5_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_579_LC_5_27_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i1_2_lut_adj_579_LC_5_27_4  (
            .in0(N__20878),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41882),
            .lcout(\c0.n41 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_219_Select_15_i3_2_lut_3_lut_LC_5_27_5 .C_ON=1'b0;
    defparam \c0.select_219_Select_15_i3_2_lut_3_lut_LC_5_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.select_219_Select_15_i3_2_lut_3_lut_LC_5_27_5 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \c0.select_219_Select_15_i3_2_lut_3_lut_LC_5_27_5  (
            .in0(N__41885),
            .in1(_gnd_net_),
            .in2(N__27831),
            .in3(N__27259),
            .lcout(\c0.n3_adj_2261 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_219_Select_11_i3_2_lut_3_lut_LC_5_27_6 .C_ON=1'b0;
    defparam \c0.select_219_Select_11_i3_2_lut_3_lut_LC_5_27_6 .SEQ_MODE=4'b0000;
    defparam \c0.select_219_Select_11_i3_2_lut_3_lut_LC_5_27_6 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \c0.select_219_Select_11_i3_2_lut_3_lut_LC_5_27_6  (
            .in0(N__27151),
            .in1(N__27786),
            .in2(_gnd_net_),
            .in3(N__41884),
            .lcout(\c0.n3_adj_2270 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_219_Select_19_i3_2_lut_3_lut_LC_5_27_7 .C_ON=1'b0;
    defparam \c0.select_219_Select_19_i3_2_lut_3_lut_LC_5_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.select_219_Select_19_i3_2_lut_3_lut_LC_5_27_7 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \c0.select_219_Select_19_i3_2_lut_3_lut_LC_5_27_7  (
            .in0(N__41886),
            .in1(_gnd_net_),
            .in2(N__27832),
            .in3(N__24994),
            .lcout(\c0.n3_adj_2252 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17_4_lut_adj_660_LC_5_28_0 .C_ON=1'b0;
    defparam \c0.i17_4_lut_adj_660_LC_5_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.i17_4_lut_adj_660_LC_5_28_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i17_4_lut_adj_660_LC_5_28_0  (
            .in0(N__25054),
            .in1(N__20946),
            .in2(N__25119),
            .in3(N__20796),
            .lcout(\c0.n42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i17_LC_5_28_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i17_LC_5_28_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i17_LC_5_28_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i17_LC_5_28_1  (
            .in0(_gnd_net_),
            .in1(N__20814),
            .in2(_gnd_net_),
            .in3(N__33235),
            .lcout(\c0.FRAME_MATCHER_i_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49741),
            .ce(),
            .sr(N__20808));
    defparam \c0.select_219_Select_17_i3_2_lut_3_lut_LC_5_28_2 .C_ON=1'b0;
    defparam \c0.select_219_Select_17_i3_2_lut_3_lut_LC_5_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.select_219_Select_17_i3_2_lut_3_lut_LC_5_28_2 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \c0.select_219_Select_17_i3_2_lut_3_lut_LC_5_28_2  (
            .in0(N__41878),
            .in1(N__27796),
            .in2(_gnd_net_),
            .in3(N__20798),
            .lcout(\c0.n3_adj_2257 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10671_2_lut_LC_5_28_3 .C_ON=1'b0;
    defparam \c0.i10671_2_lut_LC_5_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.i10671_2_lut_LC_5_28_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i10671_2_lut_LC_5_28_3  (
            .in0(N__20797),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41877),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_219_Select_21_i3_2_lut_3_lut_LC_5_28_4 .C_ON=1'b0;
    defparam \c0.select_219_Select_21_i3_2_lut_3_lut_LC_5_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.select_219_Select_21_i3_2_lut_3_lut_LC_5_28_4 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \c0.select_219_Select_21_i3_2_lut_3_lut_LC_5_28_4  (
            .in0(N__41880),
            .in1(N__27795),
            .in2(_gnd_net_),
            .in3(N__20948),
            .lcout(\c0.n3_adj_2248 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_219_Select_20_i3_2_lut_3_lut_LC_5_28_5 .C_ON=1'b0;
    defparam \c0.select_219_Select_20_i3_2_lut_3_lut_LC_5_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.select_219_Select_20_i3_2_lut_3_lut_LC_5_28_5 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \c0.select_219_Select_20_i3_2_lut_3_lut_LC_5_28_5  (
            .in0(N__27793),
            .in1(N__25055),
            .in2(_gnd_net_),
            .in3(N__41879),
            .lcout(\c0.n3_adj_2250 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_219_Select_23_i3_2_lut_3_lut_LC_5_28_6 .C_ON=1'b0;
    defparam \c0.select_219_Select_23_i3_2_lut_3_lut_LC_5_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.select_219_Select_23_i3_2_lut_3_lut_LC_5_28_6 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \c0.select_219_Select_23_i3_2_lut_3_lut_LC_5_28_6  (
            .in0(N__41881),
            .in1(_gnd_net_),
            .in2(N__25120),
            .in3(N__27794),
            .lcout(\c0.n3_adj_2244 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10667_2_lut_LC_5_28_7 .C_ON=1'b0;
    defparam \c0.i10667_2_lut_LC_5_28_7 .SEQ_MODE=4'b0000;
    defparam \c0.i10667_2_lut_LC_5_28_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i10667_2_lut_LC_5_28_7  (
            .in0(N__20947),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41876),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i6_LC_5_29_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i6_LC_5_29_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i6_LC_5_29_0 .LUT_INIT=16'b1110000011000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i6_LC_5_29_0  (
            .in0(N__45019),
            .in1(N__44811),
            .in2(N__27395),
            .in3(N__44542),
            .lcout(\c0.FRAME_MATCHER_state_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49752),
            .ce(),
            .sr(N__27363));
    defparam \c0.select_219_Select_27_i3_2_lut_3_lut_LC_5_29_1 .C_ON=1'b0;
    defparam \c0.select_219_Select_27_i3_2_lut_3_lut_LC_5_29_1 .SEQ_MODE=4'b0000;
    defparam \c0.select_219_Select_27_i3_2_lut_3_lut_LC_5_29_1 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \c0.select_219_Select_27_i3_2_lut_3_lut_LC_5_29_1  (
            .in0(N__41870),
            .in1(_gnd_net_),
            .in2(N__22693),
            .in3(N__27781),
            .lcout(\c0.n3_adj_2236 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_686_LC_5_29_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_686_LC_5_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_686_LC_5_29_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_686_LC_5_29_2  (
            .in0(_gnd_net_),
            .in1(N__22683),
            .in2(_gnd_net_),
            .in3(N__41866),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_219_Select_8_i3_2_lut_3_lut_LC_5_29_3 .C_ON=1'b0;
    defparam \c0.select_219_Select_8_i3_2_lut_3_lut_LC_5_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.select_219_Select_8_i3_2_lut_3_lut_LC_5_29_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \c0.select_219_Select_8_i3_2_lut_3_lut_LC_5_29_3  (
            .in0(N__41871),
            .in1(N__27780),
            .in2(_gnd_net_),
            .in3(N__22194),
            .lcout(\c0.n3_adj_2276 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10680_2_lut_LC_5_29_4 .C_ON=1'b0;
    defparam \c0.i10680_2_lut_LC_5_29_4 .SEQ_MODE=4'b0000;
    defparam \c0.i10680_2_lut_LC_5_29_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i10680_2_lut_LC_5_29_4  (
            .in0(_gnd_net_),
            .in1(N__22193),
            .in2(_gnd_net_),
            .in3(N__41869),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_219_Select_9_i3_2_lut_3_lut_LC_5_29_5 .C_ON=1'b0;
    defparam \c0.select_219_Select_9_i3_2_lut_3_lut_LC_5_29_5 .SEQ_MODE=4'b0000;
    defparam \c0.select_219_Select_9_i3_2_lut_3_lut_LC_5_29_5 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \c0.select_219_Select_9_i3_2_lut_3_lut_LC_5_29_5  (
            .in0(N__41872),
            .in1(N__22631),
            .in2(_gnd_net_),
            .in3(N__27782),
            .lcout(\c0.n3_adj_2274 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10679_2_lut_LC_5_29_6 .C_ON=1'b0;
    defparam \c0.i10679_2_lut_LC_5_29_6 .SEQ_MODE=4'b0000;
    defparam \c0.i10679_2_lut_LC_5_29_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i10679_2_lut_LC_5_29_6  (
            .in0(N__22630),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41868),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10657_2_lut_LC_5_29_7 .C_ON=1'b0;
    defparam \c0.i10657_2_lut_LC_5_29_7 .SEQ_MODE=4'b0000;
    defparam \c0.i10657_2_lut_LC_5_29_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i10657_2_lut_LC_5_29_7  (
            .in0(N__41867),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29564),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i25_LC_5_30_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i25_LC_5_30_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i25_LC_5_30_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i25_LC_5_30_0  (
            .in0(_gnd_net_),
            .in1(N__21030),
            .in2(_gnd_net_),
            .in3(N__33236),
            .lcout(\c0.FRAME_MATCHER_i_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49765),
            .ce(),
            .sr(N__22476));
    defparam \c0.FRAME_MATCHER_i_i26_LC_5_31_3 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i26_LC_5_31_3 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i26_LC_5_31_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i26_LC_5_31_3  (
            .in0(_gnd_net_),
            .in1(N__21024),
            .in2(_gnd_net_),
            .in3(N__33250),
            .lcout(\c0.FRAME_MATCHER_i_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49777),
            .ce(),
            .sr(N__25257));
    defparam \c0.rx.i1_4_lut_adj_396_LC_5_32_0 .C_ON=1'b0;
    defparam \c0.rx.i1_4_lut_adj_396_LC_5_32_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_4_lut_adj_396_LC_5_32_0 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \c0.rx.i1_4_lut_adj_396_LC_5_32_0  (
            .in0(N__31866),
            .in1(N__22587),
            .in2(N__25560),
            .in3(N__22512),
            .lcout(\c0.rx.n10845 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_DV_52_LC_5_32_1 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_DV_52_LC_5_32_1 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_DV_52_LC_5_32_1 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \c0.rx.r_Rx_DV_52_LC_5_32_1  (
            .in0(N__25551),
            .in1(N__31868),
            .in2(N__39059),
            .in3(N__25638),
            .lcout(rx_data_ready),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49787),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_2__I_0_56_Mux_0_i1_3_lut_LC_5_32_2 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_2__I_0_56_Mux_0_i1_3_lut_LC_5_32_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.r_SM_Main_2__I_0_56_Mux_0_i1_3_lut_LC_5_32_2 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \c0.rx.r_SM_Main_2__I_0_56_Mux_0_i1_3_lut_LC_5_32_2  (
            .in0(N__25487),
            .in1(N__45267),
            .in2(_gnd_net_),
            .in3(N__22854),
            .lcout(n1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_2_lut_LC_5_32_3 .C_ON=1'b0;
    defparam \c0.rx.i2_2_lut_LC_5_32_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_2_lut_LC_5_32_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.rx.i2_2_lut_LC_5_32_3  (
            .in0(_gnd_net_),
            .in1(N__21002),
            .in2(_gnd_net_),
            .in3(N__20990),
            .lcout(\c0.rx.n6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i15215_4_lut_LC_5_32_4 .C_ON=1'b0;
    defparam \c0.rx.i15215_4_lut_LC_5_32_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i15215_4_lut_LC_5_32_4 .LUT_INIT=16'b0000110100001111;
    LogicCell40 \c0.rx.i15215_4_lut_LC_5_32_4  (
            .in0(N__25486),
            .in1(N__25550),
            .in2(N__31869),
            .in3(N__22839),
            .lcout(\c0.rx.n10656 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i15089_2_lut_LC_5_32_5 .C_ON=1'b0;
    defparam \c0.rx.i15089_2_lut_LC_5_32_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i15089_2_lut_LC_5_32_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.rx.i15089_2_lut_LC_5_32_5  (
            .in0(_gnd_net_),
            .in1(N__25488),
            .in2(_gnd_net_),
            .in3(N__25598),
            .lcout(),
            .ltout(n17708_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_i1_LC_5_32_6 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_i1_LC_5_32_6 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_SM_Main_i1_LC_5_32_6 .LUT_INIT=16'b0000010000010101;
    LogicCell40 \c0.rx.r_SM_Main_i1_LC_5_32_6  (
            .in0(N__31867),
            .in1(N__25552),
            .in2(N__21135),
            .in3(N__22581),
            .lcout(r_SM_Main_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49787),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Bit_Index_i2_LC_5_32_7 .C_ON=1'b0;
    defparam \c0.rx.r_Bit_Index_i2_LC_5_32_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Bit_Index_i2_LC_5_32_7 .LUT_INIT=16'b1011010000000000;
    LogicCell40 \c0.rx.r_Bit_Index_i2_LC_5_32_7  (
            .in0(N__25626),
            .in1(N__21132),
            .in2(N__37907),
            .in3(N__21120),
            .lcout(r_Bit_Index_2_adj_2435),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49787),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6489_2_lut_LC_6_14_4 .C_ON=1'b0;
    defparam \c0.i6489_2_lut_LC_6_14_4 .SEQ_MODE=4'b0000;
    defparam \c0.i6489_2_lut_LC_6_14_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i6489_2_lut_LC_6_14_4  (
            .in0(_gnd_net_),
            .in1(N__28585),
            .in2(_gnd_net_),
            .in3(N__28932),
            .lcout(\c0.n9157 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_0_i22_4_lut_LC_6_16_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_0_i22_4_lut_LC_6_16_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_0_i22_4_lut_LC_6_16_0 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_0_i22_4_lut_LC_6_16_0  (
            .in0(N__32142),
            .in1(N__21108),
            .in2(N__21699),
            .in3(N__21211),
            .lcout(\c0.n22_adj_2387 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_2_i6_4_lut_LC_6_16_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_2_i6_4_lut_LC_6_16_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_2_i6_4_lut_LC_6_16_2 .LUT_INIT=16'b1011100010001000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_2_i6_4_lut_LC_6_16_2  (
            .in0(N__23787),
            .in1(N__28613),
            .in2(N__24177),
            .in3(N__29003),
            .lcout(\c0.n6_adj_2140 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15435_LC_6_16_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15435_LC_6_16_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15435_LC_6_16_3 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_15435_LC_6_16_3  (
            .in0(N__21102),
            .in1(N__32369),
            .in2(N__21087),
            .in3(N__32141),
            .lcout(),
            .ltout(\c0.n18244_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18244_bdd_4_lut_LC_6_16_4 .C_ON=1'b0;
    defparam \c0.n18244_bdd_4_lut_LC_6_16_4 .SEQ_MODE=4'b0000;
    defparam \c0.n18244_bdd_4_lut_LC_6_16_4 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n18244_bdd_4_lut_LC_6_16_4  (
            .in0(N__32370),
            .in1(N__21072),
            .in2(N__21060),
            .in3(N__21057),
            .lcout(\c0.n18247 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Bit_Index_0__bdd_4_lut_LC_6_16_6 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_0__bdd_4_lut_LC_6_16_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_Bit_Index_0__bdd_4_lut_LC_6_16_6 .LUT_INIT=16'b1010111111000000;
    LogicCell40 \c0.tx2.r_Bit_Index_0__bdd_4_lut_LC_6_16_6  (
            .in0(N__21582),
            .in1(N__22812),
            .in2(N__25794),
            .in3(N__25736),
            .lcout(),
            .ltout(\c0.tx2.n18232_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.n18232_bdd_4_lut_LC_6_16_7 .C_ON=1'b0;
    defparam \c0.tx2.n18232_bdd_4_lut_LC_6_16_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.n18232_bdd_4_lut_LC_6_16_7 .LUT_INIT=16'b1111000011001010;
    LogicCell40 \c0.tx2.n18232_bdd_4_lut_LC_6_16_7  (
            .in0(N__21399),
            .in1(N__21051),
            .in2(N__21042),
            .in3(N__25791),
            .lcout(\c0.tx2.n18235 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i0_LC_6_17_0 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i0_LC_6_17_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i0_LC_6_17_0 .LUT_INIT=16'b0011101000001010;
    LogicCell40 \c0.tx2.r_Tx_Data_i0_LC_6_17_0  (
            .in0(N__21375),
            .in1(N__32414),
            .in2(N__32276),
            .in3(N__21405),
            .lcout(\c0.tx2.r_Tx_Data_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49640),
            .ce(N__24265),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15420_LC_6_17_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15420_LC_6_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15420_LC_6_17_2 .LUT_INIT=16'b1011101111000000;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_15420_LC_6_17_2  (
            .in0(N__21393),
            .in1(N__32412),
            .in2(N__21321),
            .in3(N__32149),
            .lcout(),
            .ltout(\c0.n18226_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18226_bdd_4_lut_LC_6_17_3 .C_ON=1'b0;
    defparam \c0.n18226_bdd_4_lut_LC_6_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.n18226_bdd_4_lut_LC_6_17_3 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n18226_bdd_4_lut_LC_6_17_3  (
            .in0(N__32413),
            .in1(N__21384),
            .in2(N__21378),
            .in3(N__21246),
            .lcout(\c0.n18229 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15351_LC_6_17_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15351_LC_6_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15351_LC_6_17_4 .LUT_INIT=16'b1110110000101100;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15351_LC_6_17_4  (
            .in0(N__21368),
            .in1(N__28891),
            .in2(N__28661),
            .in3(N__24750),
            .lcout(),
            .ltout(\c0.n18148_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18148_bdd_4_lut_LC_6_17_5 .C_ON=1'b0;
    defparam \c0.n18148_bdd_4_lut_LC_6_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.n18148_bdd_4_lut_LC_6_17_5 .LUT_INIT=16'b1111000010101100;
    LogicCell40 \c0.n18148_bdd_4_lut_LC_6_17_5  (
            .in0(N__41108),
            .in1(N__24323),
            .in2(N__21324),
            .in3(N__28610),
            .lcout(\c0.n18151 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_0_i6_4_lut_LC_6_17_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_0_i6_4_lut_LC_6_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_0_i6_4_lut_LC_6_17_6 .LUT_INIT=16'b1110010010100000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_0_i6_4_lut_LC_6_17_6  (
            .in0(N__28611),
            .in1(N__21312),
            .in2(N__21267),
            .in3(N__28892),
            .lcout(\c0.n6_adj_2143 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15274_LC_6_18_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15274_LC_6_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15274_LC_6_18_0 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15274_LC_6_18_0  (
            .in0(N__21416),
            .in1(N__28614),
            .in2(N__21240),
            .in3(N__28938),
            .lcout(),
            .ltout(\c0.n18052_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18052_bdd_4_lut_LC_6_18_1 .C_ON=1'b0;
    defparam \c0.n18052_bdd_4_lut_LC_6_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.n18052_bdd_4_lut_LC_6_18_1 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n18052_bdd_4_lut_LC_6_18_1  (
            .in0(N__28615),
            .in1(N__21681),
            .in2(N__21228),
            .in3(N__24481),
            .lcout(),
            .ltout(\c0.n18055_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_3_i22_4_lut_LC_6_18_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_3_i22_4_lut_LC_6_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_3_i22_4_lut_LC_6_18_2 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_3_i22_4_lut_LC_6_18_2  (
            .in0(N__32167),
            .in1(N__21225),
            .in2(N__21216),
            .in3(N__21194),
            .lcout(\c0.n22_adj_2371 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15440_LC_6_18_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15440_LC_6_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_2__bdd_4_lut_15440_LC_6_18_3 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter2_2__bdd_4_lut_15440_LC_6_18_3  (
            .in0(N__23322),
            .in1(N__32415),
            .in2(N__21615),
            .in3(N__32168),
            .lcout(),
            .ltout(\c0.n18256_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18256_bdd_4_lut_LC_6_18_4 .C_ON=1'b0;
    defparam \c0.n18256_bdd_4_lut_LC_6_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.n18256_bdd_4_lut_LC_6_18_4 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n18256_bdd_4_lut_LC_6_18_4  (
            .in0(N__32416),
            .in1(N__28716),
            .in2(N__21600),
            .in3(N__21597),
            .lcout(),
            .ltout(\c0.n18259_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i3_LC_6_18_5 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i3_LC_6_18_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i3_LC_6_18_5 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \c0.tx2.r_Tx_Data_i3_LC_6_18_5  (
            .in0(N__21591),
            .in1(N__32417),
            .in2(N__21585),
            .in3(N__32277),
            .lcout(\c0.tx2.r_Tx_Data_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49652),
            .ce(N__24254),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i82_LC_6_19_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i82_LC_6_19_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i82_LC_6_19_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i82_LC_6_19_0  (
            .in0(N__26514),
            .in1(N__30363),
            .in2(_gnd_net_),
            .in3(N__21564),
            .lcout(data_out_frame2_10_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49658),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i42_LC_6_19_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i42_LC_6_19_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i42_LC_6_19_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_out_frame2_0___i42_LC_6_19_1  (
            .in0(N__23397),
            .in1(N__30842),
            .in2(_gnd_net_),
            .in3(N__26516),
            .lcout(data_out_frame2_5_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49658),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_680_LC_6_19_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_680_LC_6_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_680_LC_6_19_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_680_LC_6_19_2  (
            .in0(N__23137),
            .in1(N__21860),
            .in2(_gnd_net_),
            .in3(N__21895),
            .lcout(\c0.n17203 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18124_bdd_4_lut_LC_6_19_3 .C_ON=1'b0;
    defparam \c0.n18124_bdd_4_lut_LC_6_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.n18124_bdd_4_lut_LC_6_19_3 .LUT_INIT=16'b1100110011100010;
    LogicCell40 \c0.n18124_bdd_4_lut_LC_6_19_3  (
            .in0(N__21523),
            .in1(N__23103),
            .in2(N__21474),
            .in3(N__28505),
            .lcout(\c0.n18127 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i148_LC_6_19_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i148_LC_6_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i148_LC_6_19_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i148_LC_6_19_4  (
            .in0(N__26513),
            .in1(N__30169),
            .in2(_gnd_net_),
            .in3(N__21417),
            .lcout(data_out_frame2_18_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49658),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i136_LC_6_19_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i136_LC_6_19_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i136_LC_6_19_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i136_LC_6_19_5  (
            .in0(N__29931),
            .in1(N__27635),
            .in2(_gnd_net_),
            .in3(N__26515),
            .lcout(data_out_frame2_16_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49658),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18160_bdd_4_lut_LC_6_19_6 .C_ON=1'b0;
    defparam \c0.n18160_bdd_4_lut_LC_6_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.n18160_bdd_4_lut_LC_6_19_6 .LUT_INIT=16'b1101100111001000;
    LogicCell40 \c0.n18160_bdd_4_lut_LC_6_19_6  (
            .in0(N__28506),
            .in1(N__23073),
            .in2(N__21717),
            .in3(N__24941),
            .lcout(\c0.n18163 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15450_LC_6_19_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15450_LC_6_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15450_LC_6_19_7 .LUT_INIT=16'b1011101111000000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15450_LC_6_19_7  (
            .in0(N__21894),
            .in1(N__28504),
            .in2(N__24138),
            .in3(N__28999),
            .lcout(\c0.n18208 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i140_LC_6_20_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i140_LC_6_20_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i140_LC_6_20_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i140_LC_6_20_0  (
            .in0(N__30717),
            .in1(N__21680),
            .in2(_gnd_net_),
            .in3(N__26370),
            .lcout(data_out_frame2_17_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49666),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i127_LC_6_20_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i127_LC_6_20_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i127_LC_6_20_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i127_LC_6_20_1  (
            .in0(N__26366),
            .in1(N__30536),
            .in2(_gnd_net_),
            .in3(N__23012),
            .lcout(data_out_frame2_15_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49666),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i145_LC_6_20_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i145_LC_6_20_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i145_LC_6_20_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_out_frame2_0___i145_LC_6_20_2  (
            .in0(N__23085),
            .in1(N__29454),
            .in2(_gnd_net_),
            .in3(N__26371),
            .lcout(data_out_frame2_18_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49666),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i87_LC_6_20_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i87_LC_6_20_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i87_LC_6_20_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i87_LC_6_20_3  (
            .in0(N__26368),
            .in1(N__31026),
            .in2(_gnd_net_),
            .in3(N__23184),
            .lcout(data_out_frame2_10_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49666),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i106_LC_6_20_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i106_LC_6_20_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i106_LC_6_20_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i106_LC_6_20_4  (
            .in0(N__30834),
            .in1(N__23652),
            .in2(_gnd_net_),
            .in3(N__26369),
            .lcout(data_out_frame2_13_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49666),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i115_LC_6_20_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i115_LC_6_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i115_LC_6_20_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i115_LC_6_20_5  (
            .in0(N__26365),
            .in1(N__31264),
            .in2(_gnd_net_),
            .in3(N__21660),
            .lcout(data_out_frame2_14_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49666),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_4_lut_adj_724_LC_6_20_6 .C_ON=1'b0;
    defparam \c0.i5_3_lut_4_lut_adj_724_LC_6_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_4_lut_adj_724_LC_6_20_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_3_lut_4_lut_adj_724_LC_6_20_6  (
            .in0(N__41098),
            .in1(N__41149),
            .in2(N__21787),
            .in3(N__21630),
            .lcout(\c0.n17095 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i59_LC_6_20_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i59_LC_6_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i59_LC_6_20_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i59_LC_6_20_7  (
            .in0(N__26367),
            .in1(N__30782),
            .in2(_gnd_net_),
            .in3(N__23844),
            .lcout(data_out_frame2_7_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49666),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i43_LC_6_21_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i43_LC_6_21_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i43_LC_6_21_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i43_LC_6_21_0  (
            .in0(N__26353),
            .in1(N__31674),
            .in2(_gnd_net_),
            .in3(N__24163),
            .lcout(data_out_frame2_5_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49674),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i119_LC_6_21_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i119_LC_6_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i119_LC_6_21_1 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \c0.data_out_frame2_0___i119_LC_6_21_1  (
            .in0(N__24526),
            .in1(_gnd_net_),
            .in2(N__31032),
            .in3(N__26356),
            .lcout(data_out_frame2_14_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49674),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i85_LC_6_21_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i85_LC_6_21_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i85_LC_6_21_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i85_LC_6_21_2  (
            .in0(N__26355),
            .in1(N__31149),
            .in2(_gnd_net_),
            .in3(N__24133),
            .lcout(data_out_frame2_10_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49674),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_672_LC_6_21_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_672_LC_6_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_672_LC_6_21_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_672_LC_6_21_3  (
            .in0(N__23123),
            .in1(N__21893),
            .in2(N__21867),
            .in3(N__24024),
            .lcout(\c0.n10359 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i45_LC_6_21_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i45_LC_6_21_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i45_LC_6_21_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i45_LC_6_21_4  (
            .in0(N__26354),
            .in1(N__31564),
            .in2(_gnd_net_),
            .in3(N__21783),
            .lcout(data_out_frame2_5_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49674),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i95_LC_6_21_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i95_LC_6_21_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i95_LC_6_21_5 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \c0.data_out_frame2_0___i95_LC_6_21_5  (
            .in0(N__23124),
            .in1(_gnd_net_),
            .in2(N__30537),
            .in3(N__26358),
            .lcout(data_out_frame2_11_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49674),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15346_LC_6_21_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15346_LC_6_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15346_LC_6_21_6 .LUT_INIT=16'b1010111111000000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15346_LC_6_21_6  (
            .in0(N__23255),
            .in1(N__21740),
            .in2(N__28599),
            .in3(N__28960),
            .lcout(\c0.n18142 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i88_LC_6_21_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i88_LC_6_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i88_LC_6_21_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_out_frame2_0___i88_LC_6_21_7  (
            .in0(N__21741),
            .in1(N__30975),
            .in2(_gnd_net_),
            .in3(N__26357),
            .lcout(data_out_frame2_10_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49674),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i11067_2_lut_4_lut_LC_6_22_0 .C_ON=1'b0;
    defparam \c0.tx2.i11067_2_lut_4_lut_LC_6_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i11067_2_lut_4_lut_LC_6_22_0 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \c0.tx2.i11067_2_lut_4_lut_LC_6_22_0  (
            .in0(N__22145),
            .in1(N__26839),
            .in2(N__22287),
            .in3(N__22044),
            .lcout(),
            .ltout(\c0.tx2.n13748_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i1_4_lut_LC_6_22_1 .C_ON=1'b0;
    defparam \c0.tx2.i1_4_lut_LC_6_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i1_4_lut_LC_6_22_1 .LUT_INIT=16'b0000000000001110;
    LogicCell40 \c0.tx2.i1_4_lut_LC_6_22_1  (
            .in0(N__26742),
            .in1(N__25941),
            .in2(N__22008),
            .in3(N__22068),
            .lcout(\c0.tx2.n17322 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i73_LC_6_22_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i73_LC_6_22_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i73_LC_6_22_2 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \c0.data_out_frame2_0___i73_LC_6_22_2  (
            .in0(N__26374),
            .in1(N__30919),
            .in2(N__41105),
            .in3(_gnd_net_),
            .lcout(data_out_frame2_9_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49686),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i152_LC_6_22_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i152_LC_6_22_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i152_LC_6_22_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i152_LC_6_22_3  (
            .in0(N__29912),
            .in1(N__22001),
            .in2(_gnd_net_),
            .in3(N__26376),
            .lcout(data_out_frame2_18_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49686),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i139_LC_6_22_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i139_LC_6_22_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i139_LC_6_22_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i139_LC_6_22_4  (
            .in0(N__26372),
            .in1(N__30781),
            .in2(_gnd_net_),
            .in3(N__21977),
            .lcout(data_out_frame2_17_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49686),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i1_2_lut_4_lut_LC_6_22_5 .C_ON=1'b0;
    defparam \c0.tx2.i1_2_lut_4_lut_LC_6_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i1_2_lut_4_lut_LC_6_22_5 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \c0.tx2.i1_2_lut_4_lut_LC_6_22_5  (
            .in0(N__22043),
            .in1(N__22067),
            .in2(N__22146),
            .in3(N__22283),
            .lcout(r_SM_Main_2_N_2031_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i70_LC_6_22_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i70_LC_6_22_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i70_LC_6_22_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i70_LC_6_22_6  (
            .in0(N__26373),
            .in1(N__30032),
            .in2(_gnd_net_),
            .in3(N__40925),
            .lcout(data_out_frame2_8_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49686),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i109_LC_6_22_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i109_LC_6_22_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i109_LC_6_22_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i109_LC_6_22_7  (
            .in0(N__31563),
            .in1(N__41144),
            .in2(_gnd_net_),
            .in3(N__26375),
            .lcout(data_out_frame2_13_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49686),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i62_LC_6_23_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i62_LC_6_23_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i62_LC_6_23_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_out_frame2_0___i62_LC_6_23_0  (
            .in0(N__21955),
            .in1(N__30584),
            .in2(_gnd_net_),
            .in3(N__26566),
            .lcout(data_out_frame2_7_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49697),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i69_LC_6_23_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i69_LC_6_23_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i69_LC_6_23_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i69_LC_6_23_1  (
            .in0(N__26565),
            .in1(N__30104),
            .in2(_gnd_net_),
            .in3(N__24358),
            .lcout(data_out_frame2_8_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49697),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i4_4_lut_LC_6_23_2 .C_ON=1'b0;
    defparam \c0.tx2.i4_4_lut_LC_6_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i4_4_lut_LC_6_23_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.tx2.i4_4_lut_LC_6_23_2  (
            .in0(N__22058),
            .in1(N__22323),
            .in2(N__22305),
            .in3(N__22022),
            .lcout(\c0.tx2.n10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.o_Tx_Serial_45_LC_6_23_3 .C_ON=1'b0;
    defparam \c0.tx2.o_Tx_Serial_45_LC_6_23_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.o_Tx_Serial_45_LC_6_23_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.tx2.o_Tx_Serial_45_LC_6_23_3  (
            .in0(N__22114),
            .in1(N__25672),
            .in2(_gnd_net_),
            .in3(N__22719),
            .lcout(tx2_o),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49697),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i65_LC_6_23_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i65_LC_6_23_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i65_LC_6_23_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i65_LC_6_23_4  (
            .in0(N__29453),
            .in1(N__24316),
            .in2(_gnd_net_),
            .in3(N__26567),
            .lcout(data_out_frame2_8_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49697),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_613_LC_6_23_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_613_LC_6_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_613_LC_6_23_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_613_LC_6_23_5  (
            .in0(_gnd_net_),
            .in1(N__24596),
            .in2(_gnd_net_),
            .in3(N__22093),
            .lcout(\c0.n10563 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i15218_2_lut_LC_6_23_6 .C_ON=1'b0;
    defparam \c0.tx2.i15218_2_lut_LC_6_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i15218_2_lut_LC_6_23_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \c0.tx2.i15218_2_lut_LC_6_23_6  (
            .in0(_gnd_net_),
            .in1(N__22074),
            .in2(_gnd_net_),
            .in3(N__26852),
            .lcout(\c0.tx2.n10852 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i2_3_lut_LC_6_23_7 .C_ON=1'b0;
    defparam \c0.tx2.i2_3_lut_LC_6_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i2_3_lut_LC_6_23_7 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.tx2.i2_3_lut_LC_6_23_7  (
            .in0(N__22230),
            .in1(N__22262),
            .in2(_gnd_net_),
            .in3(N__22247),
            .lcout(\c0.tx2.n17018 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Clock_Count__i0_LC_6_24_0 .C_ON=1'b1;
    defparam \c0.tx2.r_Clock_Count__i0_LC_6_24_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i0_LC_6_24_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx2.r_Clock_Count__i0_LC_6_24_0  (
            .in0(_gnd_net_),
            .in1(N__22059),
            .in2(_gnd_net_),
            .in3(N__22047),
            .lcout(\c0.tx2.r_Clock_Count_0 ),
            .ltout(),
            .carryin(bfn_6_24_0_),
            .carryout(\c0.tx2.n16132 ),
            .clk(N__49708),
            .ce(N__25676),
            .sr(N__22215));
    defparam \c0.tx2.r_Clock_Count__i1_LC_6_24_1 .C_ON=1'b1;
    defparam \c0.tx2.r_Clock_Count__i1_LC_6_24_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i1_LC_6_24_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx2.r_Clock_Count__i1_LC_6_24_1  (
            .in0(_gnd_net_),
            .in1(N__22042),
            .in2(_gnd_net_),
            .in3(N__22026),
            .lcout(\c0.tx2.r_Clock_Count_1 ),
            .ltout(),
            .carryin(\c0.tx2.n16132 ),
            .carryout(\c0.tx2.n16133 ),
            .clk(N__49708),
            .ce(N__25676),
            .sr(N__22215));
    defparam \c0.tx2.r_Clock_Count__i2_LC_6_24_2 .C_ON=1'b1;
    defparam \c0.tx2.r_Clock_Count__i2_LC_6_24_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i2_LC_6_24_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx2.r_Clock_Count__i2_LC_6_24_2  (
            .in0(_gnd_net_),
            .in1(N__22023),
            .in2(_gnd_net_),
            .in3(N__22011),
            .lcout(\c0.tx2.r_Clock_Count_2 ),
            .ltout(),
            .carryin(\c0.tx2.n16133 ),
            .carryout(\c0.tx2.n16134 ),
            .clk(N__49708),
            .ce(N__25676),
            .sr(N__22215));
    defparam \c0.tx2.r_Clock_Count__i3_LC_6_24_3 .C_ON=1'b1;
    defparam \c0.tx2.r_Clock_Count__i3_LC_6_24_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i3_LC_6_24_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx2.r_Clock_Count__i3_LC_6_24_3  (
            .in0(_gnd_net_),
            .in1(N__22322),
            .in2(_gnd_net_),
            .in3(N__22308),
            .lcout(\c0.tx2.r_Clock_Count_3 ),
            .ltout(),
            .carryin(\c0.tx2.n16134 ),
            .carryout(\c0.tx2.n16135 ),
            .clk(N__49708),
            .ce(N__25676),
            .sr(N__22215));
    defparam \c0.tx2.r_Clock_Count__i4_LC_6_24_4 .C_ON=1'b1;
    defparam \c0.tx2.r_Clock_Count__i4_LC_6_24_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i4_LC_6_24_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx2.r_Clock_Count__i4_LC_6_24_4  (
            .in0(_gnd_net_),
            .in1(N__22304),
            .in2(_gnd_net_),
            .in3(N__22290),
            .lcout(\c0.tx2.r_Clock_Count_4 ),
            .ltout(),
            .carryin(\c0.tx2.n16135 ),
            .carryout(\c0.tx2.n16136 ),
            .clk(N__49708),
            .ce(N__25676),
            .sr(N__22215));
    defparam \c0.tx2.r_Clock_Count__i5_LC_6_24_5 .C_ON=1'b1;
    defparam \c0.tx2.r_Clock_Count__i5_LC_6_24_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i5_LC_6_24_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx2.r_Clock_Count__i5_LC_6_24_5  (
            .in0(_gnd_net_),
            .in1(N__22282),
            .in2(_gnd_net_),
            .in3(N__22266),
            .lcout(\c0.tx2.r_Clock_Count_5 ),
            .ltout(),
            .carryin(\c0.tx2.n16136 ),
            .carryout(\c0.tx2.n16137 ),
            .clk(N__49708),
            .ce(N__25676),
            .sr(N__22215));
    defparam \c0.tx2.r_Clock_Count__i6_LC_6_24_6 .C_ON=1'b1;
    defparam \c0.tx2.r_Clock_Count__i6_LC_6_24_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i6_LC_6_24_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx2.r_Clock_Count__i6_LC_6_24_6  (
            .in0(_gnd_net_),
            .in1(N__22263),
            .in2(_gnd_net_),
            .in3(N__22251),
            .lcout(\c0.tx2.r_Clock_Count_6 ),
            .ltout(),
            .carryin(\c0.tx2.n16137 ),
            .carryout(\c0.tx2.n16138 ),
            .clk(N__49708),
            .ce(N__25676),
            .sr(N__22215));
    defparam \c0.tx2.r_Clock_Count__i7_LC_6_24_7 .C_ON=1'b1;
    defparam \c0.tx2.r_Clock_Count__i7_LC_6_24_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i7_LC_6_24_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx2.r_Clock_Count__i7_LC_6_24_7  (
            .in0(_gnd_net_),
            .in1(N__22248),
            .in2(_gnd_net_),
            .in3(N__22236),
            .lcout(\c0.tx2.r_Clock_Count_7 ),
            .ltout(),
            .carryin(\c0.tx2.n16138 ),
            .carryout(\c0.tx2.n16139 ),
            .clk(N__49708),
            .ce(N__25676),
            .sr(N__22215));
    defparam \c0.tx2.r_Clock_Count__i8_LC_6_25_0 .C_ON=1'b0;
    defparam \c0.tx2.r_Clock_Count__i8_LC_6_25_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Clock_Count__i8_LC_6_25_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.tx2.r_Clock_Count__i8_LC_6_25_0  (
            .in0(_gnd_net_),
            .in1(N__22229),
            .in2(_gnd_net_),
            .in3(N__22233),
            .lcout(\c0.tx2.r_Clock_Count_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49721),
            .ce(N__25677),
            .sr(N__22214));
    defparam \c0.i14_4_lut_adj_668_LC_6_26_0 .C_ON=1'b0;
    defparam \c0.i14_4_lut_adj_668_LC_6_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_adj_668_LC_6_26_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i14_4_lut_adj_668_LC_6_26_0  (
            .in0(N__22694),
            .in1(N__25431),
            .in2(N__25342),
            .in3(N__27996),
            .lcout(\c0.n39_adj_2377 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_639_LC_6_26_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_639_LC_6_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_639_LC_6_26_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i1_2_lut_adj_639_LC_6_26_1  (
            .in0(_gnd_net_),
            .in1(N__37077),
            .in2(_gnd_net_),
            .in3(N__22373),
            .lcout(\c0.n10161 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_4_lut_adj_666_LC_6_26_2 .C_ON=1'b0;
    defparam \c0.i16_4_lut_adj_666_LC_6_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.i16_4_lut_adj_666_LC_6_26_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i16_4_lut_adj_666_LC_6_26_2  (
            .in0(N__22626),
            .in1(N__27928),
            .in2(N__27890),
            .in3(N__22182),
            .lcout(),
            .ltout(\c0.n41_adj_2376_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i23_4_lut_LC_6_26_3 .C_ON=1'b0;
    defparam \c0.i23_4_lut_LC_6_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.i23_4_lut_LC_6_26_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i23_4_lut_LC_6_26_3  (
            .in0(N__22416),
            .in1(N__22506),
            .in2(N__22407),
            .in3(N__22404),
            .lcout(),
            .ltout(\c0.n48_adj_2379_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_675_LC_6_26_4 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_675_LC_6_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_675_LC_6_26_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i1_4_lut_adj_675_LC_6_26_4  (
            .in0(N__22398),
            .in1(N__32791),
            .in2(N__22386),
            .in3(N__22383),
            .lcout(\c0.n9995 ),
            .ltout(\c0.n9995_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10584_4_lut_LC_6_26_5 .C_ON=1'b0;
    defparam \c0.i10584_4_lut_LC_6_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.i10584_4_lut_LC_6_26_5 .LUT_INIT=16'b0101010001010000;
    LogicCell40 \c0.i10584_4_lut_LC_6_26_5  (
            .in0(N__29560),
            .in1(N__32865),
            .in2(N__22377),
            .in3(N__32640),
            .lcout(n3779),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10579_2_lut_3_lut_LC_6_27_0 .C_ON=1'b0;
    defparam \c0.i10579_2_lut_3_lut_LC_6_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10579_2_lut_3_lut_LC_6_27_0 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \c0.i10579_2_lut_3_lut_LC_6_27_0  (
            .in0(N__37079),
            .in1(N__29558),
            .in2(_gnd_net_),
            .in3(N__22374),
            .lcout(n4408),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i2_LC_6_27_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i2_LC_6_27_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i2_LC_6_27_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i2_LC_6_27_1  (
            .in0(_gnd_net_),
            .in1(N__22362),
            .in2(_gnd_net_),
            .in3(N__33185),
            .lcout(\c0.FRAME_MATCHER_i_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49742),
            .ce(),
            .sr(N__22353));
    defparam \c0.select_219_Select_2_i3_2_lut_3_lut_LC_6_27_2 .C_ON=1'b0;
    defparam \c0.select_219_Select_2_i3_2_lut_3_lut_LC_6_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.select_219_Select_2_i3_2_lut_3_lut_LC_6_27_2 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \c0.select_219_Select_2_i3_2_lut_3_lut_LC_6_27_2  (
            .in0(N__37081),
            .in1(_gnd_net_),
            .in2(N__27833),
            .in3(N__41874),
            .lcout(\c0.n3_adj_2286 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_219_Select_31_i3_2_lut_3_lut_LC_6_27_3 .C_ON=1'b0;
    defparam \c0.select_219_Select_31_i3_2_lut_3_lut_LC_6_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.select_219_Select_31_i3_2_lut_3_lut_LC_6_27_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \c0.select_219_Select_31_i3_2_lut_3_lut_LC_6_27_3  (
            .in0(N__41875),
            .in1(N__27801),
            .in2(_gnd_net_),
            .in3(N__29559),
            .lcout(\c0.n3_adj_2226 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10686_2_lut_LC_6_27_4 .C_ON=1'b0;
    defparam \c0.i10686_2_lut_LC_6_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.i10686_2_lut_LC_6_27_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i10686_2_lut_LC_6_27_4  (
            .in0(N__37080),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41873),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_658_LC_6_27_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_658_LC_6_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_658_LC_6_27_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_658_LC_6_27_5  (
            .in0(_gnd_net_),
            .in1(N__37156),
            .in2(_gnd_net_),
            .in3(N__37078),
            .lcout(\c0.n39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_adj_661_LC_6_28_0 .C_ON=1'b0;
    defparam \c0.i15_4_lut_adj_661_LC_6_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_adj_661_LC_6_28_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i15_4_lut_adj_661_LC_6_28_0  (
            .in0(N__25218),
            .in1(N__27025),
            .in2(N__33657),
            .in3(N__25158),
            .lcout(\c0.n40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i24_LC_6_28_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i24_LC_6_28_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i24_LC_6_28_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i24_LC_6_28_1  (
            .in0(N__33186),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22497),
            .lcout(\c0.FRAME_MATCHER_i_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49753),
            .ce(),
            .sr(N__22485));
    defparam \c0.select_219_Select_24_i3_2_lut_3_lut_LC_6_28_2 .C_ON=1'b0;
    defparam \c0.select_219_Select_24_i3_2_lut_3_lut_LC_6_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.select_219_Select_24_i3_2_lut_3_lut_LC_6_28_2 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \c0.select_219_Select_24_i3_2_lut_3_lut_LC_6_28_2  (
            .in0(N__41889),
            .in1(N__27800),
            .in2(_gnd_net_),
            .in3(N__25159),
            .lcout(\c0.n3_adj_2242 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_219_Select_25_i3_2_lut_3_lut_LC_6_28_3 .C_ON=1'b0;
    defparam \c0.select_219_Select_25_i3_2_lut_3_lut_LC_6_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.select_219_Select_25_i3_2_lut_3_lut_LC_6_28_3 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \c0.select_219_Select_25_i3_2_lut_3_lut_LC_6_28_3  (
            .in0(N__27797),
            .in1(N__25219),
            .in2(_gnd_net_),
            .in3(N__41890),
            .lcout(\c0.n3_adj_2240 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_219_Select_28_i3_2_lut_3_lut_LC_6_28_4 .C_ON=1'b0;
    defparam \c0.select_219_Select_28_i3_2_lut_3_lut_LC_6_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.select_219_Select_28_i3_2_lut_3_lut_LC_6_28_4 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \c0.select_219_Select_28_i3_2_lut_3_lut_LC_6_28_4  (
            .in0(N__41888),
            .in1(N__27799),
            .in2(_gnd_net_),
            .in3(N__27026),
            .lcout(\c0.n3_adj_2234 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_219_Select_30_i3_2_lut_3_lut_LC_6_28_5 .C_ON=1'b0;
    defparam \c0.select_219_Select_30_i3_2_lut_3_lut_LC_6_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.select_219_Select_30_i3_2_lut_3_lut_LC_6_28_5 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \c0.select_219_Select_30_i3_2_lut_3_lut_LC_6_28_5  (
            .in0(N__27798),
            .in1(N__33655),
            .in2(_gnd_net_),
            .in3(N__41891),
            .lcout(\c0.n3_adj_2230 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_4_lut_LC_6_28_6 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_4_lut_LC_6_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_4_lut_LC_6_28_6 .LUT_INIT=16'b1010101111111011;
    LogicCell40 \c0.i1_3_lut_4_lut_4_lut_LC_6_28_6  (
            .in0(N__35492),
            .in1(N__33444),
            .in2(N__35766),
            .in3(N__35832),
            .lcout(\c0.n10009 ),
            .ltout(\c0.n10009_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_588_LC_6_28_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_588_LC_6_28_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_588_LC_6_28_7 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_588_LC_6_28_7  (
            .in0(N__37185),
            .in1(_gnd_net_),
            .in2(N__22440),
            .in3(N__41887),
            .lcout(\c0.n3_adj_2181 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i18_LC_6_29_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i18_LC_6_29_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i18_LC_6_29_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i18_LC_6_29_0  (
            .in0(_gnd_net_),
            .in1(N__22425),
            .in2(_gnd_net_),
            .in3(N__33187),
            .lcout(\c0.FRAME_MATCHER_i_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49766),
            .ce(),
            .sr(N__25449));
    defparam \c0.FRAME_MATCHER_i_i27_LC_6_30_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i27_LC_6_30_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i27_LC_6_30_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i27_LC_6_30_0  (
            .in0(N__33233),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22707),
            .lcout(\c0.FRAME_MATCHER_i_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49778),
            .ce(),
            .sr(N__22659));
    defparam \c0.FRAME_MATCHER_i_i9_LC_6_31_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i9_LC_6_31_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i9_LC_6_31_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i9_LC_6_31_0  (
            .in0(_gnd_net_),
            .in1(N__33234),
            .in2(_gnd_net_),
            .in3(N__22644),
            .lcout(\c0.FRAME_MATCHER_i_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49788),
            .ce(),
            .sr(N__22599));
    defparam \c0.rx.i15081_4_lut_LC_6_32_0 .C_ON=1'b0;
    defparam \c0.rx.i15081_4_lut_LC_6_32_0 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i15081_4_lut_LC_6_32_0 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \c0.rx.i15081_4_lut_LC_6_32_0  (
            .in0(N__31891),
            .in1(N__31853),
            .in2(N__31695),
            .in3(N__31939),
            .lcout(\c0.rx.n17636 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i15113_3_lut_LC_6_32_1 .C_ON=1'b0;
    defparam \c0.rx.i15113_3_lut_LC_6_32_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i15113_3_lut_LC_6_32_1 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \c0.rx.i15113_3_lut_LC_6_32_1  (
            .in0(N__22853),
            .in1(N__25508),
            .in2(_gnd_net_),
            .in3(N__45263),
            .lcout(n17707),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_4_lut_LC_6_32_2 .C_ON=1'b0;
    defparam \c0.rx.i1_4_lut_LC_6_32_2 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_4_lut_LC_6_32_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.rx.i1_4_lut_LC_6_32_2  (
            .in0(N__22575),
            .in1(N__22560),
            .in2(N__22545),
            .in3(N__22527),
            .lcout(\c0.rx.n17022 ),
            .ltout(\c0.rx.n17022_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_3_lut_4_lut_LC_6_32_3 .C_ON=1'b0;
    defparam \c0.rx.i2_3_lut_4_lut_LC_6_32_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_3_lut_4_lut_LC_6_32_3 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \c0.rx.i2_3_lut_4_lut_LC_6_32_3  (
            .in0(N__31719),
            .in1(N__31937),
            .in2(N__22521),
            .in3(N__31774),
            .lcout(\c0.rx.r_SM_Main_2_N_2094_0 ),
            .ltout(\c0.rx.r_SM_Main_2_N_2094_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i14604_2_lut_3_lut_LC_6_32_4 .C_ON=1'b0;
    defparam \c0.rx.i14604_2_lut_3_lut_LC_6_32_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i14604_2_lut_3_lut_LC_6_32_4 .LUT_INIT=16'b1010111110101010;
    LogicCell40 \c0.rx.i14604_2_lut_3_lut_LC_6_32_4  (
            .in0(N__31938),
            .in1(_gnd_net_),
            .in2(N__22518),
            .in3(N__45261),
            .lcout(),
            .ltout(\c0.rx.n17380_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i15000_4_lut_LC_6_32_5 .C_ON=1'b0;
    defparam \c0.rx.i15000_4_lut_LC_6_32_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i15000_4_lut_LC_6_32_5 .LUT_INIT=16'b0101011101010101;
    LogicCell40 \c0.rx.i15000_4_lut_LC_6_32_5  (
            .in0(N__25507),
            .in1(N__31691),
            .in2(N__22515),
            .in3(N__31890),
            .lcout(\c0.rx.n17635 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i2_2_lut_adj_395_LC_6_32_6 .C_ON=1'b0;
    defparam \c0.rx.i2_2_lut_adj_395_LC_6_32_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i2_2_lut_adj_395_LC_6_32_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.rx.i2_2_lut_adj_395_LC_6_32_6  (
            .in0(_gnd_net_),
            .in1(N__45262),
            .in2(_gnd_net_),
            .in3(N__22852),
            .lcout(\c0.rx.n6_adj_2130 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__6__2279_LC_6_32_7 .C_ON=1'b0;
    defparam \c0.data_in_1__6__2279_LC_6_32_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__6__2279_LC_6_32_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_1__6__2279_LC_6_32_7  (
            .in0(N__39030),
            .in1(N__29679),
            .in2(_gnd_net_),
            .in3(N__26973),
            .lcout(data_in_1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49798),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Data_i2_LC_7_16_1 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Data_i2_LC_7_16_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Data_i2_LC_7_16_1 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \c0.tx2.r_Tx_Data_i2_LC_7_16_1  (
            .in0(N__22833),
            .in1(N__32388),
            .in2(N__22827),
            .in3(N__32260),
            .lcout(\c0.tx2.r_Tx_Data_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49659),
            .ce(N__24264),
            .sr(_gnd_net_));
    defparam \c0.i15080_3_lut_LC_7_17_0 .C_ON=1'b0;
    defparam \c0.i15080_3_lut_LC_7_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.i15080_3_lut_LC_7_17_0 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \c0.i15080_3_lut_LC_7_17_0  (
            .in0(N__39264),
            .in1(N__28612),
            .in2(_gnd_net_),
            .in3(N__28901),
            .lcout(\c0.n17620 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Bit_Index_0__bdd_4_lut_15415_LC_7_17_1 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_0__bdd_4_lut_15415_LC_7_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_Bit_Index_0__bdd_4_lut_15415_LC_7_17_1 .LUT_INIT=16'b1110001011001100;
    LogicCell40 \c0.tx2.r_Bit_Index_0__bdd_4_lut_15415_LC_7_17_1  (
            .in0(N__22794),
            .in1(N__25729),
            .in2(N__22782),
            .in3(N__25771),
            .lcout(),
            .ltout(\c0.tx2.n18082_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.n18082_bdd_4_lut_LC_7_17_2 .C_ON=1'b0;
    defparam \c0.tx2.n18082_bdd_4_lut_LC_7_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.n18082_bdd_4_lut_LC_7_17_2 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.tx2.n18082_bdd_4_lut_LC_7_17_2  (
            .in0(N__25772),
            .in1(N__22764),
            .in2(N__22749),
            .in3(N__22746),
            .lcout(),
            .ltout(\c0.tx2.n18085_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i11130210_i1_3_lut_LC_7_17_3 .C_ON=1'b0;
    defparam \c0.tx2.i11130210_i1_3_lut_LC_7_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i11130210_i1_3_lut_LC_7_17_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \c0.tx2.i11130210_i1_3_lut_LC_7_17_3  (
            .in0(N__22868),
            .in1(_gnd_net_),
            .in2(N__22731),
            .in3(N__22728),
            .lcout(),
            .ltout(\c0.tx2.o_Tx_Serial_N_2062_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_2__I_0_56_i3_3_lut_LC_7_17_4 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_2__I_0_56_i3_3_lut_LC_7_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.r_SM_Main_2__I_0_56_i3_3_lut_LC_7_17_4 .LUT_INIT=16'b1100110011110011;
    LogicCell40 \c0.tx2.r_SM_Main_2__I_0_56_i3_3_lut_LC_7_17_4  (
            .in0(_gnd_net_),
            .in1(N__26751),
            .in2(N__22722),
            .in3(N__25936),
            .lcout(n3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i2_2_lut_3_lut_LC_7_17_6 .C_ON=1'b0;
    defparam \c0.tx2.i2_2_lut_3_lut_LC_7_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i2_2_lut_3_lut_LC_7_17_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.tx2.i2_2_lut_3_lut_LC_7_17_6  (
            .in0(N__25730),
            .in1(N__22867),
            .in2(_gnd_net_),
            .in3(N__25773),
            .lcout(\c0.tx2.n13614 ),
            .ltout(\c0.tx2.n13614_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i5661_4_lut_LC_7_17_7 .C_ON=1'b0;
    defparam \c0.tx2.i5661_4_lut_LC_7_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i5661_4_lut_LC_7_17_7 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \c0.tx2.i5661_4_lut_LC_7_17_7  (
            .in0(N__26752),
            .in1(N__35610),
            .in2(N__23064),
            .in3(N__25983),
            .lcout(n8191),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Bit_Index_i0_LC_7_18_0 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_i0_LC_7_18_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Bit_Index_i0_LC_7_18_0 .LUT_INIT=16'b1001100100000000;
    LogicCell40 \c0.tx2.r_Bit_Index_i0_LC_7_18_0  (
            .in0(N__25734),
            .in1(N__24673),
            .in2(_gnd_net_),
            .in3(N__22880),
            .lcout(r_Bit_Index_0_adj_2442),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49660),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15074_3_lut_LC_7_18_1 .C_ON=1'b0;
    defparam \c0.i15074_3_lut_LC_7_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.i15074_3_lut_LC_7_18_1 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \c0.i15074_3_lut_LC_7_18_1  (
            .in0(N__28934),
            .in1(N__28448),
            .in2(_gnd_net_),
            .in3(N__40286),
            .lcout(\c0.n17587 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Bit_Index_i1_LC_7_18_2 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_i1_LC_7_18_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Bit_Index_i1_LC_7_18_2 .LUT_INIT=16'b1101001000000000;
    LogicCell40 \c0.tx2.r_Bit_Index_i1_LC_7_18_2  (
            .in0(N__25735),
            .in1(N__24674),
            .in2(N__25792),
            .in3(N__22881),
            .lcout(r_Bit_Index_1_adj_2441),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49660),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_612_LC_7_18_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_612_LC_7_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_612_LC_7_18_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_612_LC_7_18_3  (
            .in0(_gnd_net_),
            .in1(N__39259),
            .in2(_gnd_net_),
            .in3(N__34710),
            .lcout(\c0.n17107 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15326_LC_7_18_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15326_LC_7_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15326_LC_7_18_4 .LUT_INIT=16'b1111010110001000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15326_LC_7_18_4  (
            .in0(N__28447),
            .in1(N__24527),
            .in2(N__23023),
            .in3(N__28933),
            .lcout(),
            .ltout(\c0.n18118_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18118_bdd_4_lut_LC_7_18_5 .C_ON=1'b0;
    defparam \c0.n18118_bdd_4_lut_LC_7_18_5 .SEQ_MODE=4'b0000;
    defparam \c0.n18118_bdd_4_lut_LC_7_18_5 .LUT_INIT=16'b1111001011000010;
    LogicCell40 \c0.n18118_bdd_4_lut_LC_7_18_5  (
            .in0(N__22974),
            .in1(N__28449),
            .in2(N__22941),
            .in3(N__22938),
            .lcout(\c0.n18121 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i14643_3_lut_LC_7_18_6 .C_ON=1'b0;
    defparam \c0.tx2.i14643_3_lut_LC_7_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i14643_3_lut_LC_7_18_6 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \c0.tx2.i14643_3_lut_LC_7_18_6  (
            .in0(N__26746),
            .in1(N__22890),
            .in2(_gnd_net_),
            .in3(N__24672),
            .lcout(n10976),
            .ltout(n10976_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Bit_Index_i2_LC_7_18_7 .C_ON=1'b0;
    defparam \c0.tx2.r_Bit_Index_i2_LC_7_18_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Bit_Index_i2_LC_7_18_7 .LUT_INIT=16'b1101000000100000;
    LogicCell40 \c0.tx2.r_Bit_Index_i2_LC_7_18_7  (
            .in0(N__25701),
            .in1(N__24675),
            .in2(N__22872),
            .in3(N__22869),
            .lcout(r_Bit_Index_2_adj_2440),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49660),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_1_i6_4_lut_LC_7_19_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_1_i6_4_lut_LC_7_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_1_i6_4_lut_LC_7_19_0 .LUT_INIT=16'b1100110010100000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_1_i6_4_lut_LC_7_19_0  (
            .in0(N__28925),
            .in1(N__23268),
            .in2(N__23388),
            .in3(N__28497),
            .lcout(\c0.n6_adj_2142 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18064_bdd_4_lut_LC_7_19_1 .C_ON=1'b0;
    defparam \c0.n18064_bdd_4_lut_LC_7_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.n18064_bdd_4_lut_LC_7_19_1 .LUT_INIT=16'b1101100111001000;
    LogicCell40 \c0.n18064_bdd_4_lut_LC_7_19_1  (
            .in0(N__28498),
            .in1(N__23337),
            .in2(N__24654),
            .in3(N__24850),
            .lcout(\c0.n18067 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_i0_LC_7_19_2 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_i0_LC_7_19_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_SM_Main_i0_LC_7_19_2 .LUT_INIT=16'b0000001000001110;
    LogicCell40 \c0.tx2.r_SM_Main_i0_LC_7_19_2  (
            .in0(N__23316),
            .in1(N__25939),
            .in2(N__26848),
            .in3(N__25984),
            .lcout(r_SM_Main_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49667),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_1_i5_3_lut_LC_7_19_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_1_i5_3_lut_LC_7_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_1_i5_3_lut_LC_7_19_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_1_i5_3_lut_LC_7_19_4  (
            .in0(N__28924),
            .in1(_gnd_net_),
            .in2(N__26639),
            .in3(N__23307),
            .lcout(\c0.n5_adj_2289 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_593_LC_7_19_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_593_LC_7_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_593_LC_7_19_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_593_LC_7_19_5  (
            .in0(N__26032),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23262),
            .lcout(),
            .ltout(\c0.n10413_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_653_LC_7_19_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_653_LC_7_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_653_LC_7_19_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_653_LC_7_19_6  (
            .in0(N__24137),
            .in1(N__23554),
            .in2(N__23211),
            .in3(N__23621),
            .lcout(\c0.n17282 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15331_LC_7_19_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15331_LC_7_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15331_LC_7_19_7 .LUT_INIT=16'b1110110000101100;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15331_LC_7_19_7  (
            .in0(N__23180),
            .in1(N__28923),
            .in2(N__28600),
            .in3(N__23136),
            .lcout(\c0.n18124 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i100_LC_7_20_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i100_LC_7_20_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i100_LC_7_20_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i100_LC_7_20_0  (
            .in0(N__30171),
            .in1(N__23547),
            .in2(_gnd_net_),
            .in3(N__26585),
            .lcout(data_out_frame2_12_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49675),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15395_LC_7_20_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15395_LC_7_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15395_LC_7_20_1 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15395_LC_7_20_1  (
            .in0(N__28998),
            .in1(N__23097),
            .in2(N__28601),
            .in3(N__23084),
            .lcout(\c0.n18160 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_509_LC_7_20_2 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_509_LC_7_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_509_LC_7_20_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i12_4_lut_adj_509_LC_7_20_2  (
            .in0(N__40896),
            .in1(N__23762),
            .in2(N__23748),
            .in3(N__23687),
            .lcout(\c0.n31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18016_bdd_4_lut_LC_7_20_3 .C_ON=1'b0;
    defparam \c0.n18016_bdd_4_lut_LC_7_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.n18016_bdd_4_lut_LC_7_20_3 .LUT_INIT=16'b1101100111001000;
    LogicCell40 \c0.n18016_bdd_4_lut_LC_7_20_3  (
            .in0(N__28503),
            .in1(N__23931),
            .in2(N__23653),
            .in3(N__23614),
            .lcout(\c0.n18019 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_735_LC_7_20_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_735_LC_7_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_735_LC_7_20_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_735_LC_7_20_4  (
            .in0(N__23503),
            .in1(N__23546),
            .in2(_gnd_net_),
            .in3(N__23475),
            .lcout(\c0.n6_adj_2197 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i72_LC_7_20_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i72_LC_7_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i72_LC_7_20_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \c0.data_out_frame2_0___i72_LC_7_20_5  (
            .in0(N__26584),
            .in1(_gnd_net_),
            .in2(N__23483),
            .in3(N__29929),
            .lcout(data_out_frame2_8_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49675),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i44_LC_7_20_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i44_LC_7_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i44_LC_7_20_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_out_frame2_0___i44_LC_7_20_6  (
            .in0(N__23504),
            .in1(N__31622),
            .in2(_gnd_net_),
            .in3(N__26586),
            .lcout(data_out_frame2_5_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49675),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18142_bdd_4_lut_LC_7_20_7 .C_ON=1'b0;
    defparam \c0.n18142_bdd_4_lut_LC_7_20_7 .SEQ_MODE=4'b0000;
    defparam \c0.n18142_bdd_4_lut_LC_7_20_7 .LUT_INIT=16'b1101110010011000;
    LogicCell40 \c0.n18142_bdd_4_lut_LC_7_20_7  (
            .in0(N__28499),
            .in1(N__23490),
            .in2(N__23482),
            .in3(N__23454),
            .lcout(\c0.n18145 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i114_LC_7_21_0 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i114_LC_7_21_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i114_LC_7_21_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i114_LC_7_21_0  (
            .in0(N__30359),
            .in1(N__23992),
            .in2(_gnd_net_),
            .in3(N__26511),
            .lcout(data_out_frame2_14_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49687),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i15179_4_lut_4_lut_LC_7_21_1 .C_ON=1'b0;
    defparam \c0.tx2.i15179_4_lut_4_lut_LC_7_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i15179_4_lut_4_lut_LC_7_21_1 .LUT_INIT=16'b1001100000010000;
    LogicCell40 \c0.tx2.i15179_4_lut_4_lut_LC_7_21_1  (
            .in0(N__25934),
            .in1(N__26750),
            .in2(N__35605),
            .in3(N__25968),
            .lcout(n4_adj_2484),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i2_3_lut_4_lut_LC_7_21_2 .C_ON=1'b0;
    defparam \c0.tx2.i2_3_lut_4_lut_LC_7_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i2_3_lut_4_lut_LC_7_21_2 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \c0.tx2.i2_3_lut_4_lut_LC_7_21_2  (
            .in0(N__35595),
            .in1(N__26847),
            .in2(N__26754),
            .in3(N__25935),
            .lcout(\c0.tx2.n9269 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i132_LC_7_21_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i132_LC_7_21_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i132_LC_7_21_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i132_LC_7_21_3  (
            .in0(N__26509),
            .in1(N__30170),
            .in2(_gnd_net_),
            .in3(N__24464),
            .lcout(data_out_frame2_16_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49687),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_511_LC_7_21_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_511_LC_7_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_511_LC_7_21_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_511_LC_7_21_4  (
            .in0(N__24156),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24129),
            .lcout(\c0.n10456 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i86_LC_7_21_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i86_LC_7_21_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i86_LC_7_21_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_frame2_0___i86_LC_7_21_5  (
            .in0(N__26510),
            .in1(N__31095),
            .in2(_gnd_net_),
            .in3(N__24063),
            .lcout(data_out_frame2_10_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49687),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i92_LC_7_21_6 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i92_LC_7_21_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i92_LC_7_21_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i92_LC_7_21_6  (
            .in0(N__30716),
            .in1(N__24031),
            .in2(_gnd_net_),
            .in3(N__26512),
            .lcout(data_out_frame2_11_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49687),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i117_LC_7_21_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i117_LC_7_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i117_LC_7_21_7 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \c0.data_out_frame2_0___i117_LC_7_21_7  (
            .in0(N__26508),
            .in1(_gnd_net_),
            .in2(N__31155),
            .in3(N__24778),
            .lcout(data_out_frame2_14_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49687),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15245_LC_7_22_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15245_LC_7_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_0__bdd_4_lut_15245_LC_7_22_0 .LUT_INIT=16'b1111100000111000;
    LogicCell40 \c0.byte_transmit_counter2_0__bdd_4_lut_15245_LC_7_22_0  (
            .in0(N__23985),
            .in1(N__28493),
            .in2(N__29066),
            .in3(N__23964),
            .lcout(\c0.n18016 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_681_LC_7_22_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_681_LC_7_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_681_LC_7_22_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_681_LC_7_22_2  (
            .in0(N__24315),
            .in1(N__23910),
            .in2(_gnd_net_),
            .in3(N__24357),
            .lcout(\c0.n17098 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_2_i5_3_lut_LC_7_22_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_2_i5_3_lut_LC_7_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter2_4__I_0_Mux_2_i5_3_lut_LC_7_22_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter2_4__I_0_Mux_2_i5_3_lut_LC_7_22_3  (
            .in0(N__28997),
            .in1(N__23852),
            .in2(_gnd_net_),
            .in3(N__23819),
            .lcout(\c0.n5_adj_2290 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_429_LC_7_22_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_429_LC_7_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_429_LC_7_22_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_429_LC_7_22_4  (
            .in0(_gnd_net_),
            .in1(N__24774),
            .in2(_gnd_net_),
            .in3(N__24749),
            .lcout(\c0.n17276 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i14635_3_lut_4_lut_LC_7_22_5 .C_ON=1'b0;
    defparam \c0.tx2.i14635_3_lut_4_lut_LC_7_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i14635_3_lut_4_lut_LC_7_22_5 .LUT_INIT=16'b1110111011111110;
    LogicCell40 \c0.tx2.i14635_3_lut_4_lut_LC_7_22_5  (
            .in0(N__25940),
            .in1(N__26840),
            .in2(N__26753),
            .in3(N__25962),
            .lcout(n17412),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_474_LC_7_22_6 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_474_LC_7_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_474_LC_7_22_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_474_LC_7_22_6  (
            .in0(N__24651),
            .in1(N__24609),
            .in2(N__27657),
            .in3(N__24597),
            .lcout(\c0.n17123 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_606_LC_7_22_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_606_LC_7_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_606_LC_7_22_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_606_LC_7_22_7  (
            .in0(_gnd_net_),
            .in1(N__26042),
            .in2(_gnd_net_),
            .in3(N__24525),
            .lcout(\c0.n10434 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_533_LC_7_23_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_533_LC_7_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_533_LC_7_23_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_533_LC_7_23_0  (
            .in0(_gnd_net_),
            .in1(N__24471),
            .in2(_gnd_net_),
            .in3(N__24435),
            .lcout(\c0.n10482 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_584_LC_7_23_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_584_LC_7_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_584_LC_7_23_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_584_LC_7_23_1  (
            .in0(N__24350),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24308),
            .lcout(\c0.n10513 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_514_LC_7_23_2 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_514_LC_7_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_514_LC_7_23_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_514_LC_7_23_2  (
            .in0(N__42192),
            .in1(N__45495),
            .in2(N__46647),
            .in3(N__48883),
            .lcout(\c0.n17110 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_219_Select_12_i3_2_lut_3_lut_LC_7_23_3 .C_ON=1'b0;
    defparam \c0.select_219_Select_12_i3_2_lut_3_lut_LC_7_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.select_219_Select_12_i3_2_lut_3_lut_LC_7_23_3 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \c0.select_219_Select_12_i3_2_lut_3_lut_LC_7_23_3  (
            .in0(N__27834),
            .in1(N__25866),
            .in2(_gnd_net_),
            .in3(N__41765),
            .lcout(\c0.n3_adj_2268 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__2__2267_LC_7_23_4 .C_ON=1'b0;
    defparam \c0.data_in_3__2__2267_LC_7_23_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__2__2267_LC_7_23_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_3__2__2267_LC_7_23_4  (
            .in0(N__39221),
            .in1(N__36881),
            .in2(_gnd_net_),
            .in3(N__38967),
            .lcout(data_in_3_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49709),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_597_LC_7_23_5 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_597_LC_7_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_597_LC_7_23_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i7_4_lut_adj_597_LC_7_23_5  (
            .in0(N__27579),
            .in1(N__24936),
            .in2(N__24869),
            .in3(N__24851),
            .lcout(\c0.n17_adj_2321 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__6__2271_LC_7_23_6 .C_ON=1'b0;
    defparam \c0.data_in_2__6__2271_LC_7_23_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__6__2271_LC_7_23_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_2__6__2271_LC_7_23_6  (
            .in0(N__39220),
            .in1(N__35094),
            .in2(_gnd_net_),
            .in3(N__26962),
            .lcout(data_in_2_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49709),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i19_LC_7_24_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i19_LC_7_24_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i19_LC_7_24_0 .LUT_INIT=16'b1110000011000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i19_LC_7_24_0  (
            .in0(N__44990),
            .in1(N__44777),
            .in2(N__27430),
            .in3(N__44602),
            .lcout(\c0.FRAME_MATCHER_state_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49722),
            .ce(),
            .sr(N__27408));
    defparam \c0.FRAME_MATCHER_state_i12_LC_7_25_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i12_LC_7_25_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i12_LC_7_25_0 .LUT_INIT=16'b1010101010000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i12_LC_7_25_0  (
            .in0(N__27347),
            .in1(N__44991),
            .in2(N__44618),
            .in3(N__44799),
            .lcout(\c0.FRAME_MATCHER_state_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49732),
            .ce(),
            .sr(N__27333));
    defparam \c0.i1_2_lut_adj_410_LC_7_25_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_410_LC_7_25_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_410_LC_7_25_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i1_2_lut_adj_410_LC_7_25_1  (
            .in0(_gnd_net_),
            .in1(N__33322),
            .in2(_gnd_net_),
            .in3(N__27346),
            .lcout(),
            .ltout(\c0.n30_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i22_4_lut_LC_7_25_2 .C_ON=1'b0;
    defparam \c0.i22_4_lut_LC_7_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.i22_4_lut_LC_7_25_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i22_4_lut_LC_7_25_2  (
            .in0(N__29609),
            .in1(N__27323),
            .in2(N__24786),
            .in3(N__27391),
            .lcout(\c0.n51 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15142_3_lut_LC_7_25_3 .C_ON=1'b0;
    defparam \c0.i15142_3_lut_LC_7_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.i15142_3_lut_LC_7_25_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \c0.i15142_3_lut_LC_7_25_3  (
            .in0(N__48421),
            .in1(N__42492),
            .in2(_gnd_net_),
            .in3(N__44287),
            .lcout(\c0.n17574 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15001_3_lut_LC_7_25_4 .C_ON=1'b0;
    defparam \c0.i15001_3_lut_LC_7_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.i15001_3_lut_LC_7_25_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \c0.i15001_3_lut_LC_7_25_4  (
            .in0(N__48419),
            .in1(N__47133),
            .in2(_gnd_net_),
            .in3(N__49109),
            .lcout(\c0.n17643 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15002_3_lut_LC_7_25_7 .C_ON=1'b0;
    defparam \c0.i15002_3_lut_LC_7_25_7 .SEQ_MODE=4'b0000;
    defparam \c0.i15002_3_lut_LC_7_25_7 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \c0.i15002_3_lut_LC_7_25_7  (
            .in0(N__49110),
            .in1(N__48420),
            .in2(_gnd_net_),
            .in3(N__44286),
            .lcout(\c0.n17647 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i8_LC_7_26_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i8_LC_7_26_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i8_LC_7_26_0 .LUT_INIT=16'b1110000011000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i8_LC_7_26_0  (
            .in0(N__44992),
            .in1(N__44800),
            .in2(N__33332),
            .in3(N__44610),
            .lcout(\c0.FRAME_MATCHER_state_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49743),
            .ce(),
            .sr(N__33306));
    defparam \c0.i10662_2_lut_LC_7_26_1 .C_ON=1'b0;
    defparam \c0.i10662_2_lut_LC_7_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.i10662_2_lut_LC_7_26_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i10662_2_lut_LC_7_26_1  (
            .in0(_gnd_net_),
            .in1(N__25299),
            .in2(_gnd_net_),
            .in3(N__41836),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10663_2_lut_LC_7_26_2 .C_ON=1'b0;
    defparam \c0.i10663_2_lut_LC_7_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.i10663_2_lut_LC_7_26_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i10663_2_lut_LC_7_26_2  (
            .in0(N__41837),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25220),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10664_2_lut_LC_7_26_3 .C_ON=1'b0;
    defparam \c0.i10664_2_lut_LC_7_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.i10664_2_lut_LC_7_26_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i10664_2_lut_LC_7_26_3  (
            .in0(_gnd_net_),
            .in1(N__25169),
            .in2(_gnd_net_),
            .in3(N__41838),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10665_2_lut_LC_7_26_4 .C_ON=1'b0;
    defparam \c0.i10665_2_lut_LC_7_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.i10665_2_lut_LC_7_26_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i10665_2_lut_LC_7_26_4  (
            .in0(N__41839),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25125),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10668_2_lut_LC_7_26_5 .C_ON=1'b0;
    defparam \c0.i10668_2_lut_LC_7_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.i10668_2_lut_LC_7_26_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i10668_2_lut_LC_7_26_5  (
            .in0(N__25053),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41840),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10669_2_lut_LC_7_26_6 .C_ON=1'b0;
    defparam \c0.i10669_2_lut_LC_7_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.i10669_2_lut_LC_7_26_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i10669_2_lut_LC_7_26_6  (
            .in0(N__41841),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25007),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10672_2_lut_LC_7_26_7 .C_ON=1'b0;
    defparam \c0.i10672_2_lut_LC_7_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.i10672_2_lut_LC_7_26_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i10672_2_lut_LC_7_26_7  (
            .in0(_gnd_net_),
            .in1(N__27889),
            .in2(_gnd_net_),
            .in3(N__41842),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i5_LC_7_27_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i5_LC_7_27_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i5_LC_7_27_0 .LUT_INIT=16'b1110000011000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i5_LC_7_27_0  (
            .in0(N__45020),
            .in1(N__44801),
            .in2(N__33469),
            .in3(N__44606),
            .lcout(\c0.FRAME_MATCHER_state_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49754),
            .ce(),
            .sr(N__29475));
    defparam \c0.select_219_Select_18_i3_2_lut_3_lut_LC_7_27_1 .C_ON=1'b0;
    defparam \c0.select_219_Select_18_i3_2_lut_3_lut_LC_7_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.select_219_Select_18_i3_2_lut_3_lut_LC_7_27_1 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \c0.select_219_Select_18_i3_2_lut_3_lut_LC_7_27_1  (
            .in0(N__41851),
            .in1(_gnd_net_),
            .in2(N__25437),
            .in3(N__27819),
            .lcout(\c0.n3_adj_2254 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10670_2_lut_LC_7_27_2 .C_ON=1'b0;
    defparam \c0.i10670_2_lut_LC_7_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.i10670_2_lut_LC_7_27_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i10670_2_lut_LC_7_27_2  (
            .in0(_gnd_net_),
            .in1(N__25433),
            .in2(_gnd_net_),
            .in3(N__41849),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_219_Select_1_i3_2_lut_3_lut_LC_7_27_3 .C_ON=1'b0;
    defparam \c0.select_219_Select_1_i3_2_lut_3_lut_LC_7_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.select_219_Select_1_i3_2_lut_3_lut_LC_7_27_3 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \c0.select_219_Select_1_i3_2_lut_3_lut_LC_7_27_3  (
            .in0(N__41852),
            .in1(_gnd_net_),
            .in2(N__32884),
            .in3(N__27817),
            .lcout(\c0.n3_adj_2288 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10687_2_lut_LC_7_27_4 .C_ON=1'b0;
    defparam \c0.i10687_2_lut_LC_7_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.i10687_2_lut_LC_7_27_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i10687_2_lut_LC_7_27_4  (
            .in0(_gnd_net_),
            .in1(N__32873),
            .in2(_gnd_net_),
            .in3(N__41850),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_219_Select_22_i3_2_lut_3_lut_LC_7_27_5 .C_ON=1'b0;
    defparam \c0.select_219_Select_22_i3_2_lut_3_lut_LC_7_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.select_219_Select_22_i3_2_lut_3_lut_LC_7_27_5 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \c0.select_219_Select_22_i3_2_lut_3_lut_LC_7_27_5  (
            .in0(N__41853),
            .in1(_gnd_net_),
            .in2(N__25347),
            .in3(N__27818),
            .lcout(\c0.n3_adj_2246 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10666_2_lut_LC_7_27_6 .C_ON=1'b0;
    defparam \c0.i10666_2_lut_LC_7_27_6 .SEQ_MODE=4'b0000;
    defparam \c0.i10666_2_lut_LC_7_27_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i10666_2_lut_LC_7_27_6  (
            .in0(_gnd_net_),
            .in1(N__25343),
            .in2(_gnd_net_),
            .in3(N__41848),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_219_Select_26_i3_2_lut_3_lut_LC_7_27_7 .C_ON=1'b0;
    defparam \c0.select_219_Select_26_i3_2_lut_3_lut_LC_7_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.select_219_Select_26_i3_2_lut_3_lut_LC_7_27_7 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \c0.select_219_Select_26_i3_2_lut_3_lut_LC_7_27_7  (
            .in0(N__41854),
            .in1(N__27816),
            .in2(_gnd_net_),
            .in3(N__25298),
            .lcout(\c0.n3_adj_2238 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i10_LC_7_28_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i10_LC_7_28_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i10_LC_7_28_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i10_LC_7_28_0  (
            .in0(_gnd_net_),
            .in1(N__25242),
            .in2(_gnd_net_),
            .in3(N__33184),
            .lcout(\c0.FRAME_MATCHER_i_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49767),
            .ce(),
            .sr(N__28017));
    defparam \c0.FRAME_MATCHER_state_i14_LC_7_29_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i14_LC_7_29_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i14_LC_7_29_0 .LUT_INIT=16'b1110000011000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i14_LC_7_29_0  (
            .in0(N__45021),
            .in1(N__44812),
            .in2(N__27322),
            .in3(N__44615),
            .lcout(\c0.FRAME_MATCHER_state_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49779),
            .ce(),
            .sr(N__27297));
    defparam \c0.tx2.i2615_2_lut_LC_7_29_2 .C_ON=1'b0;
    defparam \c0.tx2.i2615_2_lut_LC_7_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i2615_2_lut_LC_7_29_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.tx2.i2615_2_lut_LC_7_29_2  (
            .in0(_gnd_net_),
            .in1(N__25793),
            .in2(_gnd_net_),
            .in3(N__25740),
            .lcout(n5266),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.o_Tx_Serial_I_0_1_lut_LC_7_29_3 .C_ON=1'b0;
    defparam \c0.tx.o_Tx_Serial_I_0_1_lut_LC_7_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx.o_Tx_Serial_I_0_1_lut_LC_7_29_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \c0.tx.o_Tx_Serial_I_0_1_lut_LC_7_29_3  (
            .in0(N__43880),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(tx_enable),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.i1_1_lut_LC_7_29_4 .C_ON=1'b0;
    defparam \c0.tx2.i1_1_lut_LC_7_29_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx2.i1_1_lut_LC_7_29_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \c0.tx2.i1_1_lut_LC_7_29_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26853),
            .lcout(n10674),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__1__2199_LC_7_30_0 .C_ON=1'b0;
    defparam \c0.data_out_7__1__2199_LC_7_30_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__1__2199_LC_7_30_0 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \c0.data_out_7__1__2199_LC_7_30_0  (
            .in0(N__25647),
            .in1(N__48089),
            .in2(N__50321),
            .in3(N__29757),
            .lcout(\c0.data_out_7_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49789),
            .ce(N__46933),
            .sr(_gnd_net_));
    defparam \c0.i15053_2_lut_LC_7_30_2 .C_ON=1'b0;
    defparam \c0.i15053_2_lut_LC_7_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.i15053_2_lut_LC_7_30_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i15053_2_lut_LC_7_30_2  (
            .in0(N__30303),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48088),
            .lcout(\c0.n17626 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i13_4_lut_4_lut_LC_7_30_4 .C_ON=1'b0;
    defparam \c0.rx.i13_4_lut_4_lut_LC_7_30_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i13_4_lut_4_lut_LC_7_30_4 .LUT_INIT=16'b0100000000001111;
    LogicCell40 \c0.rx.i13_4_lut_4_lut_LC_7_30_4  (
            .in0(N__31850),
            .in1(N__25584),
            .in2(N__25509),
            .in3(N__25563),
            .lcout(\c0.rx.n10620 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i14585_4_lut_LC_7_30_5 .C_ON=1'b0;
    defparam \c0.rx.i14585_4_lut_LC_7_30_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i14585_4_lut_LC_7_30_5 .LUT_INIT=16'b1111111111001110;
    LogicCell40 \c0.rx.i14585_4_lut_LC_7_30_5  (
            .in0(N__25561),
            .in1(N__25503),
            .in2(N__25591),
            .in3(N__31849),
            .lcout(n17361),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_3_lut_4_lut_LC_7_30_6 .C_ON=1'b0;
    defparam \c0.rx.i1_3_lut_4_lut_LC_7_30_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_3_lut_4_lut_LC_7_30_6 .LUT_INIT=16'b1111111011101110;
    LogicCell40 \c0.rx.i1_3_lut_4_lut_LC_7_30_6  (
            .in0(N__31775),
            .in1(N__31735),
            .in2(N__31952),
            .in3(N__31895),
            .lcout(\c0.rx.r_SM_Main_2_N_2088_2 ),
            .ltout(\c0.rx.r_SM_Main_2_N_2088_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i3_4_lut_LC_7_30_7 .C_ON=1'b0;
    defparam \c0.rx.i3_4_lut_LC_7_30_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i3_4_lut_LC_7_30_7 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \c0.rx.i3_4_lut_LC_7_30_7  (
            .in0(N__25562),
            .in1(N__31848),
            .in2(N__25512),
            .in3(N__25502),
            .lcout(\c0.rx.n10158 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i12_LC_7_31_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i12_LC_7_31_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i12_LC_7_31_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i12_LC_7_31_0  (
            .in0(_gnd_net_),
            .in1(N__25884),
            .in2(_gnd_net_),
            .in3(N__33232),
            .lcout(\c0.FRAME_MATCHER_i_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49799),
            .ce(),
            .sr(N__25833));
    defparam \c0.FRAME_MATCHER_state_i20_LC_7_32_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i20_LC_7_32_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i20_LC_7_32_0 .LUT_INIT=16'b1110110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i20_LC_7_32_0  (
            .in0(N__45032),
            .in1(N__44813),
            .in2(N__44619),
            .in3(N__29608),
            .lcout(\c0.FRAME_MATCHER_state_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49806),
            .ce(),
            .sr(N__29586));
    defparam \c0.byte_transmit_counter2_i4_LC_9_16_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_i4_LC_9_16_0 .SEQ_MODE=4'b1001;
    defparam \c0.byte_transmit_counter2_i4_LC_9_16_0 .LUT_INIT=16'b1100101000000000;
    LogicCell40 \c0.byte_transmit_counter2_i4_LC_9_16_0  (
            .in0(N__25806),
            .in1(N__32234),
            .in2(N__39683),
            .in3(N__42086),
            .lcout(\c0.byte_transmit_counter2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49676),
            .ce(),
            .sr(N__26922));
    defparam \c0.add_2510_2_lut_LC_9_17_0 .C_ON=1'b1;
    defparam \c0.add_2510_2_lut_LC_9_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.add_2510_2_lut_LC_9_17_0 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.add_2510_2_lut_LC_9_17_0  (
            .in0(N__34110),
            .in1(N__28783),
            .in2(_gnd_net_),
            .in3(N__25818),
            .lcout(\c0.n17659 ),
            .ltout(),
            .carryin(bfn_9_17_0_),
            .carryout(\c0.n15972 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2510_3_lut_LC_9_17_1 .C_ON=1'b1;
    defparam \c0.add_2510_3_lut_LC_9_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_2510_3_lut_LC_9_17_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.add_2510_3_lut_LC_9_17_1  (
            .in0(N__34112),
            .in1(N__28465),
            .in2(_gnd_net_),
            .in3(N__25815),
            .lcout(\c0.n17589 ),
            .ltout(),
            .carryin(\c0.n15972 ),
            .carryout(\c0.n15973 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2510_4_lut_LC_9_17_2 .C_ON=1'b1;
    defparam \c0.add_2510_4_lut_LC_9_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_2510_4_lut_LC_9_17_2 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.add_2510_4_lut_LC_9_17_2  (
            .in0(N__34108),
            .in1(N__32109),
            .in2(_gnd_net_),
            .in3(N__25812),
            .lcout(\c0.n17710 ),
            .ltout(),
            .carryin(\c0.n15973 ),
            .carryout(\c0.n15974 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2510_5_lut_LC_9_17_3 .C_ON=1'b1;
    defparam \c0.add_2510_5_lut_LC_9_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_2510_5_lut_LC_9_17_3 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.add_2510_5_lut_LC_9_17_3  (
            .in0(N__34113),
            .in1(N__32334),
            .in2(_gnd_net_),
            .in3(N__25809),
            .lcout(\c0.n17711 ),
            .ltout(),
            .carryin(\c0.n15974 ),
            .carryout(\c0.n15975 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2510_6_lut_LC_9_17_4 .C_ON=1'b1;
    defparam \c0.add_2510_6_lut_LC_9_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_2510_6_lut_LC_9_17_4 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.add_2510_6_lut_LC_9_17_4  (
            .in0(N__34109),
            .in1(N__32225),
            .in2(_gnd_net_),
            .in3(N__25800),
            .lcout(\c0.n17606 ),
            .ltout(),
            .carryin(\c0.n15975 ),
            .carryout(\c0.n15976 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2510_7_lut_LC_9_17_5 .C_ON=1'b1;
    defparam \c0.add_2510_7_lut_LC_9_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_2510_7_lut_LC_9_17_5 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.add_2510_7_lut_LC_9_17_5  (
            .in0(N__34111),
            .in1(N__39623),
            .in2(_gnd_net_),
            .in3(N__25797),
            .lcout(\c0.n17712 ),
            .ltout(),
            .carryin(\c0.n15976 ),
            .carryout(\c0.n15977 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2510_8_lut_LC_9_17_6 .C_ON=1'b1;
    defparam \c0.add_2510_8_lut_LC_9_17_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_2510_8_lut_LC_9_17_6 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.add_2510_8_lut_LC_9_17_6  (
            .in0(N__34106),
            .in1(N__34446),
            .in2(_gnd_net_),
            .in3(N__26670),
            .lcout(\c0.n17713 ),
            .ltout(),
            .carryin(\c0.n15977 ),
            .carryout(\c0.n15978 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2510_9_lut_LC_9_17_7 .C_ON=1'b0;
    defparam \c0.add_2510_9_lut_LC_9_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_2510_9_lut_LC_9_17_7 .LUT_INIT=16'b1000010001001000;
    LogicCell40 \c0.add_2510_9_lut_LC_9_17_7  (
            .in0(N__34485),
            .in1(N__34107),
            .in2(_gnd_net_),
            .in3(N__26667),
            .lcout(\c0.n17714 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_i1_LC_9_18_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_i1_LC_9_18_0 .SEQ_MODE=4'b1001;
    defparam \c0.byte_transmit_counter2_i1_LC_9_18_0 .LUT_INIT=16'b1100101000000000;
    LogicCell40 \c0.byte_transmit_counter2_i1_LC_9_18_0  (
            .in0(N__26652),
            .in1(N__28362),
            .in2(N__39679),
            .in3(N__42084),
            .lcout(\c0.byte_transmit_counter2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49677),
            .ce(),
            .sr(N__28263));
    defparam \c0.i1_2_lut_adj_415_LC_9_19_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_415_LC_9_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_415_LC_9_19_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i1_2_lut_adj_415_LC_9_19_0  (
            .in0(_gnd_net_),
            .in1(N__37186),
            .in2(_gnd_net_),
            .in3(N__37105),
            .lcout(\c0.n15179 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i58_LC_9_19_1 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i58_LC_9_19_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i58_LC_9_19_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i58_LC_9_19_1  (
            .in0(N__29817),
            .in1(N__26632),
            .in2(_gnd_net_),
            .in3(N__26612),
            .lcout(data_out_frame2_7_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49688),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__0__2277_LC_9_19_3 .C_ON=1'b0;
    defparam \c0.data_in_2__0__2277_LC_9_19_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__0__2277_LC_9_19_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_2__0__2277_LC_9_19_3  (
            .in0(N__39207),
            .in1(N__29140),
            .in2(_gnd_net_),
            .in3(N__34934),
            .lcout(data_in_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49688),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_i1_LC_9_19_4 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_i1_LC_9_19_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_SM_Main_i1_LC_9_19_4 .LUT_INIT=16'b0000000001111000;
    LogicCell40 \c0.tx2.r_SM_Main_i1_LC_9_19_4  (
            .in0(N__25985),
            .in1(N__25937),
            .in2(N__26741),
            .in3(N__26818),
            .lcout(r_SM_Main_1_adj_2439),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49688),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i97_LC_9_19_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i97_LC_9_19_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i97_LC_9_19_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_frame2_0___i97_LC_9_19_5  (
            .in0(N__29458),
            .in1(N__26022),
            .in2(_gnd_net_),
            .in3(N__26613),
            .lcout(data_out_frame2_12_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49688),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_SM_Main_i2_LC_9_19_6 .C_ON=1'b0;
    defparam \c0.tx2.r_SM_Main_i2_LC_9_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_SM_Main_i2_LC_9_19_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \c0.tx2.r_SM_Main_i2_LC_9_19_6  (
            .in0(N__25986),
            .in1(N__25938),
            .in2(N__26740),
            .in3(N__26819),
            .lcout(r_SM_Main_2_adj_2438),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49688),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_2_lut_3_lut_LC_9_20_0 .C_ON=1'b0;
    defparam \c0.i6_2_lut_3_lut_LC_9_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i6_2_lut_3_lut_LC_9_20_0 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \c0.i6_2_lut_3_lut_LC_9_20_0  (
            .in0(N__48425),
            .in1(N__48167),
            .in2(_gnd_net_),
            .in3(N__50315),
            .lcout(n10705),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14597_3_lut_4_lut_LC_9_20_1 .C_ON=1'b0;
    defparam \c0.i14597_3_lut_4_lut_LC_9_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i14597_3_lut_4_lut_LC_9_20_1 .LUT_INIT=16'b1000001000101000;
    LogicCell40 \c0.i14597_3_lut_4_lut_LC_9_20_1  (
            .in0(N__32514),
            .in1(N__34773),
            .in2(N__35127),
            .in3(N__37398),
            .lcout(\c0.n17373 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i50_LC_9_20_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i50_LC_9_20_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i50_LC_9_20_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0__i50_LC_9_20_2  (
            .in0(N__39479),
            .in1(N__34673),
            .in2(_gnd_net_),
            .in3(N__32562),
            .lcout(data_in_frame_6_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49698),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2.r_Tx_Active_47_LC_9_20_3 .C_ON=1'b0;
    defparam \c0.tx2.r_Tx_Active_47_LC_9_20_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx2.r_Tx_Active_47_LC_9_20_3 .LUT_INIT=16'b1011000011110100;
    LogicCell40 \c0.tx2.r_Tx_Active_47_LC_9_20_3  (
            .in0(N__26826),
            .in1(N__26769),
            .in2(N__34395),
            .in3(N__26720),
            .lcout(tx2_active),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49698),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i55_LC_9_20_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i55_LC_9_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i55_LC_9_20_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_frame_0__i55_LC_9_20_5  (
            .in0(N__32563),
            .in1(N__39553),
            .in2(_gnd_net_),
            .in3(N__36992),
            .lcout(data_in_frame_6_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49698),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i49_LC_9_20_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i49_LC_9_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i49_LC_9_20_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_in_frame_0__i49_LC_9_20_6  (
            .in0(N__34550),
            .in1(N__36801),
            .in2(_gnd_net_),
            .in3(N__32561),
            .lcout(data_in_frame_6_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49698),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__2__2283_LC_9_20_7 .C_ON=1'b0;
    defparam \c0.data_in_1__2__2283_LC_9_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__2__2283_LC_9_20_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_1__2__2283_LC_9_20_7  (
            .in0(N__39206),
            .in1(N__28048),
            .in2(_gnd_net_),
            .in3(N__38940),
            .lcout(data_in_1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49698),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__5__2272_LC_9_21_0 .C_ON=1'b0;
    defparam \c0.data_in_2__5__2272_LC_9_21_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__5__2272_LC_9_21_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_2__5__2272_LC_9_21_0  (
            .in0(N__29180),
            .in1(N__29651),
            .in2(_gnd_net_),
            .in3(N__39211),
            .lcout(data_in_2_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49710),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__3__2290_LC_9_21_1 .C_ON=1'b0;
    defparam \c0.data_in_0__3__2290_LC_9_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__3__2290_LC_9_21_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0__3__2290_LC_9_21_1  (
            .in0(N__26868),
            .in1(N__39095),
            .in2(_gnd_net_),
            .in3(N__26901),
            .lcout(data_in_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49710),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_657_LC_9_21_2 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_657_LC_9_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_657_LC_9_21_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i7_4_lut_adj_657_LC_9_21_2  (
            .in0(N__26900),
            .in1(N__29176),
            .in2(N__29154),
            .in3(N__29280),
            .lcout(\c0.n17_adj_2370 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10774_2_lut_LC_9_21_3 .C_ON=1'b0;
    defparam \c0.i10774_2_lut_LC_9_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i10774_2_lut_LC_9_21_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i10774_2_lut_LC_9_21_3  (
            .in0(_gnd_net_),
            .in1(N__29328),
            .in2(_gnd_net_),
            .in3(N__26899),
            .lcout(\c0.n13450 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__7__2286_LC_9_21_4 .C_ON=1'b0;
    defparam \c0.data_in_0__7__2286_LC_9_21_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__7__2286_LC_9_21_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0__7__2286_LC_9_21_4  (
            .in0(N__29329),
            .in1(N__39212),
            .in2(_gnd_net_),
            .in3(N__26880),
            .lcout(data_in_0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49710),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__3__2274_LC_9_21_5 .C_ON=1'b0;
    defparam \c0.data_in_2__3__2274_LC_9_21_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__3__2274_LC_9_21_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_2__3__2274_LC_9_21_5  (
            .in0(N__39210),
            .in1(N__29213),
            .in2(_gnd_net_),
            .in3(N__35241),
            .lcout(data_in_2_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49710),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__3__2282_LC_9_21_6 .C_ON=1'b0;
    defparam \c0.data_in_1__3__2282_LC_9_21_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__3__2282_LC_9_21_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_1__3__2282_LC_9_21_6  (
            .in0(N__29214),
            .in1(N__39213),
            .in2(_gnd_net_),
            .in3(N__26867),
            .lcout(data_in_1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49710),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__0__2285_LC_9_21_7 .C_ON=1'b0;
    defparam \c0.data_in_1__0__2285_LC_9_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__0__2285_LC_9_21_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_1__0__2285_LC_9_21_7  (
            .in0(N__39209),
            .in1(N__29153),
            .in2(_gnd_net_),
            .in3(N__35051),
            .lcout(data_in_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49710),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_627_LC_9_22_0 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_627_LC_9_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_627_LC_9_22_0 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \c0.i6_4_lut_adj_627_LC_9_22_0  (
            .in0(N__27531),
            .in1(N__26943),
            .in2(N__35009),
            .in3(N__26979),
            .lcout(\c0.n10133 ),
            .ltout(\c0.n10133_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_631_LC_9_22_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_631_LC_9_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_631_LC_9_22_1 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \c0.i1_2_lut_adj_631_LC_9_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26889),
            .in3(N__27277),
            .lcout(),
            .ltout(\c0.n6_adj_2356_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_632_LC_9_22_2 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_632_LC_9_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_632_LC_9_22_2 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \c0.i4_4_lut_adj_632_LC_9_22_2  (
            .in0(N__26907),
            .in1(N__29211),
            .in2(N__26886),
            .in3(N__29232),
            .lcout(\c0.n10027 ),
            .ltout(\c0.n10027_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_642_LC_9_22_3 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_642_LC_9_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_642_LC_9_22_3 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \c0.i3_4_lut_adj_642_LC_9_22_3  (
            .in0(N__35377),
            .in1(N__28029),
            .in2(N__26883),
            .in3(N__29253),
            .lcout(n63_adj_2418),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14556_2_lut_LC_9_22_4 .C_ON=1'b0;
    defparam \c0.i14556_2_lut_LC_9_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i14556_2_lut_LC_9_22_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i14556_2_lut_LC_9_22_4  (
            .in0(_gnd_net_),
            .in1(N__26879),
            .in2(_gnd_net_),
            .in3(N__26866),
            .lcout(),
            .ltout(\c0.n17331_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14633_4_lut_LC_9_22_5 .C_ON=1'b0;
    defparam \c0.i14633_4_lut_LC_9_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i14633_4_lut_LC_9_22_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i14633_4_lut_LC_9_22_5  (
            .in0(N__35050),
            .in1(N__27546),
            .in2(N__26982),
            .in3(N__27516),
            .lcout(\c0.n17410 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__4__2281_LC_9_22_6 .C_ON=1'b0;
    defparam \c0.data_in_1__4__2281_LC_9_22_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__4__2281_LC_9_22_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_1__4__2281_LC_9_22_6  (
            .in0(N__39184),
            .in1(N__26937),
            .in2(_gnd_net_),
            .in3(N__29233),
            .lcout(data_in_1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49723),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_625_LC_9_23_0 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_625_LC_9_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_625_LC_9_23_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i5_4_lut_adj_625_LC_9_23_0  (
            .in0(N__26963),
            .in1(N__35237),
            .in2(N__35405),
            .in3(N__26935),
            .lcout(\c0.n12_adj_2355 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__4__2273_LC_9_23_1 .C_ON=1'b0;
    defparam \c0.data_in_2__4__2273_LC_9_23_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__4__2273_LC_9_23_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_2__4__2273_LC_9_23_1  (
            .in0(N__26936),
            .in1(N__39186),
            .in2(_gnd_net_),
            .in3(N__29733),
            .lcout(data_in_2_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49733),
            .ce(),
            .sr(_gnd_net_));
    defparam i14650_4_lut_LC_9_23_2.C_ON=1'b0;
    defparam i14650_4_lut_LC_9_23_2.SEQ_MODE=4'b0000;
    defparam i14650_4_lut_LC_9_23_2.LUT_INIT=16'b1111001000110000;
    LogicCell40 i14650_4_lut_LC_9_23_2 (
            .in0(N__36245),
            .in1(N__36275),
            .in2(N__36174),
            .in3(N__36203),
            .lcout(n17427),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_414_LC_9_23_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_414_LC_9_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_414_LC_9_23_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i1_2_lut_adj_414_LC_9_23_3  (
            .in0(N__32247),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33537),
            .lcout(\c0.n4_adj_2150 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__1__2276_LC_9_23_4 .C_ON=1'b0;
    defparam \c0.data_in_2__1__2276_LC_9_23_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__1__2276_LC_9_23_4 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \c0.data_in_2__1__2276_LC_9_23_4  (
            .in0(N__35401),
            .in1(_gnd_net_),
            .in2(N__39218),
            .in3(N__35010),
            .lcout(data_in_2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49733),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_646_LC_9_23_5 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_646_LC_9_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_646_LC_9_23_5 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \c0.i7_4_lut_adj_646_LC_9_23_5  (
            .in0(N__29731),
            .in1(N__26913),
            .in2(N__27282),
            .in3(N__27566),
            .lcout(\c0.n17_adj_2362 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14629_4_lut_LC_9_23_6 .C_ON=1'b0;
    defparam \c0.i14629_4_lut_LC_9_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i14629_4_lut_LC_9_23_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i14629_4_lut_LC_9_23_6  (
            .in0(N__38977),
            .in1(N__29730),
            .in2(N__27567),
            .in3(N__34933),
            .lcout(\c0.n17406 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__6__2287_LC_9_23_7 .C_ON=1'b0;
    defparam \c0.data_in_0__6__2287_LC_9_23_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__6__2287_LC_9_23_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_in_0__6__2287_LC_9_23_7  (
            .in0(N__27281),
            .in1(N__39185),
            .in2(_gnd_net_),
            .in3(N__29712),
            .lcout(data_in_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49733),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i9_LC_9_24_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i9_LC_9_24_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i9_LC_9_24_0 .LUT_INIT=16'b1110000011000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i9_LC_9_24_0  (
            .in0(N__44931),
            .in1(N__44776),
            .in2(N__33290),
            .in3(N__44601),
            .lcout(\c0.FRAME_MATCHER_state_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49744),
            .ce(),
            .sr(N__33264));
    defparam \c0.i10673_2_lut_LC_9_24_1 .C_ON=1'b0;
    defparam \c0.i10673_2_lut_LC_9_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.i10673_2_lut_LC_9_24_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i10673_2_lut_LC_9_24_1  (
            .in0(_gnd_net_),
            .in1(N__27264),
            .in2(_gnd_net_),
            .in3(N__41672),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10675_2_lut_LC_9_24_2 .C_ON=1'b0;
    defparam \c0.i10675_2_lut_LC_9_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.i10675_2_lut_LC_9_24_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i10675_2_lut_LC_9_24_2  (
            .in0(N__41673),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27210),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10677_2_lut_LC_9_24_3 .C_ON=1'b0;
    defparam \c0.i10677_2_lut_LC_9_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.i10677_2_lut_LC_9_24_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i10677_2_lut_LC_9_24_3  (
            .in0(_gnd_net_),
            .in1(N__27159),
            .in2(_gnd_net_),
            .in3(N__41674),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10681_2_lut_LC_9_24_4 .C_ON=1'b0;
    defparam \c0.i10681_2_lut_LC_9_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.i10681_2_lut_LC_9_24_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i10681_2_lut_LC_9_24_4  (
            .in0(N__41675),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27099),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_405_LC_9_24_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_405_LC_9_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_405_LC_9_24_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i1_2_lut_adj_405_LC_9_24_5  (
            .in0(N__37175),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41670),
            .lcout(\c0.n37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_701_LC_9_24_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_701_LC_9_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_701_LC_9_24_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i1_2_lut_adj_701_LC_9_24_6  (
            .in0(N__41671),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27033),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15155_2_lut_LC_9_24_7 .C_ON=1'b0;
    defparam \c0.i15155_2_lut_LC_9_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.i15155_2_lut_LC_9_24_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i15155_2_lut_LC_9_24_7  (
            .in0(_gnd_net_),
            .in1(N__36297),
            .in2(_gnd_net_),
            .in3(N__47842),
            .lcout(\c0.n17701 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i21_4_lut_LC_9_25_0 .C_ON=1'b0;
    defparam \c0.i21_4_lut_LC_9_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.i21_4_lut_LC_9_25_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i21_4_lut_LC_9_25_0  (
            .in0(N__27431),
            .in1(N__27482),
            .in2(N__38070),
            .in3(N__27451),
            .lcout(\c0.n50 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i13_LC_9_25_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i13_LC_9_25_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i13_LC_9_25_1 .LUT_INIT=16'b1010101010000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i13_LC_9_25_1  (
            .in0(N__27453),
            .in1(N__44932),
            .in2(N__44603),
            .in3(N__44768),
            .lcout(\c0.FRAME_MATCHER_state_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49755),
            .ce(),
            .sr(N__27441));
    defparam \c0.i1_2_lut_adj_712_LC_9_25_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_712_LC_9_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_712_LC_9_25_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_712_LC_9_25_2  (
            .in0(_gnd_net_),
            .in1(N__27452),
            .in2(_gnd_net_),
            .in3(N__40796),
            .lcout(\c0.n8_adj_2332 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_723_LC_9_25_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_723_LC_9_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_723_LC_9_25_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i1_2_lut_adj_723_LC_9_25_3  (
            .in0(N__40798),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27432),
            .lcout(\c0.n8_adj_2328 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_705_LC_9_25_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_705_LC_9_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_705_LC_9_25_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_705_LC_9_25_4  (
            .in0(_gnd_net_),
            .in1(N__27396),
            .in2(_gnd_net_),
            .in3(N__40793),
            .lcout(\c0.n8_adj_2334 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_709_LC_9_25_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_709_LC_9_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_709_LC_9_25_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i1_2_lut_adj_709_LC_9_25_5  (
            .in0(N__40794),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37299),
            .lcout(\c0.n8_adj_2333 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_711_LC_9_25_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_711_LC_9_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_711_LC_9_25_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_711_LC_9_25_6  (
            .in0(_gnd_net_),
            .in1(N__27351),
            .in2(_gnd_net_),
            .in3(N__40795),
            .lcout(\c0.n16708 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_713_LC_9_25_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_713_LC_9_25_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_713_LC_9_25_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i1_2_lut_adj_713_LC_9_25_7  (
            .in0(N__40797),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27324),
            .lcout(\c0.n8_adj_2331 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_718_LC_9_26_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_718_LC_9_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_718_LC_9_26_0 .LUT_INIT=16'b1000110010001000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_718_LC_9_26_0  (
            .in0(N__41332),
            .in1(N__27483),
            .in2(N__41427),
            .in3(N__41457),
            .lcout(\c0.n16716 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_594_LC_9_26_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_594_LC_9_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_594_LC_9_26_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_594_LC_9_26_1  (
            .in0(N__27656),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27606),
            .lcout(\c0.n10459 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_adj_398_LC_9_26_3 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_adj_398_LC_9_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_adj_398_LC_9_26_3 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \c0.rx.i1_2_lut_adj_398_LC_9_26_3  (
            .in0(N__37868),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37829),
            .lcout(n10010),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__5__2288_LC_9_26_4 .C_ON=1'b0;
    defparam \c0.data_in_0__5__2288_LC_9_26_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__5__2288_LC_9_26_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0__5__2288_LC_9_26_4  (
            .in0(N__27515),
            .in1(N__39131),
            .in2(_gnd_net_),
            .in3(N__27562),
            .lcout(data_in_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49768),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__4__2289_LC_9_26_5 .C_ON=1'b0;
    defparam \c0.data_in_0__4__2289_LC_9_26_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__4__2289_LC_9_26_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0__4__2289_LC_9_26_5  (
            .in0(N__39129),
            .in1(N__29241),
            .in2(_gnd_net_),
            .in3(N__27545),
            .lcout(data_in_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49768),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__2__2291_LC_9_26_6 .C_ON=1'b0;
    defparam \c0.data_in_0__2__2291_LC_9_26_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__2__2291_LC_9_26_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_0__2__2291_LC_9_26_6  (
            .in0(N__28054),
            .in1(N__39130),
            .in2(_gnd_net_),
            .in3(N__27530),
            .lcout(data_in_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49768),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__5__2280_LC_9_26_7 .C_ON=1'b0;
    defparam \c0.data_in_1__5__2280_LC_9_26_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__5__2280_LC_9_26_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_1__5__2280_LC_9_26_7  (
            .in0(N__29181),
            .in1(N__39132),
            .in2(_gnd_net_),
            .in3(N__27514),
            .lcout(data_in_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49768),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_i_i16_LC_9_27_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_i_i16_LC_9_27_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_i_i16_LC_9_27_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_i_i16_LC_9_27_0  (
            .in0(_gnd_net_),
            .in1(N__27498),
            .in2(_gnd_net_),
            .in3(N__33159),
            .lcout(\c0.FRAME_MATCHER_i_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49780),
            .ce(),
            .sr(N__27687));
    defparam \c0.FRAME_MATCHER_state_i4_LC_9_28_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i4_LC_9_28_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i4_LC_9_28_0 .LUT_INIT=16'b1110110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i4_LC_9_28_0  (
            .in0(N__44986),
            .in1(N__44798),
            .in2(N__44616),
            .in3(N__27481),
            .lcout(\c0.FRAME_MATCHER_state_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49790),
            .ce(),
            .sr(N__27462));
    defparam \c0.i2_3_lut_adj_628_LC_9_28_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_628_LC_9_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_628_LC_9_28_1 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \c0.i2_3_lut_adj_628_LC_9_28_1  (
            .in0(N__28055),
            .in1(N__35092),
            .in2(_gnd_net_),
            .in3(N__35385),
            .lcout(\c0.n10141 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14611_2_lut_LC_9_28_2 .C_ON=1'b0;
    defparam \c0.i14611_2_lut_LC_9_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.i14611_2_lut_LC_9_28_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i14611_2_lut_LC_9_28_2  (
            .in0(N__35093),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28056),
            .lcout(\c0.n17388 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_219_Select_10_i3_2_lut_3_lut_LC_9_28_3 .C_ON=1'b0;
    defparam \c0.select_219_Select_10_i3_2_lut_3_lut_LC_9_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.select_219_Select_10_i3_2_lut_3_lut_LC_9_28_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \c0.select_219_Select_10_i3_2_lut_3_lut_LC_9_28_3  (
            .in0(N__41845),
            .in1(N__27821),
            .in2(_gnd_net_),
            .in3(N__28001),
            .lcout(\c0.n3_adj_2272 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10678_2_lut_LC_9_28_4 .C_ON=1'b0;
    defparam \c0.i10678_2_lut_LC_9_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.i10678_2_lut_LC_9_28_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i10678_2_lut_LC_9_28_4  (
            .in0(_gnd_net_),
            .in1(N__28000),
            .in2(_gnd_net_),
            .in3(N__41844),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_219_Select_14_i3_2_lut_3_lut_LC_9_28_5 .C_ON=1'b0;
    defparam \c0.select_219_Select_14_i3_2_lut_3_lut_LC_9_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.select_219_Select_14_i3_2_lut_3_lut_LC_9_28_5 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \c0.select_219_Select_14_i3_2_lut_3_lut_LC_9_28_5  (
            .in0(N__41846),
            .in1(_gnd_net_),
            .in2(N__27942),
            .in3(N__27820),
            .lcout(\c0.n3_adj_2264 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10674_2_lut_LC_9_28_6 .C_ON=1'b0;
    defparam \c0.i10674_2_lut_LC_9_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.i10674_2_lut_LC_9_28_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i10674_2_lut_LC_9_28_6  (
            .in0(_gnd_net_),
            .in1(N__27937),
            .in2(_gnd_net_),
            .in3(N__41843),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_219_Select_16_i3_2_lut_3_lut_LC_9_28_7 .C_ON=1'b0;
    defparam \c0.select_219_Select_16_i3_2_lut_3_lut_LC_9_28_7 .SEQ_MODE=4'b0000;
    defparam \c0.select_219_Select_16_i3_2_lut_3_lut_LC_9_28_7 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \c0.select_219_Select_16_i3_2_lut_3_lut_LC_9_28_7  (
            .in0(N__41847),
            .in1(N__27873),
            .in2(_gnd_net_),
            .in3(N__27822),
            .lcout(\c0.n3_adj_2259 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2360__i0_LC_9_29_0.C_ON=1'b1;
    defparam blink_counter_2360__i0_LC_9_29_0.SEQ_MODE=4'b1000;
    defparam blink_counter_2360__i0_LC_9_29_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2360__i0_LC_9_29_0 (
            .in0(_gnd_net_),
            .in1(N__27675),
            .in2(_gnd_net_),
            .in3(N__27669),
            .lcout(n26_adj_2423),
            .ltout(),
            .carryin(bfn_9_29_0_),
            .carryout(n16041),
            .clk(N__49800),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2360__i1_LC_9_29_1.C_ON=1'b1;
    defparam blink_counter_2360__i1_LC_9_29_1.SEQ_MODE=4'b1000;
    defparam blink_counter_2360__i1_LC_9_29_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2360__i1_LC_9_29_1 (
            .in0(_gnd_net_),
            .in1(N__27666),
            .in2(_gnd_net_),
            .in3(N__27660),
            .lcout(n25_adj_2424),
            .ltout(),
            .carryin(n16041),
            .carryout(n16042),
            .clk(N__49800),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2360__i2_LC_9_29_2.C_ON=1'b1;
    defparam blink_counter_2360__i2_LC_9_29_2.SEQ_MODE=4'b1000;
    defparam blink_counter_2360__i2_LC_9_29_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2360__i2_LC_9_29_2 (
            .in0(_gnd_net_),
            .in1(N__28137),
            .in2(_gnd_net_),
            .in3(N__28131),
            .lcout(n24),
            .ltout(),
            .carryin(n16042),
            .carryout(n16043),
            .clk(N__49800),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2360__i3_LC_9_29_3.C_ON=1'b1;
    defparam blink_counter_2360__i3_LC_9_29_3.SEQ_MODE=4'b1000;
    defparam blink_counter_2360__i3_LC_9_29_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2360__i3_LC_9_29_3 (
            .in0(_gnd_net_),
            .in1(N__28128),
            .in2(_gnd_net_),
            .in3(N__28122),
            .lcout(n23_adj_2425),
            .ltout(),
            .carryin(n16043),
            .carryout(n16044),
            .clk(N__49800),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2360__i4_LC_9_29_4.C_ON=1'b1;
    defparam blink_counter_2360__i4_LC_9_29_4.SEQ_MODE=4'b1000;
    defparam blink_counter_2360__i4_LC_9_29_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2360__i4_LC_9_29_4 (
            .in0(_gnd_net_),
            .in1(N__28119),
            .in2(_gnd_net_),
            .in3(N__28113),
            .lcout(n22_adj_2426),
            .ltout(),
            .carryin(n16044),
            .carryout(n16045),
            .clk(N__49800),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2360__i5_LC_9_29_5.C_ON=1'b1;
    defparam blink_counter_2360__i5_LC_9_29_5.SEQ_MODE=4'b1000;
    defparam blink_counter_2360__i5_LC_9_29_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2360__i5_LC_9_29_5 (
            .in0(_gnd_net_),
            .in1(N__28110),
            .in2(_gnd_net_),
            .in3(N__28104),
            .lcout(n21),
            .ltout(),
            .carryin(n16045),
            .carryout(n16046),
            .clk(N__49800),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2360__i6_LC_9_29_6.C_ON=1'b1;
    defparam blink_counter_2360__i6_LC_9_29_6.SEQ_MODE=4'b1000;
    defparam blink_counter_2360__i6_LC_9_29_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2360__i6_LC_9_29_6 (
            .in0(_gnd_net_),
            .in1(N__28101),
            .in2(_gnd_net_),
            .in3(N__28095),
            .lcout(n20),
            .ltout(),
            .carryin(n16046),
            .carryout(n16047),
            .clk(N__49800),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2360__i7_LC_9_29_7.C_ON=1'b1;
    defparam blink_counter_2360__i7_LC_9_29_7.SEQ_MODE=4'b1000;
    defparam blink_counter_2360__i7_LC_9_29_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2360__i7_LC_9_29_7 (
            .in0(_gnd_net_),
            .in1(N__28092),
            .in2(_gnd_net_),
            .in3(N__28086),
            .lcout(n19),
            .ltout(),
            .carryin(n16047),
            .carryout(n16048),
            .clk(N__49800),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2360__i8_LC_9_30_0.C_ON=1'b1;
    defparam blink_counter_2360__i8_LC_9_30_0.SEQ_MODE=4'b1000;
    defparam blink_counter_2360__i8_LC_9_30_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2360__i8_LC_9_30_0 (
            .in0(_gnd_net_),
            .in1(N__28083),
            .in2(_gnd_net_),
            .in3(N__28077),
            .lcout(n18),
            .ltout(),
            .carryin(bfn_9_30_0_),
            .carryout(n16049),
            .clk(N__49807),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2360__i9_LC_9_30_1.C_ON=1'b1;
    defparam blink_counter_2360__i9_LC_9_30_1.SEQ_MODE=4'b1000;
    defparam blink_counter_2360__i9_LC_9_30_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2360__i9_LC_9_30_1 (
            .in0(_gnd_net_),
            .in1(N__28074),
            .in2(_gnd_net_),
            .in3(N__28068),
            .lcout(n17),
            .ltout(),
            .carryin(n16049),
            .carryout(n16050),
            .clk(N__49807),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2360__i10_LC_9_30_2.C_ON=1'b1;
    defparam blink_counter_2360__i10_LC_9_30_2.SEQ_MODE=4'b1000;
    defparam blink_counter_2360__i10_LC_9_30_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2360__i10_LC_9_30_2 (
            .in0(_gnd_net_),
            .in1(N__28065),
            .in2(_gnd_net_),
            .in3(N__28059),
            .lcout(n16),
            .ltout(),
            .carryin(n16050),
            .carryout(n16051),
            .clk(N__49807),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2360__i11_LC_9_30_3.C_ON=1'b1;
    defparam blink_counter_2360__i11_LC_9_30_3.SEQ_MODE=4'b1000;
    defparam blink_counter_2360__i11_LC_9_30_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2360__i11_LC_9_30_3 (
            .in0(_gnd_net_),
            .in1(N__28209),
            .in2(_gnd_net_),
            .in3(N__28203),
            .lcout(n15),
            .ltout(),
            .carryin(n16051),
            .carryout(n16052),
            .clk(N__49807),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2360__i12_LC_9_30_4.C_ON=1'b1;
    defparam blink_counter_2360__i12_LC_9_30_4.SEQ_MODE=4'b1000;
    defparam blink_counter_2360__i12_LC_9_30_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2360__i12_LC_9_30_4 (
            .in0(_gnd_net_),
            .in1(N__28200),
            .in2(_gnd_net_),
            .in3(N__28194),
            .lcout(n14),
            .ltout(),
            .carryin(n16052),
            .carryout(n16053),
            .clk(N__49807),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2360__i13_LC_9_30_5.C_ON=1'b1;
    defparam blink_counter_2360__i13_LC_9_30_5.SEQ_MODE=4'b1000;
    defparam blink_counter_2360__i13_LC_9_30_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2360__i13_LC_9_30_5 (
            .in0(_gnd_net_),
            .in1(N__28191),
            .in2(_gnd_net_),
            .in3(N__28185),
            .lcout(n13),
            .ltout(),
            .carryin(n16053),
            .carryout(n16054),
            .clk(N__49807),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2360__i14_LC_9_30_6.C_ON=1'b1;
    defparam blink_counter_2360__i14_LC_9_30_6.SEQ_MODE=4'b1000;
    defparam blink_counter_2360__i14_LC_9_30_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2360__i14_LC_9_30_6 (
            .in0(_gnd_net_),
            .in1(N__28182),
            .in2(_gnd_net_),
            .in3(N__28176),
            .lcout(n12),
            .ltout(),
            .carryin(n16054),
            .carryout(n16055),
            .clk(N__49807),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2360__i15_LC_9_30_7.C_ON=1'b1;
    defparam blink_counter_2360__i15_LC_9_30_7.SEQ_MODE=4'b1000;
    defparam blink_counter_2360__i15_LC_9_30_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2360__i15_LC_9_30_7 (
            .in0(_gnd_net_),
            .in1(N__28173),
            .in2(_gnd_net_),
            .in3(N__28167),
            .lcout(n11),
            .ltout(),
            .carryin(n16055),
            .carryout(n16056),
            .clk(N__49807),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2360__i16_LC_9_31_0.C_ON=1'b1;
    defparam blink_counter_2360__i16_LC_9_31_0.SEQ_MODE=4'b1000;
    defparam blink_counter_2360__i16_LC_9_31_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2360__i16_LC_9_31_0 (
            .in0(_gnd_net_),
            .in1(N__28164),
            .in2(_gnd_net_),
            .in3(N__28158),
            .lcout(n10_adj_2420),
            .ltout(),
            .carryin(bfn_9_31_0_),
            .carryout(n16057),
            .clk(N__49815),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2360__i17_LC_9_31_1.C_ON=1'b1;
    defparam blink_counter_2360__i17_LC_9_31_1.SEQ_MODE=4'b1000;
    defparam blink_counter_2360__i17_LC_9_31_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2360__i17_LC_9_31_1 (
            .in0(_gnd_net_),
            .in1(N__28155),
            .in2(_gnd_net_),
            .in3(N__28149),
            .lcout(n9_adj_2421),
            .ltout(),
            .carryin(n16057),
            .carryout(n16058),
            .clk(N__49815),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2360__i18_LC_9_31_2.C_ON=1'b1;
    defparam blink_counter_2360__i18_LC_9_31_2.SEQ_MODE=4'b1000;
    defparam blink_counter_2360__i18_LC_9_31_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2360__i18_LC_9_31_2 (
            .in0(_gnd_net_),
            .in1(N__28146),
            .in2(_gnd_net_),
            .in3(N__28140),
            .lcout(n8_adj_2412),
            .ltout(),
            .carryin(n16058),
            .carryout(n16059),
            .clk(N__49815),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2360__i19_LC_9_31_3.C_ON=1'b1;
    defparam blink_counter_2360__i19_LC_9_31_3.SEQ_MODE=4'b1000;
    defparam blink_counter_2360__i19_LC_9_31_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2360__i19_LC_9_31_3 (
            .in0(_gnd_net_),
            .in1(N__28248),
            .in2(_gnd_net_),
            .in3(N__28242),
            .lcout(n7),
            .ltout(),
            .carryin(n16059),
            .carryout(n16060),
            .clk(N__49815),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2360__i20_LC_9_31_4.C_ON=1'b1;
    defparam blink_counter_2360__i20_LC_9_31_4.SEQ_MODE=4'b1000;
    defparam blink_counter_2360__i20_LC_9_31_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2360__i20_LC_9_31_4 (
            .in0(_gnd_net_),
            .in1(N__28239),
            .in2(_gnd_net_),
            .in3(N__28233),
            .lcout(n6_adj_2429),
            .ltout(),
            .carryin(n16060),
            .carryout(n16061),
            .clk(N__49815),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2360__i21_LC_9_31_5.C_ON=1'b1;
    defparam blink_counter_2360__i21_LC_9_31_5.SEQ_MODE=4'b1000;
    defparam blink_counter_2360__i21_LC_9_31_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2360__i21_LC_9_31_5 (
            .in0(_gnd_net_),
            .in1(N__36154),
            .in2(_gnd_net_),
            .in3(N__28230),
            .lcout(blink_counter_21),
            .ltout(),
            .carryin(n16061),
            .carryout(n16062),
            .clk(N__49815),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2360__i22_LC_9_31_6.C_ON=1'b1;
    defparam blink_counter_2360__i22_LC_9_31_6.SEQ_MODE=4'b1000;
    defparam blink_counter_2360__i22_LC_9_31_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2360__i22_LC_9_31_6 (
            .in0(_gnd_net_),
            .in1(N__36190),
            .in2(_gnd_net_),
            .in3(N__28227),
            .lcout(blink_counter_22),
            .ltout(),
            .carryin(n16062),
            .carryout(n16063),
            .clk(N__49815),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2360__i23_LC_9_31_7.C_ON=1'b1;
    defparam blink_counter_2360__i23_LC_9_31_7.SEQ_MODE=4'b1000;
    defparam blink_counter_2360__i23_LC_9_31_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2360__i23_LC_9_31_7 (
            .in0(_gnd_net_),
            .in1(N__36226),
            .in2(_gnd_net_),
            .in3(N__28224),
            .lcout(blink_counter_23),
            .ltout(),
            .carryin(n16063),
            .carryout(n16064),
            .clk(N__49815),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2360__i24_LC_9_32_0.C_ON=1'b1;
    defparam blink_counter_2360__i24_LC_9_32_0.SEQ_MODE=4'b1000;
    defparam blink_counter_2360__i24_LC_9_32_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2360__i24_LC_9_32_0 (
            .in0(_gnd_net_),
            .in1(N__36257),
            .in2(_gnd_net_),
            .in3(N__28221),
            .lcout(blink_counter_24),
            .ltout(),
            .carryin(bfn_9_32_0_),
            .carryout(n16065),
            .clk(N__49823),
            .ce(),
            .sr(_gnd_net_));
    defparam blink_counter_2360__i25_LC_9_32_1.C_ON=1'b0;
    defparam blink_counter_2360__i25_LC_9_32_1.SEQ_MODE=4'b1000;
    defparam blink_counter_2360__i25_LC_9_32_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 blink_counter_2360__i25_LC_9_32_1 (
            .in0(_gnd_net_),
            .in1(N__36005),
            .in2(_gnd_net_),
            .in3(N__28218),
            .lcout(blink_counter_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49823),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_i3_LC_10_16_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_i3_LC_10_16_0 .SEQ_MODE=4'b1001;
    defparam \c0.byte_transmit_counter2_i3_LC_10_16_0 .LUT_INIT=16'b1100101000000000;
    LogicCell40 \c0.byte_transmit_counter2_i3_LC_10_16_0  (
            .in0(N__28215),
            .in1(N__32363),
            .in2(N__39678),
            .in3(N__42096),
            .lcout(\c0.byte_transmit_counter2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49679),
            .ce(),
            .sr(N__29079));
    defparam \c0.i10493_2_lut_LC_10_17_0 .C_ON=1'b0;
    defparam \c0.i10493_2_lut_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10493_2_lut_LC_10_17_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i10493_2_lut_LC_10_17_0  (
            .in0(_gnd_net_),
            .in1(N__35606),
            .in2(_gnd_net_),
            .in3(N__34398),
            .lcout(\c0.n11867 ),
            .ltout(\c0.n11867_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_i0_LC_10_17_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_i0_LC_10_17_1 .SEQ_MODE=4'b1001;
    defparam \c0.byte_transmit_counter2_i0_LC_10_17_1 .LUT_INIT=16'b1100101000000000;
    LogicCell40 \c0.byte_transmit_counter2_i0_LC_10_17_1  (
            .in0(N__29097),
            .in1(N__28818),
            .in2(N__29091),
            .in3(N__42093),
            .lcout(\c0.byte_transmit_counter2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49668),
            .ce(),
            .sr(N__29088));
    defparam \c0.i1_2_lut_adj_763_LC_10_17_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_763_LC_10_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_763_LC_10_17_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i1_2_lut_adj_763_LC_10_17_2  (
            .in0(N__28817),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33535),
            .lcout(\c0.n4_adj_2187 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_412_LC_10_17_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_412_LC_10_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_412_LC_10_17_5 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \c0.i1_2_lut_adj_412_LC_10_17_5  (
            .in0(N__33534),
            .in1(N__32362),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.n4_adj_2152 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15170_3_lut_LC_10_17_7 .C_ON=1'b0;
    defparam \c0.i15170_3_lut_LC_10_17_7 .SEQ_MODE=4'b0000;
    defparam \c0.i15170_3_lut_LC_10_17_7 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \c0.i15170_3_lut_LC_10_17_7  (
            .in0(N__37580),
            .in1(N__28360),
            .in2(_gnd_net_),
            .in3(N__28816),
            .lcout(\c0.n17761 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i47_LC_10_18_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i47_LC_10_18_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i47_LC_10_18_0 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \c0.data_in_frame_0__i47_LC_10_18_0  (
            .in0(N__40421),
            .in1(N__32492),
            .in2(N__39554),
            .in3(N__32706),
            .lcout(\c0.data_in_frame_5_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49680),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i31_LC_10_18_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i31_LC_10_18_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i31_LC_10_18_1 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0__i31_LC_10_18_1  (
            .in0(N__28257),
            .in1(N__39545),
            .in2(N__40623),
            .in3(N__39394),
            .lcout(\c0.data_in_frame_3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49680),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_408_LC_10_18_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_408_LC_10_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_408_LC_10_18_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_408_LC_10_18_4  (
            .in0(_gnd_net_),
            .in1(N__28361),
            .in2(_gnd_net_),
            .in3(N__33536),
            .lcout(\c0.n4_adj_2155 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i12_LC_10_18_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i12_LC_10_18_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i12_LC_10_18_5 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i12_LC_10_18_5  (
            .in0(N__40606),
            .in1(N__35276),
            .in2(N__38899),
            .in3(N__40422),
            .lcout(\c0.data_in_frame_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49680),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_562_LC_10_18_7 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_562_LC_10_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_562_LC_10_18_7 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \c0.i5_4_lut_adj_562_LC_10_18_7  (
            .in0(N__28256),
            .in1(N__37010),
            .in2(N__29301),
            .in3(N__34832),
            .lcout(\c0.n19_adj_2303 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i3_LC_10_19_0 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i3_LC_10_19_0 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i3_LC_10_19_0 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.rx.r_Rx_Byte_i3_LC_10_19_0  (
            .in0(N__37983),
            .in1(N__45260),
            .in2(N__35297),
            .in3(N__36710),
            .lcout(rx_data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49689),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i52_LC_10_19_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i52_LC_10_19_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i52_LC_10_19_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0__i52_LC_10_19_2  (
            .in0(N__35287),
            .in1(N__32936),
            .in2(_gnd_net_),
            .in3(N__32564),
            .lcout(data_in_frame_6_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49689),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i32_LC_10_19_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i32_LC_10_19_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i32_LC_10_19_3 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i32_LC_10_19_3  (
            .in0(N__40619),
            .in1(N__40504),
            .in2(N__37523),
            .in3(N__39386),
            .lcout(\c0.data_in_frame_3_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49689),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_574_LC_10_19_4 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_574_LC_10_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_574_LC_10_19_4 .LUT_INIT=16'b1111011001101111;
    LogicCell40 \c0.i1_4_lut_adj_574_LC_10_19_4  (
            .in0(N__29108),
            .in1(N__32765),
            .in2(N__39288),
            .in3(N__32619),
            .lcout(),
            .ltout(\c0.n15_adj_2310_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_595_LC_10_19_5 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_595_LC_10_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_595_LC_10_19_5 .LUT_INIT=16'b1111110111110111;
    LogicCell40 \c0.i8_4_lut_adj_595_LC_10_19_5  (
            .in0(N__34161),
            .in1(N__36906),
            .in2(N__29112),
            .in3(N__37471),
            .lcout(\c0.n22_adj_2319 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__5__2264_LC_10_19_6 .C_ON=1'b0;
    defparam \c0.data_in_3__5__2264_LC_10_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__5__2264_LC_10_19_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_3__5__2264_LC_10_19_6  (
            .in0(N__36675),
            .in1(N__39208),
            .in2(_gnd_net_),
            .in3(N__29646),
            .lcout(data_in_3_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49689),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i28_LC_10_19_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i28_LC_10_19_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i28_LC_10_19_7 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0__i28_LC_10_19_7  (
            .in0(N__29109),
            .in1(N__35288),
            .in2(N__40626),
            .in3(N__39385),
            .lcout(\c0.data_in_frame_3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49689),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i14_LC_10_20_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i14_LC_10_20_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i14_LC_10_20_0 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0__i14_LC_10_20_0  (
            .in0(N__40600),
            .in1(N__34521),
            .in2(N__36689),
            .in3(N__40419),
            .lcout(\c0.data_in_frame_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49699),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i45_LC_10_20_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i45_LC_10_20_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i45_LC_10_20_1 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \c0.data_in_frame_0__i45_LC_10_20_1  (
            .in0(N__40418),
            .in1(N__38849),
            .in2(N__45133),
            .in3(N__32680),
            .lcout(\c0.data_in_frame_5_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49699),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i51_LC_10_20_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i51_LC_10_20_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i51_LC_10_20_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0__i51_LC_10_20_2  (
            .in0(N__36877),
            .in1(N__34343),
            .in2(_gnd_net_),
            .in3(N__32559),
            .lcout(data_in_frame_6_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49699),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_696_LC_10_20_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_696_LC_10_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_696_LC_10_20_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_696_LC_10_20_3  (
            .in0(N__34767),
            .in1(N__37397),
            .in2(_gnd_net_),
            .in3(N__34574),
            .lcout(\c0.n2137 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i42_LC_10_20_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i42_LC_10_20_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i42_LC_10_20_4 .LUT_INIT=16'b1010101011001010;
    LogicCell40 \c0.data_in_frame_0__i42_LC_10_20_4  (
            .in0(N__34655),
            .in1(N__39476),
            .in2(N__32695),
            .in3(N__40420),
            .lcout(\c0.data_in_frame_5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49699),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i54_LC_10_20_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i54_LC_10_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i54_LC_10_20_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_frame_0__i54_LC_10_20_5  (
            .in0(N__32560),
            .in1(N__36680),
            .in2(_gnd_net_),
            .in3(N__34253),
            .lcout(data_in_frame_6_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49699),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_616_LC_10_20_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_616_LC_10_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_616_LC_10_20_6 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \c0.i2_3_lut_adj_616_LC_10_20_6  (
            .in0(N__37113),
            .in1(N__37187),
            .in2(_gnd_net_),
            .in3(N__39362),
            .lcout(n17075),
            .ltout(n17075_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i56_LC_10_20_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i56_LC_10_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i56_LC_10_20_7 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \c0.data_in_frame_0__i56_LC_10_20_7  (
            .in0(N__40505),
            .in1(_gnd_net_),
            .in2(N__29184),
            .in3(N__34974),
            .lcout(data_in_frame_6_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49699),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__7__2270_LC_10_21_0 .C_ON=1'b0;
    defparam \c0.data_in_2__7__2270_LC_10_21_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__7__2270_LC_10_21_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_2__7__2270_LC_10_21_0  (
            .in0(N__39217),
            .in1(N__29392),
            .in2(_gnd_net_),
            .in3(N__32921),
            .lcout(data_in_2_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49712),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14623_3_lut_LC_10_21_1 .C_ON=1'b0;
    defparam \c0.i14623_3_lut_LC_10_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i14623_3_lut_LC_10_21_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.i14623_3_lut_LC_10_21_1  (
            .in0(N__29391),
            .in1(N__29175),
            .in2(_gnd_net_),
            .in3(N__29278),
            .lcout(),
            .ltout(\c0.n17400_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_637_LC_10_21_2 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_637_LC_10_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_637_LC_10_21_2 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \c0.i3_4_lut_adj_637_LC_10_21_2  (
            .in0(N__29149),
            .in1(N__38932),
            .in2(N__29124),
            .in3(N__32898),
            .lcout(),
            .ltout(\c0.n8_adj_2359_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_640_LC_10_21_3 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_640_LC_10_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_640_LC_10_21_3 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \c0.i1_4_lut_adj_640_LC_10_21_3  (
            .in0(N__29647),
            .in1(N__29710),
            .in2(N__29121),
            .in3(N__29118),
            .lcout(\c0.n10136 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__7__2278_LC_10_21_4 .C_ON=1'b0;
    defparam \c0.data_in_1__7__2278_LC_10_21_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__7__2278_LC_10_21_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_1__7__2278_LC_10_21_4  (
            .in0(N__39216),
            .in1(N__29333),
            .in2(_gnd_net_),
            .in3(N__29393),
            .lcout(data_in_1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49712),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i29_LC_10_21_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i29_LC_10_21_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i29_LC_10_21_5 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i29_LC_10_21_5  (
            .in0(N__40599),
            .in1(N__45134),
            .in2(N__29300),
            .in3(N__39361),
            .lcout(\c0.data_in_frame_3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49712),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__7__2262_LC_10_21_6 .C_ON=1'b0;
    defparam \c0.data_in_3__7__2262_LC_10_21_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__7__2262_LC_10_21_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_3__7__2262_LC_10_21_6  (
            .in0(N__40503),
            .in1(N__39215),
            .in2(_gnd_net_),
            .in3(N__32920),
            .lcout(data_in_3_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49712),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__1__2292_LC_10_21_7 .C_ON=1'b0;
    defparam \c0.data_in_0__1__2292_LC_10_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__1__2292_LC_10_21_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_0__1__2292_LC_10_21_7  (
            .in0(N__39214),
            .in1(N__35384),
            .in2(_gnd_net_),
            .in3(N__29279),
            .lcout(data_in_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49712),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i18_3_lut_4_lut_LC_10_22_0 .C_ON=1'b0;
    defparam \c0.i18_3_lut_4_lut_LC_10_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i18_3_lut_4_lut_LC_10_22_0 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \c0.i18_3_lut_4_lut_LC_10_22_0  (
            .in0(N__36091),
            .in1(N__44862),
            .in2(N__41976),
            .in3(N__41700),
            .lcout(),
            .ltout(\c0.n7_adj_2384_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i3_LC_10_22_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i3_LC_10_22_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i3_LC_10_22_1 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i3_LC_10_22_1  (
            .in0(N__33488),
            .in1(N__33669),
            .in2(N__29265),
            .in3(N__35757),
            .lcout(\c0.FRAME_MATCHER_state_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49724),
            .ce(),
            .sr(N__29262));
    defparam \c0.i1_2_lut_adj_700_LC_10_22_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_700_LC_10_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_700_LC_10_22_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_700_LC_10_22_2  (
            .in0(_gnd_net_),
            .in1(N__33487),
            .in2(_gnd_net_),
            .in3(N__41297),
            .lcout(\c0.n6_adj_2336 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_LC_10_22_3 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_LC_10_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_LC_10_22_3 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \c0.i1_3_lut_4_lut_LC_10_22_3  (
            .in0(N__33384),
            .in1(N__41606),
            .in2(N__33740),
            .in3(N__33359),
            .lcout(\c0.n9369 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_645_LC_10_22_4 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_645_LC_10_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_645_LC_10_22_4 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \c0.i6_4_lut_adj_645_LC_10_22_4  (
            .in0(N__29252),
            .in1(N__38978),
            .in2(N__29240),
            .in3(N__34935),
            .lcout(),
            .ltout(\c0.n16_adj_2361_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_647_LC_10_22_5 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_647_LC_10_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_647_LC_10_22_5 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \c0.i9_4_lut_adj_647_LC_10_22_5  (
            .in0(N__29212),
            .in1(N__29375),
            .in2(N__29193),
            .in3(N__29190),
            .lcout(n63),
            .ltout(n63_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_793_LC_10_22_6.C_ON=1'b0;
    defparam i1_4_lut_adj_793_LC_10_22_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_793_LC_10_22_6.LUT_INIT=16'b1011000000110000;
    LogicCell40 i1_4_lut_adj_793_LC_10_22_6 (
            .in0(N__36090),
            .in1(N__33383),
            .in2(N__29400),
            .in3(N__33732),
            .lcout(FRAME_MATCHER_state_31_N_1406_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_649_LC_10_23_0 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_649_LC_10_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_649_LC_10_23_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i6_4_lut_adj_649_LC_10_23_0  (
            .in0(N__38939),
            .in1(N__29397),
            .in2(N__29376),
            .in3(N__29355),
            .lcout(),
            .ltout(\c0.n16_adj_2366_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_670_LC_10_23_1 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_670_LC_10_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_670_LC_10_23_1 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \c0.i9_4_lut_adj_670_LC_10_23_1  (
            .in0(N__29622),
            .in1(N__29349),
            .in2(N__29337),
            .in3(N__29334),
            .lcout(n63_adj_2428),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i16_4_lut_LC_10_23_2 .C_ON=1'b0;
    defparam \c0.i16_4_lut_LC_10_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i16_4_lut_LC_10_23_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i16_4_lut_LC_10_23_2  (
            .in0(N__41268),
            .in1(N__33280),
            .in2(N__41235),
            .in3(N__37335),
            .lcout(\c0.n45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_638_LC_10_23_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_638_LC_10_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_638_LC_10_23_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_638_LC_10_23_3  (
            .in0(N__33354),
            .in1(N__33728),
            .in2(_gnd_net_),
            .in3(N__33380),
            .lcout(n9378),
            .ltout(n9378_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_618_LC_10_23_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_618_LC_10_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_618_LC_10_23_4 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_618_LC_10_23_4  (
            .in0(_gnd_net_),
            .in1(N__33554),
            .in2(N__29310),
            .in3(N__33012),
            .lcout(\c0.n47_adj_2347 ),
            .ltout(\c0.n47_adj_2347_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_762_LC_10_23_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_762_LC_10_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_762_LC_10_23_5 .LUT_INIT=16'b1111010011110000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_762_LC_10_23_5  (
            .in0(N__35941),
            .in1(N__35892),
            .in2(N__29307),
            .in3(N__41669),
            .lcout(\c0.n17069 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_673_LC_10_23_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_673_LC_10_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_673_LC_10_23_6 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \c0.i2_3_lut_adj_673_LC_10_23_6  (
            .in0(N__33381),
            .in1(_gnd_net_),
            .in2(N__33739),
            .in3(N__33355),
            .lcout(\c0.n13146 ),
            .ltout(\c0.n13146_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_LC_10_23_7 .C_ON=1'b0;
    defparam \c0.i1_3_lut_LC_10_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_LC_10_23_7 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \c0.i1_3_lut_LC_10_23_7  (
            .in0(N__35940),
            .in1(_gnd_net_),
            .in2(N__29304),
            .in3(N__35891),
            .lcout(\c0.n4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__4__2265_LC_10_24_0 .C_ON=1'b0;
    defparam \c0.data_in_3__4__2265_LC_10_24_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__4__2265_LC_10_24_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_3__4__2265_LC_10_24_0  (
            .in0(N__45120),
            .in1(N__39190),
            .in2(_gnd_net_),
            .in3(N__29732),
            .lcout(data_in_3_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49745),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14625_4_lut_LC_10_24_1 .C_ON=1'b0;
    defparam \c0.i14625_4_lut_LC_10_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.i14625_4_lut_LC_10_24_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.i14625_4_lut_LC_10_24_1  (
            .in0(N__29711),
            .in1(N__35034),
            .in2(N__29655),
            .in3(N__32922),
            .lcout(\c0.n17402 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_725_LC_10_24_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_725_LC_10_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_725_LC_10_24_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_725_LC_10_24_2  (
            .in0(_gnd_net_),
            .in1(N__29616),
            .in2(_gnd_net_),
            .in3(N__40792),
            .lcout(\c0.n8_adj_2327 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10589_4_lut_LC_10_24_4 .C_ON=1'b0;
    defparam \c0.i10589_4_lut_LC_10_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.i10589_4_lut_LC_10_24_4 .LUT_INIT=16'b0000111100001000;
    LogicCell40 \c0.i10589_4_lut_LC_10_24_4  (
            .in0(N__32880),
            .in1(N__37174),
            .in2(N__29571),
            .in3(N__29508),
            .lcout(n2061),
            .ltout(n2061_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_LC_10_24_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_LC_10_24_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_LC_10_24_5 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \c0.i1_2_lut_LC_10_24_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29496),
            .in3(N__41668),
            .lcout(\c0.n9334 ),
            .ltout(\c0.n9334_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_adj_739_LC_10_24_6 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_adj_739_LC_10_24_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_adj_739_LC_10_24_6 .LUT_INIT=16'b1111111111011100;
    LogicCell40 \c0.i1_3_lut_4_lut_adj_739_LC_10_24_6  (
            .in0(N__41362),
            .in1(N__29493),
            .in2(N__29487),
            .in3(N__29484),
            .lcout(\c0.n15821 ),
            .ltout(\c0.n15821_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_704_LC_10_24_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_704_LC_10_24_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_704_LC_10_24_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \c0.i1_2_lut_adj_704_LC_10_24_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29478),
            .in3(N__33471),
            .lcout(\c0.n8_adj_2335 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2359__i0_LC_10_25_0.C_ON=1'b1;
    defparam rand_setpoint_2359__i0_LC_10_25_0.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2359__i0_LC_10_25_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2359__i0_LC_10_25_0 (
            .in0(_gnd_net_),
            .in1(N__29460),
            .in2(N__38018),
            .in3(_gnd_net_),
            .lcout(rand_setpoint_0),
            .ltout(),
            .carryin(bfn_10_25_0_),
            .carryout(n16010),
            .clk(N__49756),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2359__i1_LC_10_25_1.C_ON=1'b1;
    defparam rand_setpoint_2359__i1_LC_10_25_1.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2359__i1_LC_10_25_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2359__i1_LC_10_25_1 (
            .in0(_gnd_net_),
            .in1(N__30279),
            .in2(N__36410),
            .in3(N__30219),
            .lcout(rand_setpoint_1),
            .ltout(),
            .carryin(n16010),
            .carryout(n16011),
            .clk(N__49756),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2359__i2_LC_10_25_2.C_ON=1'b1;
    defparam rand_setpoint_2359__i2_LC_10_25_2.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2359__i2_LC_10_25_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2359__i2_LC_10_25_2 (
            .in0(_gnd_net_),
            .in1(N__30216),
            .in2(N__33831),
            .in3(N__30174),
            .lcout(rand_setpoint_2),
            .ltout(),
            .carryin(n16011),
            .carryout(n16012),
            .clk(N__49756),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2359__i3_LC_10_25_3.C_ON=1'b1;
    defparam rand_setpoint_2359__i3_LC_10_25_3.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2359__i3_LC_10_25_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2359__i3_LC_10_25_3 (
            .in0(_gnd_net_),
            .in1(N__30162),
            .in2(N__33815),
            .in3(N__30114),
            .lcout(rand_setpoint_3),
            .ltout(),
            .carryin(n16012),
            .carryout(n16013),
            .clk(N__49756),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2359__i4_LC_10_25_4.C_ON=1'b1;
    defparam rand_setpoint_2359__i4_LC_10_25_4.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2359__i4_LC_10_25_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2359__i4_LC_10_25_4 (
            .in0(_gnd_net_),
            .in1(N__30111),
            .in2(N__36338),
            .in3(N__30057),
            .lcout(rand_setpoint_4),
            .ltout(),
            .carryin(n16013),
            .carryout(n16014),
            .clk(N__49756),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2359__i5_LC_10_25_5.C_ON=1'b1;
    defparam rand_setpoint_2359__i5_LC_10_25_5.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2359__i5_LC_10_25_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2359__i5_LC_10_25_5 (
            .in0(_gnd_net_),
            .in1(N__30053),
            .in2(N__43736),
            .in3(N__29997),
            .lcout(rand_setpoint_5),
            .ltout(),
            .carryin(n16014),
            .carryout(n16015),
            .clk(N__49756),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2359__i6_LC_10_25_6.C_ON=1'b1;
    defparam rand_setpoint_2359__i6_LC_10_25_6.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2359__i6_LC_10_25_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2359__i6_LC_10_25_6 (
            .in0(_gnd_net_),
            .in1(N__29994),
            .in2(N__36314),
            .in3(N__29934),
            .lcout(rand_setpoint_6),
            .ltout(),
            .carryin(n16015),
            .carryout(n16016),
            .clk(N__49756),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2359__i7_LC_10_25_7.C_ON=1'b1;
    defparam rand_setpoint_2359__i7_LC_10_25_7.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2359__i7_LC_10_25_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2359__i7_LC_10_25_7 (
            .in0(_gnd_net_),
            .in1(N__29930),
            .in2(N__38153),
            .in3(N__29877),
            .lcout(rand_setpoint_7),
            .ltout(),
            .carryin(n16016),
            .carryout(n16017),
            .clk(N__49756),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2359__i8_LC_10_26_0.C_ON=1'b1;
    defparam rand_setpoint_2359__i8_LC_10_26_0.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2359__i8_LC_10_26_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2359__i8_LC_10_26_0 (
            .in0(_gnd_net_),
            .in1(N__29873),
            .in2(N__42167),
            .in3(N__29820),
            .lcout(rand_setpoint_8),
            .ltout(),
            .carryin(bfn_10_26_0_),
            .carryout(n16018),
            .clk(N__49769),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2359__i9_LC_10_26_1.C_ON=1'b1;
    defparam rand_setpoint_2359__i9_LC_10_26_1.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2359__i9_LC_10_26_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2359__i9_LC_10_26_1 (
            .in0(_gnd_net_),
            .in1(N__29816),
            .in2(N__29753),
            .in3(N__29736),
            .lcout(rand_setpoint_9),
            .ltout(),
            .carryin(n16018),
            .carryout(n16019),
            .clk(N__49769),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2359__i10_LC_10_26_2.C_ON=1'b1;
    defparam rand_setpoint_2359__i10_LC_10_26_2.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2359__i10_LC_10_26_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2359__i10_LC_10_26_2 (
            .in0(_gnd_net_),
            .in1(N__30779),
            .in2(N__31973),
            .in3(N__30720),
            .lcout(rand_setpoint_10),
            .ltout(),
            .carryin(n16019),
            .carryout(n16020),
            .clk(N__49769),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2359__i11_LC_10_26_3.C_ON=1'b1;
    defparam rand_setpoint_2359__i11_LC_10_26_3.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2359__i11_LC_10_26_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2359__i11_LC_10_26_3 (
            .in0(_gnd_net_),
            .in1(N__30707),
            .in2(N__32012),
            .in3(N__30660),
            .lcout(rand_setpoint_11),
            .ltout(),
            .carryin(n16020),
            .carryout(n16021),
            .clk(N__49769),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2359__i12_LC_10_26_4.C_ON=1'b1;
    defparam rand_setpoint_2359__i12_LC_10_26_4.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2359__i12_LC_10_26_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2359__i12_LC_10_26_4 (
            .in0(_gnd_net_),
            .in1(N__30655),
            .in2(N__33983),
            .in3(N__30603),
            .lcout(rand_setpoint_12),
            .ltout(),
            .carryin(n16021),
            .carryout(n16022),
            .clk(N__49769),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2359__i13_LC_10_26_5.C_ON=1'b1;
    defparam rand_setpoint_2359__i13_LC_10_26_5.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2359__i13_LC_10_26_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2359__i13_LC_10_26_5 (
            .in0(_gnd_net_),
            .in1(N__30600),
            .in2(N__43646),
            .in3(N__30540),
            .lcout(rand_setpoint_13),
            .ltout(),
            .carryin(n16022),
            .carryout(n16023),
            .clk(N__49769),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2359__i14_LC_10_26_6.C_ON=1'b1;
    defparam rand_setpoint_2359__i14_LC_10_26_6.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2359__i14_LC_10_26_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2359__i14_LC_10_26_6 (
            .in0(_gnd_net_),
            .in1(N__30535),
            .in2(N__34067),
            .in3(N__30471),
            .lcout(rand_setpoint_14),
            .ltout(),
            .carryin(n16023),
            .carryout(n16024),
            .clk(N__49769),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2359__i15_LC_10_26_7.C_ON=1'b1;
    defparam rand_setpoint_2359__i15_LC_10_26_7.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2359__i15_LC_10_26_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2359__i15_LC_10_26_7 (
            .in0(_gnd_net_),
            .in1(N__30468),
            .in2(N__38099),
            .in3(N__30417),
            .lcout(rand_setpoint_15),
            .ltout(),
            .carryin(n16024),
            .carryout(n16025),
            .clk(N__49769),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2359__i16_LC_10_27_0.C_ON=1'b1;
    defparam rand_setpoint_2359__i16_LC_10_27_0.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2359__i16_LC_10_27_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2359__i16_LC_10_27_0 (
            .in0(_gnd_net_),
            .in1(N__30414),
            .in2(N__38120),
            .in3(N__30366),
            .lcout(rand_setpoint_16),
            .ltout(),
            .carryin(bfn_10_27_0_),
            .carryout(n16026),
            .clk(N__49781),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2359__i17_LC_10_27_1.C_ON=1'b1;
    defparam rand_setpoint_2359__i17_LC_10_27_1.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2359__i17_LC_10_27_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2359__i17_LC_10_27_1 (
            .in0(_gnd_net_),
            .in1(N__30355),
            .in2(N__30299),
            .in3(N__30282),
            .lcout(rand_setpoint_17),
            .ltout(),
            .carryin(n16026),
            .carryout(n16027),
            .clk(N__49781),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2359__i18_LC_10_27_2.C_ON=1'b1;
    defparam rand_setpoint_2359__i18_LC_10_27_2.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2359__i18_LC_10_27_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2359__i18_LC_10_27_2 (
            .in0(_gnd_net_),
            .in1(N__31268),
            .in2(N__33882),
            .in3(N__31212),
            .lcout(rand_setpoint_18),
            .ltout(),
            .carryin(n16027),
            .carryout(n16028),
            .clk(N__49781),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2359__i19_LC_10_27_3.C_ON=1'b1;
    defparam rand_setpoint_2359__i19_LC_10_27_3.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2359__i19_LC_10_27_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2359__i19_LC_10_27_3 (
            .in0(_gnd_net_),
            .in1(N__31201),
            .in2(N__33900),
            .in3(N__31158),
            .lcout(rand_setpoint_19),
            .ltout(),
            .carryin(n16028),
            .carryout(n16029),
            .clk(N__49781),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2359__i20_LC_10_27_4.C_ON=1'b1;
    defparam rand_setpoint_2359__i20_LC_10_27_4.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2359__i20_LC_10_27_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2359__i20_LC_10_27_4 (
            .in0(_gnd_net_),
            .in1(N__31154),
            .in2(N__33945),
            .in3(N__31098),
            .lcout(rand_setpoint_20),
            .ltout(),
            .carryin(n16029),
            .carryout(n16030),
            .clk(N__49781),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2359__i21_LC_10_27_5.C_ON=1'b1;
    defparam rand_setpoint_2359__i21_LC_10_27_5.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2359__i21_LC_10_27_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2359__i21_LC_10_27_5 (
            .in0(_gnd_net_),
            .in1(N__31094),
            .in2(N__33864),
            .in3(N__31035),
            .lcout(rand_setpoint_21),
            .ltout(),
            .carryin(n16030),
            .carryout(n16031),
            .clk(N__49781),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2359__i22_LC_10_27_6.C_ON=1'b1;
    defparam rand_setpoint_2359__i22_LC_10_27_6.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2359__i22_LC_10_27_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2359__i22_LC_10_27_6 (
            .in0(_gnd_net_),
            .in1(N__31031),
            .in2(N__33930),
            .in3(N__30978),
            .lcout(rand_setpoint_22),
            .ltout(),
            .carryin(n16031),
            .carryout(n16032),
            .clk(N__49781),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2359__i23_LC_10_27_7.C_ON=1'b1;
    defparam rand_setpoint_2359__i23_LC_10_27_7.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2359__i23_LC_10_27_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2359__i23_LC_10_27_7 (
            .in0(_gnd_net_),
            .in1(N__30974),
            .in2(N__33764),
            .in3(N__30924),
            .lcout(rand_setpoint_23),
            .ltout(),
            .carryin(n16032),
            .carryout(n16033),
            .clk(N__49781),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2359__i24_LC_10_28_0.C_ON=1'b1;
    defparam rand_setpoint_2359__i24_LC_10_28_0.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2359__i24_LC_10_28_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2359__i24_LC_10_28_0 (
            .in0(_gnd_net_),
            .in1(N__30920),
            .in2(N__30863),
            .in3(N__30846),
            .lcout(rand_setpoint_24),
            .ltout(),
            .carryin(bfn_10_28_0_),
            .carryout(n16034),
            .clk(N__49791),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2359__i25_LC_10_28_1.C_ON=1'b1;
    defparam rand_setpoint_2359__i25_LC_10_28_1.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2359__i25_LC_10_28_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2359__i25_LC_10_28_1 (
            .in0(_gnd_net_),
            .in1(N__30838),
            .in2(N__47894),
            .in3(N__30786),
            .lcout(rand_setpoint_25),
            .ltout(),
            .carryin(n16034),
            .carryout(n16035),
            .clk(N__49791),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2359__i26_LC_10_28_2.C_ON=1'b1;
    defparam rand_setpoint_2359__i26_LC_10_28_2.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2359__i26_LC_10_28_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2359__i26_LC_10_28_2 (
            .in0(_gnd_net_),
            .in1(N__31677),
            .in2(N__31319),
            .in3(N__31626),
            .lcout(rand_setpoint_26),
            .ltout(),
            .carryin(n16035),
            .carryout(n16036),
            .clk(N__49791),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2359__i27_LC_10_28_3.C_ON=1'b1;
    defparam rand_setpoint_2359__i27_LC_10_28_3.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2359__i27_LC_10_28_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2359__i27_LC_10_28_3 (
            .in0(_gnd_net_),
            .in1(N__31614),
            .in2(N__31287),
            .in3(N__31569),
            .lcout(rand_setpoint_27),
            .ltout(),
            .carryin(n16036),
            .carryout(n16037),
            .clk(N__49791),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2359__i28_LC_10_28_4.C_ON=1'b1;
    defparam rand_setpoint_2359__i28_LC_10_28_4.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2359__i28_LC_10_28_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2359__i28_LC_10_28_4 (
            .in0(_gnd_net_),
            .in1(N__31566),
            .in2(N__32031),
            .in3(N__31518),
            .lcout(rand_setpoint_28),
            .ltout(),
            .carryin(n16037),
            .carryout(n16038),
            .clk(N__49791),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2359__i29_LC_10_28_5.C_ON=1'b1;
    defparam rand_setpoint_2359__i29_LC_10_28_5.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2359__i29_LC_10_28_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2359__i29_LC_10_28_5 (
            .in0(_gnd_net_),
            .in1(N__31513),
            .in2(N__31302),
            .in3(N__31461),
            .lcout(rand_setpoint_29),
            .ltout(),
            .carryin(n16038),
            .carryout(n16039),
            .clk(N__49791),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2359__i30_LC_10_28_6.C_ON=1'b1;
    defparam rand_setpoint_2359__i30_LC_10_28_6.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2359__i30_LC_10_28_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 rand_setpoint_2359__i30_LC_10_28_6 (
            .in0(_gnd_net_),
            .in1(N__31454),
            .in2(N__42293),
            .in3(N__31404),
            .lcout(rand_setpoint_30),
            .ltout(),
            .carryin(n16039),
            .carryout(n16040),
            .clk(N__49791),
            .ce(),
            .sr(_gnd_net_));
    defparam rand_setpoint_2359__i31_LC_10_28_7.C_ON=1'b0;
    defparam rand_setpoint_2359__i31_LC_10_28_7.SEQ_MODE=4'b1000;
    defparam rand_setpoint_2359__i31_LC_10_28_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 rand_setpoint_2359__i31_LC_10_28_7 (
            .in0(N__31401),
            .in1(N__31334),
            .in2(_gnd_net_),
            .in3(N__31347),
            .lcout(rand_setpoint_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49791),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_5__2__2214_LC_10_29_0 .C_ON=1'b0;
    defparam \c0.data_out_5__2__2214_LC_10_29_0 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_5__2__2214_LC_10_29_0 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \c0.data_out_5__2__2214_LC_10_29_0  (
            .in0(N__48153),
            .in1(N__31320),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.data_out_5_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49801),
            .ce(N__50575),
            .sr(N__42806));
    defparam \c0.data_out_5__5__2211_LC_10_29_1 .C_ON=1'b0;
    defparam \c0.data_out_5__5__2211_LC_10_29_1 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_5__5__2211_LC_10_29_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.data_out_5__5__2211_LC_10_29_1  (
            .in0(_gnd_net_),
            .in1(N__48152),
            .in2(_gnd_net_),
            .in3(N__31301),
            .lcout(\c0.data_out_5_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49801),
            .ce(N__50575),
            .sr(N__42806));
    defparam \c0.data_out_5__3__2213_LC_10_29_3 .C_ON=1'b0;
    defparam \c0.data_out_5__3__2213_LC_10_29_3 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_5__3__2213_LC_10_29_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.data_out_5__3__2213_LC_10_29_3  (
            .in0(_gnd_net_),
            .in1(N__48151),
            .in2(_gnd_net_),
            .in3(N__31286),
            .lcout(\c0.data_out_5_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49801),
            .ce(N__50575),
            .sr(N__42806));
    defparam \c0.data_out_5__4__2212_LC_10_29_4 .C_ON=1'b0;
    defparam \c0.data_out_5__4__2212_LC_10_29_4 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_5__4__2212_LC_10_29_4 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \c0.data_out_5__4__2212_LC_10_29_4  (
            .in0(N__48154),
            .in1(N__32030),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.data_out_5_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49801),
            .ce(N__50575),
            .sr(N__42806));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_3_i5_3_lut_LC_10_30_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_3_i5_3_lut_LC_10_30_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_3_i5_3_lut_LC_10_30_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_3_i5_3_lut_LC_10_30_1  (
            .in0(N__47156),
            .in1(N__46695),
            .in2(_gnd_net_),
            .in3(N__47819),
            .lcout(\c0.n5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14998_2_lut_LC_10_30_2 .C_ON=1'b0;
    defparam \c0.i14998_2_lut_LC_10_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.i14998_2_lut_LC_10_30_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i14998_2_lut_LC_10_30_2  (
            .in0(_gnd_net_),
            .in1(N__32016),
            .in2(_gnd_net_),
            .in3(N__48130),
            .lcout(\c0.n17585 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14993_2_lut_LC_10_30_5 .C_ON=1'b0;
    defparam \c0.i14993_2_lut_LC_10_30_5 .SEQ_MODE=4'b0000;
    defparam \c0.i14993_2_lut_LC_10_30_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i14993_2_lut_LC_10_30_5  (
            .in0(N__48132),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31977),
            .lcout(),
            .ltout(\c0.n17583_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__2__2198_LC_10_30_6 .C_ON=1'b0;
    defparam \c0.data_out_7__2__2198_LC_10_30_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__2__2198_LC_10_30_6 .LUT_INIT=16'b1010000011100100;
    LogicCell40 \c0.data_out_7__2__2198_LC_10_30_6  (
            .in0(N__50261),
            .in1(N__48409),
            .in2(N__31956),
            .in3(N__47321),
            .lcout(\c0.data_out_7_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49808),
            .ce(N__46923),
            .sr(_gnd_net_));
    defparam \c0.i15230_2_lut_3_lut_LC_10_30_7 .C_ON=1'b0;
    defparam \c0.i15230_2_lut_3_lut_LC_10_30_7 .SEQ_MODE=4'b0000;
    defparam \c0.i15230_2_lut_3_lut_LC_10_30_7 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \c0.i15230_2_lut_3_lut_LC_10_30_7  (
            .in0(N__48131),
            .in1(N__48405),
            .in2(_gnd_net_),
            .in3(N__50260),
            .lcout(\c0.n10594 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_SM_Main_i2_LC_10_31_0 .C_ON=1'b0;
    defparam \c0.rx.r_SM_Main_i2_LC_10_31_0 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_SM_Main_i2_LC_10_31_0 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \c0.rx.r_SM_Main_i2_LC_10_31_0  (
            .in0(N__31737),
            .in1(N__31953),
            .in2(N__31785),
            .in3(N__31899),
            .lcout(r_SM_Main_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49816),
            .ce(),
            .sr(N__31800));
    defparam \c0.rx.i1_2_lut_LC_10_31_1 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_LC_10_31_1 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_LC_10_31_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.rx.i1_2_lut_LC_10_31_1  (
            .in0(_gnd_net_),
            .in1(N__31781),
            .in2(_gnd_net_),
            .in3(N__31736),
            .lcout(\c0.rx.n17080 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_2_i2_3_lut_LC_10_31_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_2_i2_3_lut_LC_10_31_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_2_i2_3_lut_LC_10_31_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_2_i2_3_lut_LC_10_31_2  (
            .in0(N__47818),
            .in1(N__34172),
            .in2(_gnd_net_),
            .in3(N__34214),
            .lcout(\c0.n2_adj_2145 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15122_2_lut_LC_10_31_7 .C_ON=1'b0;
    defparam \c0.i15122_2_lut_LC_10_31_7 .SEQ_MODE=4'b0000;
    defparam \c0.i15122_2_lut_LC_10_31_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i15122_2_lut_LC_10_31_7  (
            .in0(_gnd_net_),
            .in1(N__34226),
            .in2(_gnd_net_),
            .in3(N__47817),
            .lcout(\c0.n17622 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10610_3_lut_LC_11_16_0 .C_ON=1'b0;
    defparam \c0.i10610_3_lut_LC_11_16_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10610_3_lut_LC_11_16_0 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \c0.i10610_3_lut_LC_11_16_0  (
            .in0(N__32333),
            .in1(N__32235),
            .in2(_gnd_net_),
            .in3(N__32069),
            .lcout(\c0.n13284 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_i2_LC_11_16_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_i2_LC_11_16_3 .SEQ_MODE=4'b1001;
    defparam \c0.byte_transmit_counter2_i2_LC_11_16_3 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \c0.byte_transmit_counter2_i2_LC_11_16_3  (
            .in0(N__32071),
            .in1(N__32187),
            .in2(N__39693),
            .in3(N__42085),
            .lcout(\c0.byte_transmit_counter2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49690),
            .ce(),
            .sr(N__32049));
    defparam \c0.i1_2_lut_adj_411_LC_11_16_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_411_LC_11_16_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_411_LC_11_16_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_411_LC_11_16_4  (
            .in0(_gnd_net_),
            .in1(N__32070),
            .in2(_gnd_net_),
            .in3(N__33519),
            .lcout(\c0.n4_adj_2154 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_605_LC_11_16_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_605_LC_11_16_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_605_LC_11_16_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i1_2_lut_adj_605_LC_11_16_5  (
            .in0(N__33521),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34441),
            .lcout(\c0.n4_adj_2325 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_679_LC_11_16_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_679_LC_11_16_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_679_LC_11_16_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_679_LC_11_16_6  (
            .in0(_gnd_net_),
            .in1(N__34476),
            .in2(_gnd_net_),
            .in3(N__33522),
            .lcout(\c0.n4_adj_2345 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_465_LC_11_16_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_465_LC_11_16_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_465_LC_11_16_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i1_2_lut_adj_465_LC_11_16_7  (
            .in0(N__33520),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39624),
            .lcout(\c0.n4_adj_2147 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_585_LC_11_17_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_585_LC_11_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_585_LC_11_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_585_LC_11_17_0  (
            .in0(N__32474),
            .in1(N__38822),
            .in2(_gnd_net_),
            .in3(N__39994),
            .lcout(\c0.n16475 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i48_LC_11_17_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i48_LC_11_17_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i48_LC_11_17_1 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \c0.data_in_frame_0__i48_LC_11_17_1  (
            .in0(N__32708),
            .in1(N__34628),
            .in2(N__40509),
            .in3(N__40429),
            .lcout(\c0.data_in_frame_5_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49678),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i46_LC_11_17_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i46_LC_11_17_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i46_LC_11_17_3 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \c0.data_in_frame_0__i46_LC_11_17_3  (
            .in0(N__32707),
            .in1(N__32601),
            .in2(N__36690),
            .in3(N__40428),
            .lcout(\c0.data_in_frame_5_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49678),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1010_2_lut_LC_11_17_4 .C_ON=1'b0;
    defparam \c0.i1010_2_lut_LC_11_17_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1010_2_lut_LC_11_17_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1010_2_lut_LC_11_17_4  (
            .in0(_gnd_net_),
            .in1(N__32751),
            .in2(_gnd_net_),
            .in3(N__34896),
            .lcout(\c0.n2122 ),
            .ltout(\c0.n2122_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_464_LC_11_17_5 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_464_LC_11_17_5 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_464_LC_11_17_5 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \c0.i4_4_lut_adj_464_LC_11_17_5  (
            .in0(N__32506),
            .in1(N__35324),
            .in2(N__32517),
            .in3(N__32766),
            .lcout(\c0.n20_adj_2195 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i22_LC_11_17_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i22_LC_11_17_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i22_LC_11_17_6 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0__i22_LC_11_17_6  (
            .in0(N__37736),
            .in1(N__36687),
            .in2(N__39396),
            .in3(N__32507),
            .lcout(\c0.data_in_frame_2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49678),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i11_LC_11_17_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i11_LC_11_17_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i11_LC_11_17_7 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0__i11_LC_11_17_7  (
            .in0(N__38823),
            .in1(N__36863),
            .in2(N__40625),
            .in3(N__40427),
            .lcout(\c0.data_in_frame_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49678),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i43_LC_11_18_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i43_LC_11_18_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i43_LC_11_18_0 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \c0.data_in_frame_0__i43_LC_11_18_0  (
            .in0(N__32702),
            .in1(N__40050),
            .in2(N__36882),
            .in3(N__40424),
            .lcout(\c0.data_in_frame_5_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49691),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_611_LC_11_18_1 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_611_LC_11_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_611_LC_11_18_1 .LUT_INIT=16'b1001011011111111;
    LogicCell40 \c0.i8_4_lut_adj_611_LC_11_18_1  (
            .in0(N__34528),
            .in1(N__34609),
            .in2(N__32493),
            .in3(N__34491),
            .lcout(\c0.n24_adj_2340 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1012_2_lut_LC_11_18_2 .C_ON=1'b0;
    defparam \c0.i1012_2_lut_LC_11_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1012_2_lut_LC_11_18_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1012_2_lut_LC_11_18_2  (
            .in0(_gnd_net_),
            .in1(N__32749),
            .in2(_gnd_net_),
            .in3(N__34799),
            .lcout(\c0.n2124 ),
            .ltout(\c0.n2124_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_498_LC_11_18_3 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_498_LC_11_18_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_498_LC_11_18_3 .LUT_INIT=16'b0111101111011110;
    LogicCell40 \c0.i1_4_lut_adj_498_LC_11_18_3  (
            .in0(N__34160),
            .in1(N__35120),
            .in2(N__32478),
            .in3(N__37472),
            .lcout(\c0.n17_adj_2214 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i44_LC_11_18_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i44_LC_11_18_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i44_LC_11_18_4 .LUT_INIT=16'b1010101011001010;
    LogicCell40 \c0.data_in_frame_0__i44_LC_11_18_4  (
            .in0(N__32475),
            .in1(N__35277),
            .in2(N__32709),
            .in3(N__40425),
            .lcout(\c0.data_in_frame_5_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49691),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_654_LC_11_18_6 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_654_LC_11_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_654_LC_11_18_6 .LUT_INIT=16'b1111111110111110;
    LogicCell40 \c0.i10_4_lut_adj_654_LC_11_18_6  (
            .in0(N__32607),
            .in1(N__34833),
            .in2(N__32532),
            .in3(N__34944),
            .lcout(\c0.n26_adj_2368 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_634_LC_11_18_7 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_634_LC_11_18_7 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_634_LC_11_18_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_634_LC_11_18_7  (
            .in0(N__32600),
            .in1(N__38885),
            .in2(_gnd_net_),
            .in3(N__34608),
            .lcout(\c0.n16474 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_589_LC_11_19_0 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_589_LC_11_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_589_LC_11_19_0 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \c0.i10_4_lut_adj_589_LC_11_19_0  (
            .in0(N__35325),
            .in1(N__33416),
            .in2(N__32589),
            .in3(N__32574),
            .lcout(\c0.n24_adj_2317 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i4_LC_11_19_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i4_LC_11_19_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i4_LC_11_19_1 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i4_LC_11_19_1  (
            .in0(N__37690),
            .in1(N__40408),
            .in2(N__35292),
            .in3(N__34895),
            .lcout(\c0.data_in_frame_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49700),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i6_LC_11_19_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i6_LC_11_19_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i6_LC_11_19_2 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i6_LC_11_19_2  (
            .in0(N__40406),
            .in1(N__37692),
            .in2(N__36688),
            .in3(N__34800),
            .lcout(\c0.data_in_frame_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49700),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i13_LC_11_19_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i13_LC_11_19_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i13_LC_11_19_3 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i13_LC_11_19_3  (
            .in0(N__40578),
            .in1(N__45131),
            .in2(N__34614),
            .in3(N__40409),
            .lcout(\c0.data_in_frame_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49700),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_adj_730_LC_11_19_4 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_adj_730_LC_11_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_adj_730_LC_11_19_4 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \c0.i1_3_lut_4_lut_adj_730_LC_11_19_4  (
            .in0(N__32892),
            .in1(N__32810),
            .in2(N__39219),
            .in3(N__33039),
            .lcout(\c0.n17076 ),
            .ltout(\c0.n17076_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i5_LC_11_19_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i5_LC_11_19_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i5_LC_11_19_5 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0__i5_LC_11_19_5  (
            .in0(N__37691),
            .in1(N__45132),
            .in2(N__32568),
            .in3(N__32750),
            .lcout(\c0.data_in_frame_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49700),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i53_LC_11_19_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i53_LC_11_19_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i53_LC_11_19_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.data_in_frame_0__i53_LC_11_19_6  (
            .in0(N__45130),
            .in1(N__32531),
            .in2(_gnd_net_),
            .in3(N__32565),
            .lcout(data_in_frame_6_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49700),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i10_LC_11_19_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i10_LC_11_19_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i10_LC_11_19_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i10_LC_11_19_7  (
            .in0(N__40577),
            .in1(N__40407),
            .in2(N__39998),
            .in3(N__39477),
            .lcout(\c0.data_in_frame_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49700),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_539_LC_11_20_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_539_LC_11_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_539_LC_11_20_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_539_LC_11_20_0  (
            .in0(_gnd_net_),
            .in1(N__34854),
            .in2(_gnd_net_),
            .in3(N__36947),
            .lcout(\c0.n10215 ),
            .ltout(\c0.n10215_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_526_LC_11_20_1 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_526_LC_11_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_526_LC_11_20_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_526_LC_11_20_1  (
            .in0(N__32745),
            .in1(N__34890),
            .in2(N__32724),
            .in3(N__34796),
            .lcout(\c0.n17206 ),
            .ltout(\c0.n17206_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1026_2_lut_3_lut_4_lut_LC_11_20_2 .C_ON=1'b0;
    defparam \c0.i1026_2_lut_3_lut_4_lut_LC_11_20_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1026_2_lut_3_lut_4_lut_LC_11_20_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1026_2_lut_3_lut_4_lut_LC_11_20_2  (
            .in0(N__37376),
            .in1(N__41030),
            .in2(N__32721),
            .in3(N__34763),
            .lcout(\c0.n2138 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i7_LC_11_20_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i7_LC_11_20_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i7_LC_11_20_3 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \c0.data_in_frame_0__i7_LC_11_20_3  (
            .in0(N__37730),
            .in1(N__34772),
            .in2(N__40433),
            .in3(N__39552),
            .lcout(\c0.data_in_frame_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49713),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_495_LC_11_20_4 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_495_LC_11_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_495_LC_11_20_4 .LUT_INIT=16'b1110111111011111;
    LogicCell40 \c0.i10_4_lut_adj_495_LC_11_20_4  (
            .in0(N__34980),
            .in1(N__32718),
            .in2(N__34522),
            .in3(N__40021),
            .lcout(\c0.n26_adj_2210 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i41_LC_11_20_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i41_LC_11_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i41_LC_11_20_5 .LUT_INIT=16'b1110111101000000;
    LogicCell40 \c0.data_in_frame_0__i41_LC_11_20_5  (
            .in0(N__40410),
            .in1(N__36802),
            .in2(N__32696),
            .in3(N__34959),
            .lcout(\c0.data_in_frame_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49713),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i3_LC_11_20_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i3_LC_11_20_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i3_LC_11_20_6 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i3_LC_11_20_6  (
            .in0(N__36876),
            .in1(N__40411),
            .in2(N__34865),
            .in3(N__37729),
            .lcout(\c0.data_in_frame_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49713),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i9_LC_11_20_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i9_LC_11_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i9_LC_11_20_7 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0__i9_LC_11_20_7  (
            .in0(N__40022),
            .in1(N__36803),
            .in2(N__40434),
            .in3(N__40618),
            .lcout(\c0.data_in_frame_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49713),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_491_LC_11_21_0 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_491_LC_11_21_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_491_LC_11_21_0 .LUT_INIT=16'b1011111001111101;
    LogicCell40 \c0.i2_4_lut_adj_491_LC_11_21_0  (
            .in0(N__37443),
            .in1(N__34820),
            .in2(N__33417),
            .in3(N__32618),
            .lcout(\c0.n18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_480_LC_11_21_1 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_480_LC_11_21_1 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_480_LC_11_21_1 .LUT_INIT=16'b1111011001101111;
    LogicCell40 \c0.i7_4_lut_adj_480_LC_11_21_1  (
            .in0(N__37396),
            .in1(N__39993),
            .in2(N__40989),
            .in3(N__37464),
            .lcout(),
            .ltout(\c0.n23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14_4_lut_LC_11_21_2 .C_ON=1'b0;
    defparam \c0.i14_4_lut_LC_11_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i14_4_lut_LC_11_21_2 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \c0.i14_4_lut_LC_11_21_2  (
            .in0(N__38892),
            .in1(N__34613),
            .in2(N__32967),
            .in3(N__34806),
            .lcout(),
            .ltout(\c0.n30_adj_2213_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15_4_lut_adj_517_LC_11_21_3 .C_ON=1'b0;
    defparam \c0.i15_4_lut_adj_517_LC_11_21_3 .SEQ_MODE=4'b0000;
    defparam \c0.i15_4_lut_adj_517_LC_11_21_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i15_4_lut_adj_517_LC_11_21_3  (
            .in0(N__32964),
            .in1(N__32958),
            .in2(N__32952),
            .in3(N__32949),
            .lcout(n31_adj_2415),
            .ltout(n31_adj_2415_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_3_lut_LC_11_21_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_3_lut_LC_11_21_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_3_lut_LC_11_21_4 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \c0.i1_2_lut_3_lut_3_lut_LC_11_21_4  (
            .in0(N__35743),
            .in1(_gnd_net_),
            .in2(N__32940),
            .in3(N__33437),
            .lcout(n1_adj_2486),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_651_LC_11_21_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_651_LC_11_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_651_LC_11_21_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_651_LC_11_21_5  (
            .in0(N__40988),
            .in1(N__32937),
            .in2(N__34869),
            .in3(N__36949),
            .lcout(\c0.n16352 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_635_LC_11_22_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_635_LC_11_22_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_635_LC_11_22_0 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \c0.i1_2_lut_adj_635_LC_11_22_0  (
            .in0(N__32916),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35026),
            .lcout(\c0.n6_adj_2358 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i27_LC_11_22_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i27_LC_11_22_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i27_LC_11_22_1 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0__i27_LC_11_22_1  (
            .in0(N__40610),
            .in1(N__34364),
            .in2(N__36862),
            .in3(N__39359),
            .lcout(\c0.data_in_frame_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49734),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_adj_726_LC_11_22_2 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_adj_726_LC_11_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_adj_726_LC_11_22_2 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \c0.i1_3_lut_4_lut_adj_726_LC_11_22_2  (
            .in0(N__32888),
            .in1(N__39200),
            .in2(N__32811),
            .in3(N__33013),
            .lcout(\c0.n17072 ),
            .ltout(\c0.n17072_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i21_LC_11_22_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i21_LC_11_22_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i21_LC_11_22_3 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0__i21_LC_11_22_3  (
            .in0(N__37733),
            .in1(N__45135),
            .in2(N__32769),
            .in3(N__33412),
            .lcout(\c0.data_in_frame_2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49734),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_620_LC_11_22_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_620_LC_11_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_adj_620_LC_11_22_4 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_adj_620_LC_11_22_4  (
            .in0(N__36072),
            .in1(N__40197),
            .in2(N__35745),
            .in3(N__35532),
            .lcout(FRAME_MATCHER_i_31__N_1273),
            .ltout(FRAME_MATCHER_i_31__N_1273_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_630_LC_11_22_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_630_LC_11_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_630_LC_11_22_5 .LUT_INIT=16'b1111000011110011;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_630_LC_11_22_5  (
            .in0(_gnd_net_),
            .in1(N__35723),
            .in2(N__33390),
            .in3(N__35817),
            .lcout(n17086),
            .ltout(n17086_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_626_LC_11_22_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_626_LC_11_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_626_LC_11_22_6 .LUT_INIT=16'b1111010111110000;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_626_LC_11_22_6  (
            .in0(N__35818),
            .in1(_gnd_net_),
            .in2(N__33387),
            .in3(N__35725),
            .lcout(\c0.n1034 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_641_LC_11_22_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_641_LC_11_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_641_LC_11_22_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.i1_2_lut_adj_641_LC_11_22_7  (
            .in0(_gnd_net_),
            .in1(N__35724),
            .in2(_gnd_net_),
            .in3(N__35819),
            .lcout(FRAME_MATCHER_i_31__N_1275),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4980_2_lut_LC_11_23_0 .C_ON=1'b0;
    defparam \c0.i4980_2_lut_LC_11_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i4980_2_lut_LC_11_23_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i4980_2_lut_LC_11_23_0  (
            .in0(_gnd_net_),
            .in1(N__33382),
            .in2(_gnd_net_),
            .in3(N__33360),
            .lcout(n10088),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_707_LC_11_23_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_707_LC_11_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_707_LC_11_23_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_707_LC_11_23_1  (
            .in0(_gnd_net_),
            .in1(N__33336),
            .in2(_gnd_net_),
            .in3(N__40702),
            .lcout(\c0.n16666 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_708_LC_11_23_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_708_LC_11_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_708_LC_11_23_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \c0.i1_2_lut_adj_708_LC_11_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__40711),
            .in3(N__33291),
            .lcout(\c0.n16674 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_644_LC_11_23_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_644_LC_11_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_644_LC_11_23_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i1_2_lut_adj_644_LC_11_23_3  (
            .in0(_gnd_net_),
            .in1(N__33553),
            .in2(_gnd_net_),
            .in3(N__33011),
            .lcout(n10140),
            .ltout(n10140_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_LC_11_23_4.C_ON=1'b0;
    defparam i1_3_lut_LC_11_23_4.SEQ_MODE=4'b0000;
    defparam i1_3_lut_LC_11_23_4.LUT_INIT=16'b0011111100001111;
    LogicCell40 i1_3_lut_LC_11_23_4 (
            .in0(_gnd_net_),
            .in1(N__41592),
            .in2(N__32970),
            .in3(N__44414),
            .lcout(n17089),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_629_LC_11_23_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_629_LC_11_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_629_LC_11_23_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \c0.i1_2_lut_adj_629_LC_11_23_5  (
            .in0(N__35704),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35820),
            .lcout(n44),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_753_LC_11_23_6 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_753_LC_11_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_753_LC_11_23_6 .LUT_INIT=16'b1111111100000100;
    LogicCell40 \c0.i1_4_lut_adj_753_LC_11_23_6  (
            .in0(N__35821),
            .in1(N__41445),
            .in2(N__35746),
            .in3(N__41296),
            .lcout(\c0.n8_adj_2385 ),
            .ltout(\c0.n8_adj_2385_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_716_LC_11_23_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_716_LC_11_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_716_LC_11_23_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \c0.i1_2_lut_adj_716_LC_11_23_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33585),
            .in3(N__37809),
            .lcout(\c0.n16670 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14591_2_lut_LC_11_24_0 .C_ON=1'b0;
    defparam \c0.i14591_2_lut_LC_11_24_0 .SEQ_MODE=4'b0000;
    defparam \c0.i14591_2_lut_LC_11_24_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i14591_2_lut_LC_11_24_0  (
            .in0(_gnd_net_),
            .in1(N__40198),
            .in2(_gnd_net_),
            .in3(N__35534),
            .lcout(),
            .ltout(\c0.n17367_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_418_LC_11_24_1 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_418_LC_11_24_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_418_LC_11_24_1 .LUT_INIT=16'b1010111110101110;
    LogicCell40 \c0.i1_4_lut_adj_418_LC_11_24_1  (
            .in0(N__42014),
            .in1(N__35702),
            .in2(N__33561),
            .in3(N__36061),
            .lcout(\c0.n10139 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_751_LC_11_24_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_751_LC_11_24_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_751_LC_11_24_2 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_751_LC_11_24_2  (
            .in0(N__36062),
            .in1(N__40199),
            .in2(_gnd_net_),
            .in3(N__35535),
            .lcout(n9),
            .ltout(n9_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_adj_698_LC_11_24_3 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_adj_698_LC_11_24_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_adj_698_LC_11_24_3 .LUT_INIT=16'b0000100011111111;
    LogicCell40 \c0.i1_3_lut_4_lut_adj_698_LC_11_24_3  (
            .in0(N__39753),
            .in1(N__35703),
            .in2(N__33558),
            .in3(N__33555),
            .lcout(\c0.n11833 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i20_4_lut_LC_11_24_4 .C_ON=1'b0;
    defparam \c0.i20_4_lut_LC_11_24_4 .SEQ_MODE=4'b0000;
    defparam \c0.i20_4_lut_LC_11_24_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i20_4_lut_LC_11_24_4  (
            .in0(N__33489),
            .in1(N__33793),
            .in2(N__40761),
            .in3(N__33470),
            .lcout(\c0.n49 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_797_LC_11_24_5.C_ON=1'b0;
    defparam i1_4_lut_adj_797_LC_11_24_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_797_LC_11_24_5.LUT_INIT=16'b1111000000010000;
    LogicCell40 i1_4_lut_adj_797_LC_11_24_5 (
            .in0(N__39754),
            .in1(N__33436),
            .in2(N__35744),
            .in3(N__35463),
            .lcout(),
            .ltout(n21_adj_2487_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i1_LC_11_24_6 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i1_LC_11_24_6 .SEQ_MODE=4'b1000;
    defparam \c0.FRAME_MATCHER_state_i1_LC_11_24_6 .LUT_INIT=16'b1111111111110100;
    LogicCell40 \c0.FRAME_MATCHER_state_i1_LC_11_24_6  (
            .in0(N__41389),
            .in1(N__33702),
            .in2(N__33747),
            .in3(N__33708),
            .lcout(FRAME_MATCHER_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49757),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_adj_798_LC_11_24_7.C_ON=1'b0;
    defparam i2_4_lut_adj_798_LC_11_24_7.SEQ_MODE=4'b0000;
    defparam i2_4_lut_adj_798_LC_11_24_7.LUT_INIT=16'b1010000011101100;
    LogicCell40 i2_4_lut_adj_798_LC_11_24_7 (
            .in0(N__35904),
            .in1(N__35462),
            .in2(N__35958),
            .in3(N__33744),
            .lcout(n6_adj_2410),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i7_LC_11_25_2 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i7_LC_11_25_2 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i7_LC_11_25_2 .LUT_INIT=16'b1110000011000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i7_LC_11_25_2  (
            .in0(N__44945),
            .in1(N__44772),
            .in2(N__33798),
            .in3(N__44564),
            .lcout(\c0.FRAME_MATCHER_state_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49770),
            .ce(),
            .sr(N__33777));
    defparam i14574_2_lut_3_lut_LC_11_25_4.C_ON=1'b0;
    defparam i14574_2_lut_3_lut_LC_11_25_4.SEQ_MODE=4'b0000;
    defparam i14574_2_lut_3_lut_LC_11_25_4.LUT_INIT=16'b1111111111101110;
    LogicCell40 i14574_2_lut_3_lut_LC_11_25_4 (
            .in0(N__35712),
            .in1(N__33698),
            .in2(_gnd_net_),
            .in3(N__35828),
            .lcout(n17349),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_428_LC_11_25_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_428_LC_11_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_428_LC_11_25_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.i1_2_lut_adj_428_LC_11_25_5  (
            .in0(_gnd_net_),
            .in1(N__35711),
            .in2(_gnd_net_),
            .in3(N__35551),
            .lcout(\c0.n51_adj_2173 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_420_LC_11_25_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_420_LC_11_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_420_LC_11_25_6 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \c0.i1_2_lut_adj_420_LC_11_25_6  (
            .in0(N__35552),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40239),
            .lcout(\c0.n10166 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10658_2_lut_LC_11_25_7 .C_ON=1'b0;
    defparam \c0.i10658_2_lut_LC_11_25_7 .SEQ_MODE=4'b0000;
    defparam \c0.i10658_2_lut_LC_11_25_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i10658_2_lut_LC_11_25_7  (
            .in0(_gnd_net_),
            .in1(N__33656),
            .in2(_gnd_net_),
            .in3(N__41741),
            .lcout(\c0.FRAME_MATCHER_i_31_N_1310_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_765_LC_11_26_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_765_LC_11_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_765_LC_11_26_0 .LUT_INIT=16'b1010101000001000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_765_LC_11_26_0  (
            .in0(N__35210),
            .in1(N__41472),
            .in2(N__41423),
            .in3(N__41333),
            .lcout(\c0.n16696 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i1_LC_11_26_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i1_LC_11_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i1_LC_11_26_1 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \c0.byte_transmit_counter__i1_LC_11_26_1  (
            .in0(N__47438),
            .in1(N__42912),
            .in2(N__42446),
            .in3(N__42367),
            .lcout(byte_transmit_counter_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49782),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_745_LC_11_26_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_745_LC_11_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_745_LC_11_26_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_745_LC_11_26_2  (
            .in0(N__49170),
            .in1(N__47120),
            .in2(_gnd_net_),
            .in3(N__49099),
            .lcout(\c0.n17270 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i6_LC_11_26_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i6_LC_11_26_3 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i6_LC_11_26_3 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \c0.byte_transmit_counter__i6_LC_11_26_3  (
            .in0(N__42716),
            .in1(N__42945),
            .in2(N__42448),
            .in3(N__42369),
            .lcout(byte_transmit_counter_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49782),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_8__2__2190_LC_11_26_4 .C_ON=1'b0;
    defparam \c0.data_out_8__2__2190_LC_11_26_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_8__2__2190_LC_11_26_4 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_out_8__2__2190_LC_11_26_4  (
            .in0(N__33830),
            .in1(_gnd_net_),
            .in2(N__49962),
            .in3(N__48718),
            .lcout(data_out_8_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49782),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i3_LC_11_26_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i3_LC_11_26_5 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i3_LC_11_26_5 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \c0.byte_transmit_counter__i3_LC_11_26_5  (
            .in0(N__43050),
            .in1(N__46379),
            .in2(N__42447),
            .in3(N__42368),
            .lcout(byte_transmit_counter_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49782),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_8__3__2189_LC_11_26_6 .C_ON=1'b0;
    defparam \c0.data_out_8__3__2189_LC_11_26_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_8__3__2189_LC_11_26_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_8__3__2189_LC_11_26_6  (
            .in0(N__49930),
            .in1(N__33816),
            .in2(_gnd_net_),
            .in3(N__48825),
            .lcout(data_out_8_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49782),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13368_2_lut_LC_11_26_7 .C_ON=1'b0;
    defparam \c0.i13368_2_lut_LC_11_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.i13368_2_lut_LC_11_26_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i13368_2_lut_LC_11_26_7  (
            .in0(_gnd_net_),
            .in1(N__33794),
            .in2(_gnd_net_),
            .in3(N__40807),
            .lcout(\c0.n16141 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__7__2201_LC_11_27_0 .C_ON=1'b0;
    defparam \c0.data_out_6__7__2201_LC_11_27_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__7__2201_LC_11_27_0 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \c0.data_out_6__7__2201_LC_11_27_0  (
            .in0(N__50150),
            .in1(N__33765),
            .in2(N__48157),
            .in3(N__42474),
            .lcout(\c0.data_out_6_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49792),
            .ce(N__50588),
            .sr(_gnd_net_));
    defparam \c0.data_out_1__1__2247_LC_11_27_1 .C_ON=1'b0;
    defparam \c0.data_out_1__1__2247_LC_11_27_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_1__1__2247_LC_11_27_1 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \c0.data_out_1__1__2247_LC_11_27_1  (
            .in0(N__48381),
            .in1(N__48121),
            .in2(_gnd_net_),
            .in3(N__50151),
            .lcout(\c0.data_out_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49792),
            .ce(N__50588),
            .sr(_gnd_net_));
    defparam \c0.i15145_3_lut_LC_11_27_3 .C_ON=1'b0;
    defparam \c0.i15145_3_lut_LC_11_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.i15145_3_lut_LC_11_27_3 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \c0.i15145_3_lut_LC_11_27_3  (
            .in0(N__45733),
            .in1(N__48380),
            .in2(_gnd_net_),
            .in3(N__47119),
            .lcout(),
            .ltout(\c0.n17639_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__4__2204_LC_11_27_4 .C_ON=1'b0;
    defparam \c0.data_out_6__4__2204_LC_11_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__4__2204_LC_11_27_4 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \c0.data_out_6__4__2204_LC_11_27_4  (
            .in0(N__48123),
            .in1(N__50153),
            .in2(N__33948),
            .in3(N__33944),
            .lcout(\c0.data_out_6_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49792),
            .ce(N__50588),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__6__2202_LC_11_27_5 .C_ON=1'b0;
    defparam \c0.data_out_6__6__2202_LC_11_27_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__6__2202_LC_11_27_5 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \c0.data_out_6__6__2202_LC_11_27_5  (
            .in0(N__33929),
            .in1(N__48122),
            .in2(N__33915),
            .in3(N__50152),
            .lcout(\c0.data_out_6_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49792),
            .ce(N__50588),
            .sr(_gnd_net_));
    defparam \c0.i15088_2_lut_LC_11_27_6 .C_ON=1'b0;
    defparam \c0.i15088_2_lut_LC_11_27_6 .SEQ_MODE=4'b0000;
    defparam \c0.i15088_2_lut_LC_11_27_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i15088_2_lut_LC_11_27_6  (
            .in0(_gnd_net_),
            .in1(N__45732),
            .in2(_gnd_net_),
            .in3(N__47700),
            .lcout(\c0.n17671 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14999_3_lut_LC_11_28_0 .C_ON=1'b0;
    defparam \c0.i14999_3_lut_LC_11_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.i14999_3_lut_LC_11_28_0 .LUT_INIT=16'b0101000010100000;
    LogicCell40 \c0.i14999_3_lut_LC_11_28_0  (
            .in0(N__45728),
            .in1(_gnd_net_),
            .in2(N__48418),
            .in3(N__47877),
            .lcout(),
            .ltout(\c0.n17631_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__3__2205_LC_11_28_1 .C_ON=1'b0;
    defparam \c0.data_out_6__3__2205_LC_11_28_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__3__2205_LC_11_28_1 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \c0.data_out_6__3__2205_LC_11_28_1  (
            .in0(N__33899),
            .in1(N__48128),
            .in2(N__33885),
            .in3(N__50157),
            .lcout(\c0.data_out_6_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49802),
            .ce(N__50566),
            .sr(_gnd_net_));
    defparam \c0.i15033_3_lut_LC_11_28_2 .C_ON=1'b0;
    defparam \c0.i15033_3_lut_LC_11_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.i15033_3_lut_LC_11_28_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \c0.i15033_3_lut_LC_11_28_2  (
            .in0(N__48392),
            .in1(N__43362),
            .in2(_gnd_net_),
            .in3(N__47876),
            .lcout(),
            .ltout(\c0.n17627_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__2__2206_LC_11_28_3 .C_ON=1'b0;
    defparam \c0.data_out_6__2__2206_LC_11_28_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__2__2206_LC_11_28_3 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \c0.data_out_6__2__2206_LC_11_28_3  (
            .in0(N__33881),
            .in1(N__48127),
            .in2(N__33867),
            .in3(N__50156),
            .lcout(\c0.data_out_6_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49802),
            .ce(N__50566),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__5__2203_LC_11_28_5 .C_ON=1'b0;
    defparam \c0.data_out_6__5__2203_LC_11_28_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__5__2203_LC_11_28_5 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \c0.data_out_6__5__2203_LC_11_28_5  (
            .in0(N__33863),
            .in1(N__48129),
            .in2(N__33849),
            .in3(N__50158),
            .lcout(\c0.data_out_6_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49802),
            .ce(N__50566),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_720_LC_11_28_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_720_LC_11_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_720_LC_11_28_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_720_LC_11_28_6  (
            .in0(N__45727),
            .in1(N__43361),
            .in2(_gnd_net_),
            .in3(N__47875),
            .lcout(\c0.n10326 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_LC_11_29_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_LC_11_29_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_LC_11_29_0 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter_1__bdd_4_lut_LC_11_29_0  (
            .in0(N__33954),
            .in1(N__46252),
            .in2(N__33993),
            .in3(N__47482),
            .lcout(),
            .ltout(\c0.n18268_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18268_bdd_4_lut_LC_11_29_1 .C_ON=1'b0;
    defparam \c0.n18268_bdd_4_lut_LC_11_29_1 .SEQ_MODE=4'b0000;
    defparam \c0.n18268_bdd_4_lut_LC_11_29_1 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n18268_bdd_4_lut_LC_11_29_1  (
            .in0(N__46253),
            .in1(N__34035),
            .in2(N__33999),
            .in3(N__34080),
            .lcout(n18271),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_2_lut_3_lut_LC_11_29_2 .C_ON=1'b0;
    defparam \c0.tx.i1_2_lut_3_lut_LC_11_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_2_lut_3_lut_LC_11_29_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.tx.i1_2_lut_3_lut_LC_11_29_2  (
            .in0(N__42640),
            .in1(N__42583),
            .in2(_gnd_net_),
            .in3(N__36370),
            .lcout(),
            .ltout(\c0.tx.n55_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_i2_LC_11_29_3 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_i2_LC_11_29_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Bit_Index_i2_LC_11_29_3 .LUT_INIT=16'b0001110111000000;
    LogicCell40 \c0.tx.r_Bit_Index_i2_LC_11_29_3  (
            .in0(N__36371),
            .in1(N__44214),
            .in2(N__33996),
            .in3(N__42550),
            .lcout(r_Bit_Index_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49809),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i5_3_lut_LC_11_29_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i5_3_lut_LC_11_29_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i5_3_lut_LC_11_29_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_4_i5_3_lut_LC_11_29_4  (
            .in0(N__48963),
            .in1(N__45646),
            .in2(_gnd_net_),
            .in3(N__47670),
            .lcout(\c0.n5_adj_2136 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_1_i8_3_lut_LC_11_29_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_1_i8_3_lut_LC_11_29_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_1_i8_3_lut_LC_11_29_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_1_i8_3_lut_LC_11_29_5  (
            .in0(N__47669),
            .in1(N__48573),
            .in2(_gnd_net_),
            .in3(N__42129),
            .lcout(n8_adj_2447),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__4__2196_LC_11_29_6 .C_ON=1'b0;
    defparam \c0.data_out_7__4__2196_LC_11_29_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__4__2196_LC_11_29_6 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \c0.data_out_7__4__2196_LC_11_29_6  (
            .in0(N__48964),
            .in1(N__33984),
            .in2(N__43718),
            .in3(N__46905),
            .lcout(\c0.data_out_7_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49809),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15376_LC_11_30_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15376_LC_11_30_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15376_LC_11_30_0 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter_1__bdd_4_lut_15376_LC_11_30_0  (
            .in0(N__34050),
            .in1(N__46250),
            .in2(N__33966),
            .in3(N__47481),
            .lcout(),
            .ltout(\c0.n18172_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18172_bdd_4_lut_LC_11_30_1 .C_ON=1'b0;
    defparam \c0.n18172_bdd_4_lut_LC_11_30_1 .SEQ_MODE=4'b0000;
    defparam \c0.n18172_bdd_4_lut_LC_11_30_1 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n18172_bdd_4_lut_LC_11_30_1  (
            .in0(N__46251),
            .in1(N__36444),
            .in2(N__33957),
            .in3(N__34029),
            .lcout(n18175),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15173_2_lut_LC_11_30_2 .C_ON=1'b0;
    defparam \c0.i15173_2_lut_LC_11_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.i15173_2_lut_LC_11_30_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i15173_2_lut_LC_11_30_2  (
            .in0(N__47673),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49065),
            .lcout(\c0.n17764 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15100_2_lut_LC_11_30_3 .C_ON=1'b0;
    defparam \c0.i15100_2_lut_LC_11_30_3 .SEQ_MODE=4'b0000;
    defparam \c0.i15100_2_lut_LC_11_30_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i15100_2_lut_LC_11_30_3  (
            .in0(_gnd_net_),
            .in1(N__47675),
            .in2(_gnd_net_),
            .in3(N__34200),
            .lcout(\c0.n17676 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__6__2194_LC_11_30_4 .C_ON=1'b0;
    defparam \c0.data_out_7__6__2194_LC_11_30_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__6__2194_LC_11_30_4 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \c0.data_out_7__6__2194_LC_11_30_4  (
            .in0(N__47230),
            .in1(N__43693),
            .in2(N__34074),
            .in3(N__46918),
            .lcout(\c0.data_out_7_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49817),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15108_2_lut_LC_11_30_5 .C_ON=1'b0;
    defparam \c0.i15108_2_lut_LC_11_30_5 .SEQ_MODE=4'b0000;
    defparam \c0.i15108_2_lut_LC_11_30_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i15108_2_lut_LC_11_30_5  (
            .in0(_gnd_net_),
            .in1(N__47672),
            .in2(_gnd_net_),
            .in3(N__47085),
            .lcout(\c0.n17703 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_1__4__2244_LC_11_30_6 .C_ON=1'b0;
    defparam \c0.data_out_1__4__2244_LC_11_30_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_1__4__2244_LC_11_30_6 .LUT_INIT=16'b0000101000111010;
    LogicCell40 \c0.data_out_1__4__2244_LC_11_30_6  (
            .in0(N__34044),
            .in1(N__48388),
            .in2(N__50576),
            .in3(N__50266),
            .lcout(\c0.data_out_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49817),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15103_2_lut_LC_11_30_7 .C_ON=1'b0;
    defparam \c0.i15103_2_lut_LC_11_30_7 .SEQ_MODE=4'b0000;
    defparam \c0.i15103_2_lut_LC_11_30_7 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \c0.i15103_2_lut_LC_11_30_7  (
            .in0(_gnd_net_),
            .in1(N__47674),
            .in2(_gnd_net_),
            .in3(N__34043),
            .lcout(\c0.n17675 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15101_2_lut_LC_11_31_0 .C_ON=1'b0;
    defparam \c0.i15101_2_lut_LC_11_31_0 .SEQ_MODE=4'b0000;
    defparam \c0.i15101_2_lut_LC_11_31_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \c0.i15101_2_lut_LC_11_31_0  (
            .in0(N__47740),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34007),
            .lcout(\c0.n17697 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_4_lut_adj_784_LC_11_31_4.C_ON=1'b0;
    defparam i24_4_lut_adj_784_LC_11_31_4.SEQ_MODE=4'b0000;
    defparam i24_4_lut_adj_784_LC_11_31_4.LUT_INIT=16'b0010001011100010;
    LogicCell40 i24_4_lut_adj_784_LC_11_31_4 (
            .in0(N__34020),
            .in1(N__46400),
            .in2(N__47352),
            .in3(N__46288),
            .lcout(),
            .ltout(n10_adj_2408_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i4_LC_11_31_5 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i4_LC_11_31_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i4_LC_11_31_5 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \c0.tx.r_Tx_Data_i4_LC_11_31_5  (
            .in0(N__44104),
            .in1(N__38249),
            .in2(N__34011),
            .in3(N__43841),
            .lcout(r_Tx_Data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49824),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_2__3__2237_LC_11_31_7 .C_ON=1'b0;
    defparam \c0.data_out_2__3__2237_LC_11_31_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_2__3__2237_LC_11_31_7 .LUT_INIT=16'b0010001000101110;
    LogicCell40 \c0.data_out_2__3__2237_LC_11_31_7  (
            .in0(N__34008),
            .in1(N__50505),
            .in2(N__48417),
            .in3(N__50320),
            .lcout(\c0.data_out_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49824),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_3__0__2232_LC_11_32_0 .C_ON=1'b0;
    defparam \c0.data_out_3__0__2232_LC_11_32_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_3__0__2232_LC_11_32_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \c0.data_out_3__0__2232_LC_11_32_0  (
            .in0(N__35858),
            .in1(N__50555),
            .in2(_gnd_net_),
            .in3(N__34184),
            .lcout(data_out_3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49830),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__5__2251_LC_11_32_1 .C_ON=1'b0;
    defparam \c0.data_out_0__5__2251_LC_11_32_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__5__2251_LC_11_32_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_out_0__5__2251_LC_11_32_1  (
            .in0(N__34183),
            .in1(N__50552),
            .in2(_gnd_net_),
            .in3(N__34227),
            .lcout(data_out_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49830),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_2__2__2238_LC_11_32_2 .C_ON=1'b0;
    defparam \c0.data_out_2__2__2238_LC_11_32_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_2__2__2238_LC_11_32_2 .LUT_INIT=16'b0111011101000100;
    LogicCell40 \c0.data_out_2__2__2238_LC_11_32_2  (
            .in0(N__50329),
            .in1(N__50554),
            .in2(_gnd_net_),
            .in3(N__34215),
            .lcout(data_out_2_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49830),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.mux_1195_i1_3_lut_LC_11_32_3 .C_ON=1'b0;
    defparam \c0.mux_1195_i1_3_lut_LC_11_32_3 .SEQ_MODE=4'b0000;
    defparam \c0.mux_1195_i1_3_lut_LC_11_32_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.mux_1195_i1_3_lut_LC_11_32_3  (
            .in0(N__48384),
            .in1(N__48133),
            .in2(_gnd_net_),
            .in3(N__50328),
            .lcout(n2699),
            .ltout(n2699_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_3__4__2228_LC_11_32_4 .C_ON=1'b0;
    defparam \c0.data_out_3__4__2228_LC_11_32_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_3__4__2228_LC_11_32_4 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \c0.data_out_3__4__2228_LC_11_32_4  (
            .in0(_gnd_net_),
            .in1(N__50556),
            .in2(N__34203),
            .in3(N__34199),
            .lcout(data_out_3_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49830),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_3__2__2230_LC_11_32_7 .C_ON=1'b0;
    defparam \c0.data_out_3__2__2230_LC_11_32_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_3__2__2230_LC_11_32_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_out_3__2__2230_LC_11_32_7  (
            .in0(N__34185),
            .in1(N__50553),
            .in2(_gnd_net_),
            .in3(N__34173),
            .lcout(data_out_3_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49830),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i23_LC_12_15_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i23_LC_12_15_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i23_LC_12_15_7 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0__i23_LC_12_15_7  (
            .in0(N__37745),
            .in1(N__34153),
            .in2(N__39555),
            .in3(N__39390),
            .lcout(\c0.data_in_frame_2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49714),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_i6_LC_12_16_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_i6_LC_12_16_0 .SEQ_MODE=4'b1001;
    defparam \c0.byte_transmit_counter2_i6_LC_12_16_0 .LUT_INIT=16'b1100101000000000;
    LogicCell40 \c0.byte_transmit_counter2_i6_LC_12_16_0  (
            .in0(N__34131),
            .in1(N__34442),
            .in2(N__39701),
            .in3(N__42053),
            .lcout(\c0.byte_transmit_counter2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49701),
            .ce(),
            .sr(N__34119));
    defparam \c0.i10953_1_lut_LC_12_17_0 .C_ON=1'b0;
    defparam \c0.i10953_1_lut_LC_12_17_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10953_1_lut_LC_12_17_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \c0.i10953_1_lut_LC_12_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34409),
            .lcout(\c0.tx2_transmit_N_1996 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_756_LC_12_17_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_756_LC_12_17_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_756_LC_12_17_1 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_756_LC_12_17_1  (
            .in0(N__34410),
            .in1(N__34397),
            .in2(N__35765),
            .in3(N__35583),
            .lcout(\c0.n16261 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_537_LC_12_17_2 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_537_LC_12_17_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_537_LC_12_17_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i3_4_lut_adj_537_LC_12_17_2  (
            .in0(N__34484),
            .in1(N__34437),
            .in2(N__39622),
            .in3(N__34416),
            .lcout(\c0.n13628 ),
            .ltout(\c0.n13628_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_687_LC_12_17_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_687_LC_12_17_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_687_LC_12_17_3 .LUT_INIT=16'b1111111111001111;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_687_LC_12_17_3  (
            .in0(_gnd_net_),
            .in1(N__35582),
            .in2(N__34401),
            .in3(N__34396),
            .lcout(n488),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_4_lut_adj_601_LC_12_18_0 .C_ON=1'b0;
    defparam \c0.i7_4_lut_adj_601_LC_12_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.i7_4_lut_adj_601_LC_12_18_0 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \c0.i7_4_lut_adj_601_LC_12_18_0  (
            .in0(N__34368),
            .in1(N__34238),
            .in2(N__35346),
            .in3(N__36921),
            .lcout(\c0.n21_adj_2323 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_624_LC_12_18_1 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_624_LC_12_18_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_624_LC_12_18_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_624_LC_12_18_1  (
            .in0(N__41033),
            .in1(N__37045),
            .in2(N__34350),
            .in3(N__36954),
            .lcout(\c0.n16353 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14698_4_lut_LC_12_18_2 .C_ON=1'b0;
    defparam \c0.i14698_4_lut_LC_12_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.i14698_4_lut_LC_12_18_2 .LUT_INIT=16'b1111110010110000;
    LogicCell40 \c0.i14698_4_lut_LC_12_18_2  (
            .in0(N__40316),
            .in1(N__39825),
            .in2(N__34314),
            .in3(N__40144),
            .lcout(),
            .ltout(\c0.n17475_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i6_LC_12_18_3 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i6_LC_12_18_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i6_LC_12_18_3 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \c0.data_out_frame2_0___i6_LC_12_18_3  (
            .in0(N__39826),
            .in1(N__39934),
            .in2(N__34329),
            .in3(N__39877),
            .lcout(\c0.data_out_frame2_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49702),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_662_LC_12_18_4 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_662_LC_12_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_662_LC_12_18_4 .LUT_INIT=16'b1101111111111101;
    LogicCell40 \c0.i12_4_lut_adj_662_LC_12_18_4  (
            .in0(N__34281),
            .in1(N__34269),
            .in2(N__34263),
            .in3(N__34239),
            .lcout(\c0.n28_adj_2374 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14692_4_lut_LC_12_18_6 .C_ON=1'b0;
    defparam \c0.i14692_4_lut_LC_12_18_6 .SEQ_MODE=4'b0000;
    defparam \c0.i14692_4_lut_LC_12_18_6 .LUT_INIT=16'b1111110010110000;
    LogicCell40 \c0.i14692_4_lut_LC_12_18_6  (
            .in0(N__40315),
            .in1(N__39824),
            .in2(N__34714),
            .in3(N__40143),
            .lcout(),
            .ltout(\c0.n17469_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i8_LC_12_18_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i8_LC_12_18_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i8_LC_12_18_7 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \c0.data_out_frame2_0___i8_LC_12_18_7  (
            .in0(N__39827),
            .in1(N__39935),
            .in2(N__34728),
            .in3(N__39878),
            .lcout(\c0.data_out_frame2_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49702),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_563_LC_12_19_0 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_563_LC_12_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_563_LC_12_19_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_4_lut_adj_563_LC_12_19_0  (
            .in0(N__37043),
            .in1(N__34529),
            .in2(N__34680),
            .in3(N__34562),
            .lcout(),
            .ltout(\c0.n17114_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_643_LC_12_19_1 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_643_LC_12_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_643_LC_12_19_1 .LUT_INIT=16'b1111100111110110;
    LogicCell40 \c0.i2_4_lut_adj_643_LC_12_19_1  (
            .in0(N__37378),
            .in1(N__34659),
            .in2(N__34641),
            .in3(N__40020),
            .lcout(\c0.n18_adj_2360 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_623_LC_12_19_2 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_623_LC_12_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_623_LC_12_19_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_623_LC_12_19_2  (
            .in0(N__37044),
            .in1(N__40953),
            .in2(N__34638),
            .in3(N__34563),
            .lcout(\c0.n17214 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_546_LC_12_19_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_546_LC_12_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_546_LC_12_19_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_546_LC_12_19_3  (
            .in0(_gnd_net_),
            .in1(N__40019),
            .in2(_gnd_net_),
            .in3(N__39983),
            .lcout(),
            .ltout(\c0.n17101_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_547_LC_12_19_4 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_547_LC_12_19_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_547_LC_12_19_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_547_LC_12_19_4  (
            .in0(N__34607),
            .in1(N__34771),
            .in2(N__34581),
            .in3(N__37377),
            .lcout(),
            .ltout(\c0.n10_adj_2299_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_554_LC_12_19_5 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_554_LC_12_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_554_LC_12_19_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_554_LC_12_19_5  (
            .in0(N__38828),
            .in1(N__38900),
            .in2(N__34578),
            .in3(N__34575),
            .lcout(\c0.n10407 ),
            .ltout(\c0.n10407_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_604_LC_12_19_6 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_604_LC_12_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_604_LC_12_19_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_4_lut_adj_604_LC_12_19_6  (
            .in0(N__34554),
            .in1(N__40952),
            .in2(N__34533),
            .in3(N__34530),
            .lcout(\c0.n17215 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i8_LC_12_19_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i8_LC_12_19_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i8_LC_12_19_7 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.data_in_frame_0__i8_LC_12_19_7  (
            .in0(N__37379),
            .in1(N__37728),
            .in2(N__40502),
            .in3(N__40426),
            .lcout(\c0.data_in_frame_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49715),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1016_2_lut_LC_12_20_0 .C_ON=1'b0;
    defparam \c0.i1016_2_lut_LC_12_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1016_2_lut_LC_12_20_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1016_2_lut_LC_12_20_0  (
            .in0(_gnd_net_),
            .in1(N__34764),
            .in2(_gnd_net_),
            .in3(N__37380),
            .lcout(\c0.n2128 ),
            .ltout(\c0.n2128_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_602_LC_12_20_1 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_602_LC_12_20_1 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_602_LC_12_20_1 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \c0.i3_4_lut_adj_602_LC_12_20_1  (
            .in0(N__34973),
            .in1(N__34958),
            .in2(N__34947),
            .in3(N__37502),
            .lcout(\c0.n19_adj_2324 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__0__2269_LC_12_20_2 .C_ON=1'b0;
    defparam \c0.data_in_3__0__2269_LC_12_20_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__0__2269_LC_12_20_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_3__0__2269_LC_12_20_2  (
            .in0(N__36804),
            .in1(N__39194),
            .in2(_gnd_net_),
            .in3(N__34923),
            .lcout(data_in_3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49725),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1008_2_lut_LC_12_20_3 .C_ON=1'b0;
    defparam \c0.i1008_2_lut_LC_12_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1008_2_lut_LC_12_20_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1008_2_lut_LC_12_20_3  (
            .in0(_gnd_net_),
            .in1(N__34894),
            .in2(_gnd_net_),
            .in3(N__34855),
            .lcout(\c0.n2120 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_3_lut_4_lut_LC_12_20_4 .C_ON=1'b0;
    defparam \c0.i6_3_lut_4_lut_LC_12_20_4 .SEQ_MODE=4'b0000;
    defparam \c0.i6_3_lut_4_lut_LC_12_20_4 .LUT_INIT=16'b1001111101101111;
    LogicCell40 \c0.i6_3_lut_4_lut_LC_12_20_4  (
            .in0(N__34797),
            .in1(N__36898),
            .in2(N__37047),
            .in3(N__34765),
            .lcout(),
            .ltout(\c0.n22_adj_2201_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_482_LC_12_20_5 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_482_LC_12_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_482_LC_12_20_5 .LUT_INIT=16'b1111011111111011;
    LogicCell40 \c0.i11_4_lut_adj_482_LC_12_20_5  (
            .in0(N__37417),
            .in1(N__38827),
            .in2(N__34809),
            .in3(N__36917),
            .lcout(\c0.n27_adj_2202 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1014_2_lut_LC_12_20_6 .C_ON=1'b0;
    defparam \c0.i1014_2_lut_LC_12_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1014_2_lut_LC_12_20_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1014_2_lut_LC_12_20_6  (
            .in0(N__34798),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34766),
            .lcout(\c0.n2126 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i2_LC_12_20_7 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i2_LC_12_20_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i2_LC_12_20_7 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \c0.data_in_frame_0__i2_LC_12_20_7  (
            .in0(N__37731),
            .in1(N__40423),
            .in2(N__39469),
            .in3(N__36953),
            .lcout(\c0.data_in_frame_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49725),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i17_LC_12_21_0 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i17_LC_12_21_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i17_LC_12_21_0 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i17_LC_12_21_0  (
            .in0(N__37732),
            .in1(N__36798),
            .in2(N__35119),
            .in3(N__39360),
            .lcout(\c0.data_in_frame_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49735),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i2_LC_12_21_1 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i2_LC_12_21_1 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i2_LC_12_21_1 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.rx.r_Rx_Byte_i2_LC_12_21_1  (
            .in0(N__37973),
            .in1(N__45258),
            .in2(N__36861),
            .in3(N__45156),
            .lcout(rx_data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49735),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_4_lut_adj_677_LC_12_21_2 .C_ON=1'b0;
    defparam \c0.i1_3_lut_4_lut_adj_677_LC_12_21_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_4_lut_adj_677_LC_12_21_2 .LUT_INIT=16'b0100000001000100;
    LogicCell40 \c0.i1_3_lut_4_lut_adj_677_LC_12_21_2  (
            .in0(N__35550),
            .in1(N__35750),
            .in2(N__36093),
            .in3(N__40235),
            .lcout(\c0.n5817 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__6__2263_LC_12_21_4 .C_ON=1'b0;
    defparam \c0.data_in_3__6__2263_LC_12_21_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__6__2263_LC_12_21_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_3__6__2263_LC_12_21_4  (
            .in0(N__39541),
            .in1(N__39094),
            .in2(_gnd_net_),
            .in3(N__35074),
            .lcout(data_in_3_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49735),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_691_LC_12_21_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_691_LC_12_21_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_691_LC_12_21_5 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_691_LC_12_21_5  (
            .in0(N__40234),
            .in1(N__36086),
            .in2(N__35758),
            .in3(N__35549),
            .lcout(\c0.n5815 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10706_2_lut_LC_12_21_6 .C_ON=1'b0;
    defparam \c0.i10706_2_lut_LC_12_21_6 .SEQ_MODE=4'b0000;
    defparam \c0.i10706_2_lut_LC_12_21_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i10706_2_lut_LC_12_21_6  (
            .in0(_gnd_net_),
            .in1(N__37327),
            .in2(_gnd_net_),
            .in3(N__40814),
            .lcout(\c0.n13381 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_0__0__2293_LC_12_21_7 .C_ON=1'b0;
    defparam \c0.data_in_0__0__2293_LC_12_21_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_0__0__2293_LC_12_21_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_0__0__2293_LC_12_21_7  (
            .in0(N__39093),
            .in1(N__35030),
            .in2(_gnd_net_),
            .in3(N__35055),
            .lcout(data_in_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49735),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_794_LC_12_22_0.C_ON=1'b0;
    defparam i1_4_lut_adj_794_LC_12_22_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_794_LC_12_22_0.LUT_INIT=16'b1110111011101010;
    LogicCell40 i1_4_lut_adj_794_LC_12_22_0 (
            .in0(N__35786),
            .in1(N__44424),
            .in2(N__41613),
            .in3(N__36109),
            .lcout(n6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__1__2268_LC_12_22_1 .C_ON=1'b0;
    defparam \c0.data_in_3__1__2268_LC_12_22_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__1__2268_LC_12_22_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \c0.data_in_3__1__2268_LC_12_22_1  (
            .in0(N__39205),
            .in1(_gnd_net_),
            .in2(N__39478),
            .in3(N__34999),
            .lcout(data_in_3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49746),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i1_LC_12_22_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i1_LC_12_22_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i1_LC_12_22_2 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i1_LC_12_22_2  (
            .in0(N__37734),
            .in1(N__36799),
            .in2(N__41034),
            .in3(N__40432),
            .lcout(\c0.data_in_frame_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49746),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_1__1__2284_LC_12_22_3 .C_ON=1'b0;
    defparam \c0.data_in_1__1__2284_LC_12_22_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_1__1__2284_LC_12_22_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_in_1__1__2284_LC_12_22_3  (
            .in0(N__39204),
            .in1(N__35370),
            .in2(_gnd_net_),
            .in3(N__35409),
            .lcout(data_in_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49746),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i25_LC_12_22_4 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i25_LC_12_22_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i25_LC_12_22_4 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0__i25_LC_12_22_4  (
            .in0(N__37487),
            .in1(N__36800),
            .in2(N__40624),
            .in3(N__39372),
            .lcout(\c0.data_in_frame_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49746),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i30_LC_12_22_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i30_LC_12_22_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i30_LC_12_22_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \c0.data_in_frame_0__i30_LC_12_22_5  (
            .in0(N__39370),
            .in1(N__40614),
            .in2(N__35345),
            .in3(N__36679),
            .lcout(\c0.data_in_frame_3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49746),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i20_LC_12_22_6 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i20_LC_12_22_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i20_LC_12_22_6 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0__i20_LC_12_22_6  (
            .in0(N__37735),
            .in1(N__35317),
            .in2(N__35298),
            .in3(N__39371),
            .lcout(\c0.data_in_frame_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49746),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_3__3__2266_LC_12_23_0 .C_ON=1'b0;
    defparam \c0.data_in_3__3__2266_LC_12_23_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_3__3__2266_LC_12_23_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.data_in_3__3__2266_LC_12_23_0  (
            .in0(N__35293),
            .in1(N__39142),
            .in2(_gnd_net_),
            .in3(N__35233),
            .lcout(data_in_3_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49758),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i18_4_lut_LC_12_23_1 .C_ON=1'b0;
    defparam \c0.i18_4_lut_LC_12_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i18_4_lut_LC_12_23_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i18_4_lut_LC_12_23_1  (
            .in0(N__43191),
            .in1(N__37285),
            .in2(N__43119),
            .in3(N__35214),
            .lcout(),
            .ltout(\c0.n47_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i27_4_lut_LC_12_23_2 .C_ON=1'b0;
    defparam \c0.i27_4_lut_LC_12_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i27_4_lut_LC_12_23_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i27_4_lut_LC_12_23_2  (
            .in0(N__35178),
            .in1(N__37773),
            .in2(N__35166),
            .in3(N__35163),
            .lcout(),
            .ltout(\c0.n56_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i28_4_lut_LC_12_23_3 .C_ON=1'b0;
    defparam \c0.i28_4_lut_LC_12_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i28_4_lut_LC_12_23_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i28_4_lut_LC_12_23_3  (
            .in0(N__35157),
            .in1(N__40689),
            .in2(N__35145),
            .in3(N__35142),
            .lcout(\c0.n10018 ),
            .ltout(\c0.n10018_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_4_lut_LC_12_23_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_4_lut_LC_12_23_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_4_lut_LC_12_23_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \c0.i1_2_lut_3_lut_4_lut_LC_12_23_4  (
            .in0(N__36071),
            .in1(N__35682),
            .in2(N__35130),
            .in3(N__40193),
            .lcout(FRAME_MATCHER_i_31__N_1272),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_636_LC_12_23_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_636_LC_12_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_636_LC_12_23_5 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_636_LC_12_23_5  (
            .in0(N__40192),
            .in1(N__36070),
            .in2(_gnd_net_),
            .in3(N__35533),
            .lcout(n5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i0_LC_12_23_7 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i0_LC_12_23_7 .SEQ_MODE=4'b1000;
    defparam \c0.FRAME_MATCHER_state_i0_LC_12_23_7 .LUT_INIT=16'b1111101110101010;
    LogicCell40 \c0.FRAME_MATCHER_state_i0_LC_12_23_7  (
            .in0(N__35790),
            .in1(N__35775),
            .in2(N__40220),
            .in3(N__35445),
            .lcout(FRAME_MATCHER_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49758),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx2_transmit_2261_LC_12_24_1 .C_ON=1'b0;
    defparam \c0.tx2_transmit_2261_LC_12_24_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx2_transmit_2261_LC_12_24_1 .LUT_INIT=16'b0011111100100010;
    LogicCell40 \c0.tx2_transmit_2261_LC_12_24_1  (
            .in0(N__35719),
            .in1(N__40219),
            .in2(N__35622),
            .in3(N__36069),
            .lcout(\c0.r_SM_Main_2_N_2034_0_adj_2167 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49771),
            .ce(),
            .sr(N__35553));
    defparam i1_4_lut_adj_796_LC_12_24_4.C_ON=1'b0;
    defparam i1_4_lut_adj_796_LC_12_24_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_796_LC_12_24_4.LUT_INIT=16'b1100110011001000;
    LogicCell40 i1_4_lut_adj_796_LC_12_24_4 (
            .in0(N__35438),
            .in1(N__35499),
            .in2(N__35493),
            .in3(N__35453),
            .lcout(n17063),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_LC_12_24_5.C_ON=1'b0;
    defparam i2_4_lut_LC_12_24_5.SEQ_MODE=4'b0000;
    defparam i2_4_lut_LC_12_24_5.LUT_INIT=16'b1111111011111111;
    LogicCell40 i2_4_lut_LC_12_24_5 (
            .in0(N__35454),
            .in1(N__35439),
            .in2(N__35871),
            .in3(N__35421),
            .lcout(n17090),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_LC_12_24_6.C_ON=1'b0;
    defparam i1_2_lut_LC_12_24_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_LC_12_24_6.LUT_INIT=16'b1010101000000000;
    LogicCell40 i1_2_lut_LC_12_24_6 (
            .in0(N__41967),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42015),
            .lcout(n3_adj_2485),
            .ltout(n3_adj_2485_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_4_lut_adj_795_LC_12_24_7.C_ON=1'b0;
    defparam i3_4_lut_adj_795_LC_12_24_7.SEQ_MODE=4'b0000;
    defparam i3_4_lut_adj_795_LC_12_24_7.LUT_INIT=16'b1111101110101010;
    LogicCell40 i3_4_lut_adj_795_LC_12_24_7 (
            .in0(N__35430),
            .in1(N__35420),
            .in2(N__35412),
            .in3(N__36120),
            .lcout(n8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_689_LC_12_25_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_689_LC_12_25_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_689_LC_12_25_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_689_LC_12_25_0  (
            .in0(N__48713),
            .in1(N__42143),
            .in2(_gnd_net_),
            .in3(N__48815),
            .lcout(\c0.n10188 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i14651_4_lut_LC_12_25_1.C_ON=1'b0;
    defparam i14651_4_lut_LC_12_25_1.SEQ_MODE=4'b0000;
    defparam i14651_4_lut_LC_12_25_1.LUT_INIT=16'b1111111010001100;
    LogicCell40 i14651_4_lut_LC_12_25_1 (
            .in0(N__36279),
            .in1(N__36246),
            .in2(N__36210),
            .in3(N__36170),
            .lcout(n17428),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.select_217_Select_2_i4_3_lut_LC_12_25_2 .C_ON=1'b0;
    defparam \c0.select_217_Select_2_i4_3_lut_LC_12_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.select_217_Select_2_i4_3_lut_LC_12_25_2 .LUT_INIT=16'b1111101000000000;
    LogicCell40 \c0.select_217_Select_2_i4_3_lut_LC_12_25_2  (
            .in0(N__36118),
            .in1(_gnd_net_),
            .in2(N__35957),
            .in3(N__35903),
            .lcout(),
            .ltout(n4_adj_2417_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i2_LC_12_25_3 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i2_LC_12_25_3 .SEQ_MODE=4'b1000;
    defparam \c0.FRAME_MATCHER_state_i2_LC_12_25_3 .LUT_INIT=16'b1111110111111100;
    LogicCell40 \c0.FRAME_MATCHER_state_i2_LC_12_25_3  (
            .in0(N__36138),
            .in1(N__36129),
            .in2(N__36123),
            .in3(N__36119),
            .lcout(FRAME_MATCHER_state_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49783),
            .ce(),
            .sr(_gnd_net_));
    defparam i14652_3_lut_LC_12_25_4.C_ON=1'b0;
    defparam i14652_3_lut_LC_12_25_4.SEQ_MODE=4'b0000;
    defparam i14652_3_lut_LC_12_25_4.LUT_INIT=16'b0010001001110111;
    LogicCell40 i14652_3_lut_LC_12_25_4 (
            .in0(N__36015),
            .in1(N__35994),
            .in2(_gnd_net_),
            .in3(N__35988),
            .lcout(LED_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_792_LC_12_25_5.C_ON=1'b0;
    defparam i1_2_lut_adj_792_LC_12_25_5.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_792_LC_12_25_5.LUT_INIT=16'b0011001100000000;
    LogicCell40 i1_2_lut_adj_792_LC_12_25_5 (
            .in0(_gnd_net_),
            .in1(N__35950),
            .in2(_gnd_net_),
            .in3(N__35902),
            .lcout(n6_adj_2488),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i2_3_lut_LC_12_25_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i2_3_lut_LC_12_25_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_0_i2_3_lut_LC_12_25_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_0_i2_3_lut_LC_12_25_7  (
            .in0(N__37994),
            .in1(N__35862),
            .in2(_gnd_net_),
            .in3(N__47787),
            .lcout(n2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_460_LC_12_26_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_460_LC_12_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_460_LC_12_26_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_460_LC_12_26_0  (
            .in0(_gnd_net_),
            .in1(N__43469),
            .in2(_gnd_net_),
            .in3(N__44285),
            .lcout(\c0.n17264 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_4_lut_adj_782_LC_12_26_2.C_ON=1'b0;
    defparam i24_4_lut_adj_782_LC_12_26_2.SEQ_MODE=4'b0000;
    defparam i24_4_lut_adj_782_LC_12_26_2.LUT_INIT=16'b0010001011100010;
    LogicCell40 i24_4_lut_adj_782_LC_12_26_2 (
            .in0(N__35844),
            .in1(N__46375),
            .in2(N__42207),
            .in3(N__46290),
            .lcout(),
            .ltout(n10_adj_2409_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i3_LC_12_26_3 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i3_LC_12_26_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i3_LC_12_26_3 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \c0.tx.r_Tx_Data_i3_LC_12_26_3  (
            .in0(N__43814),
            .in1(N__44105),
            .in2(N__36357),
            .in3(N__36392),
            .lcout(r_Tx_Data_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49793),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_2_i8_3_lut_LC_12_26_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_2_i8_3_lut_LC_12_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_2_i8_3_lut_LC_12_26_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_2_i8_3_lut_LC_12_26_5  (
            .in0(N__49169),
            .in1(N__48717),
            .in2(_gnd_net_),
            .in3(N__47794),
            .lcout(),
            .ltout(\c0.n8_adj_2183_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_2_i10_4_lut_LC_12_26_6 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_2_i10_4_lut_LC_12_26_6 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_2_i10_4_lut_LC_12_26_6 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_2_i10_4_lut_LC_12_26_6  (
            .in0(N__47795),
            .in1(N__45465),
            .in2(N__36354),
            .in3(N__47458),
            .lcout(n10_adj_2450),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i4_LC_12_26_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i4_LC_12_26_7 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i4_LC_12_26_7 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \c0.byte_transmit_counter__i4_LC_12_26_7  (
            .in0(N__43813),
            .in1(N__42993),
            .in2(N__42452),
            .in3(N__42366),
            .lcout(byte_transmit_counter_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49793),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15366_LC_12_27_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15366_LC_12_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15366_LC_12_27_0 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter_1__bdd_4_lut_15366_LC_12_27_0  (
            .in0(N__36351),
            .in1(N__46289),
            .in2(N__38274),
            .in3(N__47431),
            .lcout(\c0.n18166 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15212_2_lut_3_lut_LC_12_27_1 .C_ON=1'b0;
    defparam \c0.i15212_2_lut_3_lut_LC_12_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.i15212_2_lut_3_lut_LC_12_27_1 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \c0.i15212_2_lut_3_lut_LC_12_27_1  (
            .in0(N__48276),
            .in1(N__48114),
            .in2(_gnd_net_),
            .in3(N__50135),
            .lcout(data_out_10__7__N_110),
            .ltout(data_out_10__7__N_110_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_8__4__2188_LC_12_27_2 .C_ON=1'b0;
    defparam \c0.data_out_8__4__2188_LC_12_27_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_8__4__2188_LC_12_27_2 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_out_8__4__2188_LC_12_27_2  (
            .in0(N__36345),
            .in1(_gnd_net_),
            .in2(N__36321),
            .in3(N__48472),
            .lcout(data_out_8_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49803),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.UART_TRANSMITTER_state__i2_LC_12_27_4 .C_ON=1'b0;
    defparam \c0.UART_TRANSMITTER_state__i2_LC_12_27_4 .SEQ_MODE=4'b1000;
    defparam \c0.UART_TRANSMITTER_state__i2_LC_12_27_4 .LUT_INIT=16'b1001101011010010;
    LogicCell40 \c0.UART_TRANSMITTER_state__i2_LC_12_27_4  (
            .in0(N__50136),
            .in1(N__48278),
            .in2(N__48155),
            .in3(N__38343),
            .lcout(UART_TRANSMITTER_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49803),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_8__6__2186_LC_12_27_5 .C_ON=1'b0;
    defparam \c0.data_out_8__6__2186_LC_12_27_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_8__6__2186_LC_12_27_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_8__6__2186_LC_12_27_5  (
            .in0(N__49929),
            .in1(N__36318),
            .in2(_gnd_net_),
            .in3(N__43386),
            .lcout(data_out_8_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49803),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_1__2__2246_LC_12_27_6 .C_ON=1'b0;
    defparam \c0.data_out_1__2__2246_LC_12_27_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_1__2__2246_LC_12_27_6 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \c0.data_out_1__2__2246_LC_12_27_6  (
            .in0(N__50137),
            .in1(N__48277),
            .in2(N__50587),
            .in3(N__36293),
            .lcout(\c0.data_out_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49803),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15075_2_lut_LC_12_27_7 .C_ON=1'b0;
    defparam \c0.i15075_2_lut_LC_12_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.i15075_2_lut_LC_12_27_7 .LUT_INIT=16'b1110111011101110;
    LogicCell40 \c0.i15075_2_lut_LC_12_27_7  (
            .in0(N__47802),
            .in1(N__42768),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.n17696 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n18070_bdd_4_lut_LC_12_28_0.C_ON=1'b0;
    defparam n18070_bdd_4_lut_LC_12_28_0.SEQ_MODE=4'b0000;
    defparam n18070_bdd_4_lut_LC_12_28_0.LUT_INIT=16'b1110111001010000;
    LogicCell40 n18070_bdd_4_lut_LC_12_28_0 (
            .in0(N__42626),
            .in1(N__38694),
            .in2(N__36426),
            .in3(N__36378),
            .lcout(),
            .ltout(n18073_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i33_3_lut_LC_12_28_1 .C_ON=1'b0;
    defparam \c0.tx.i33_3_lut_LC_12_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i33_3_lut_LC_12_28_1 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \c0.tx.i33_3_lut_LC_12_28_1  (
            .in0(_gnd_net_),
            .in1(N__42578),
            .in2(N__36432),
            .in3(N__38232),
            .lcout(\c0.tx.n31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_4_lut_LC_12_28_2 .C_ON=1'b0;
    defparam \c0.tx.i1_4_lut_LC_12_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_4_lut_LC_12_28_2 .LUT_INIT=16'b0001000100000001;
    LogicCell40 \c0.tx.i1_4_lut_LC_12_28_2  (
            .in0(N__45927),
            .in1(N__44014),
            .in2(N__44212),
            .in3(N__43950),
            .lcout(\c0.tx.n10688 ),
            .ltout(\c0.tx.n10688_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_i0_LC_12_28_3 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_i0_LC_12_28_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Bit_Index_i0_LC_12_28_3 .LUT_INIT=16'b0000111111000000;
    LogicCell40 \c0.tx.r_Bit_Index_i0_LC_12_28_3  (
            .in0(_gnd_net_),
            .in1(N__44203),
            .in2(N__36429),
            .in3(N__42579),
            .lcout(\c0.tx.r_Bit_Index_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49810),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i1_LC_12_28_4 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i1_LC_12_28_4 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i1_LC_12_28_4 .LUT_INIT=16'b0000110010101010;
    LogicCell40 \c0.tx.r_Tx_Data_i1_LC_12_28_4  (
            .in0(N__36425),
            .in1(N__42231),
            .in2(N__43842),
            .in3(N__44099),
            .lcout(r_Tx_Data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49810),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_8__1__2191_LC_12_28_5 .C_ON=1'b0;
    defparam \c0.data_out_8__1__2191_LC_12_28_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_8__1__2191_LC_12_28_5 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \c0.data_out_8__1__2191_LC_12_28_5  (
            .in0(N__36414),
            .in1(_gnd_net_),
            .in2(N__49963),
            .in3(N__42136),
            .lcout(data_out_8_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49810),
            .ce(),
            .sr(_gnd_net_));
    defparam r_Bit_Index_2__bdd_4_lut_15385_LC_12_28_6.C_ON=1'b0;
    defparam r_Bit_Index_2__bdd_4_lut_15385_LC_12_28_6.SEQ_MODE=4'b0000;
    defparam r_Bit_Index_2__bdd_4_lut_15385_LC_12_28_6.LUT_INIT=16'b1111010110001000;
    LogicCell40 r_Bit_Index_2__bdd_4_lut_15385_LC_12_28_6 (
            .in0(N__42625),
            .in1(N__36393),
            .in2(N__43608),
            .in3(N__42546),
            .lcout(n18070),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Bit_Index_i1_LC_12_28_7 .C_ON=1'b0;
    defparam \c0.tx.r_Bit_Index_i1_LC_12_28_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Bit_Index_i1_LC_12_28_7 .LUT_INIT=16'b0100100011110000;
    LogicCell40 \c0.tx.r_Bit_Index_i1_LC_12_28_7  (
            .in0(N__42584),
            .in1(N__44204),
            .in2(N__42641),
            .in3(N__36372),
            .lcout(r_Bit_Index_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49810),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i0_LC_12_29_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i0_LC_12_29_0 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i0_LC_12_29_0 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \c0.byte_transmit_counter__i0_LC_12_29_0  (
            .in0(N__47677),
            .in1(N__42894),
            .in2(N__42461),
            .in3(N__42350),
            .lcout(byte_transmit_counter_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49818),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_607_LC_12_29_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_607_LC_12_29_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_607_LC_12_29_1 .LUT_INIT=16'b0000111000001111;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_607_LC_12_29_1  (
            .in0(N__50719),
            .in1(N__38664),
            .in2(N__48099),
            .in3(N__38558),
            .lcout(n4_adj_2419),
            .ltout(n4_adj_2419_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_2_lut_LC_12_29_2.C_ON=1'b0;
    defparam i2_2_lut_LC_12_29_2.SEQ_MODE=4'b0000;
    defparam i2_2_lut_LC_12_29_2.LUT_INIT=16'b1010000010100000;
    LogicCell40 i2_2_lut_LC_12_29_2 (
            .in0(N__50205),
            .in1(_gnd_net_),
            .in2(N__36465),
            .in3(_gnd_net_),
            .lcout(n5_adj_2407),
            .ltout(n5_adj_2407_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_4_lut_adj_788_LC_12_29_3.C_ON=1'b0;
    defparam i24_4_lut_adj_788_LC_12_29_3.SEQ_MODE=4'b0000;
    defparam i24_4_lut_adj_788_LC_12_29_3.LUT_INIT=16'b0111010000110000;
    LogicCell40 i24_4_lut_adj_788_LC_12_29_3 (
            .in0(N__48020),
            .in1(N__48298),
            .in2(N__36462),
            .in3(N__38214),
            .lcout(n10_adj_2444),
            .ltout(n10_adj_2444_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i2_LC_12_29_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i2_LC_12_29_4 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i2_LC_12_29_4 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \c0.byte_transmit_counter__i2_LC_12_29_4  (
            .in0(N__42456),
            .in1(N__42852),
            .in2(N__36459),
            .in3(N__46255),
            .lcout(byte_transmit_counter_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49818),
            .ce(),
            .sr(_gnd_net_));
    defparam i52_4_lut_LC_12_29_5.C_ON=1'b0;
    defparam i52_4_lut_LC_12_29_5.SEQ_MODE=4'b0000;
    defparam i52_4_lut_LC_12_29_5.LUT_INIT=16'b0010001011100010;
    LogicCell40 i52_4_lut_LC_12_29_5 (
            .in0(N__36456),
            .in1(N__47497),
            .in2(N__48759),
            .in3(N__47676),
            .lcout(n25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15147_4_lut_LC_12_29_6.C_ON=1'b0;
    defparam i15147_4_lut_LC_12_29_6.SEQ_MODE=4'b0000;
    defparam i15147_4_lut_LC_12_29_6.LUT_INIT=16'b1111100010101000;
    LogicCell40 i15147_4_lut_LC_12_29_6 (
            .in0(N__50206),
            .in1(N__36450),
            .in2(N__48371),
            .in3(N__38340),
            .lcout(n17765),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_i2_LC_12_30_1 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_i2_LC_12_30_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_SM_Main_i2_LC_12_30_1 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \c0.tx.r_SM_Main_i2_LC_12_30_1  (
            .in0(N__44016),
            .in1(N__45894),
            .in2(N__44213),
            .in3(N__43956),
            .lcout(\c0.tx.r_SM_Main_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49825),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10536_2_lut_3_lut_4_lut_LC_12_30_2 .C_ON=1'b0;
    defparam \c0.i10536_2_lut_3_lut_4_lut_LC_12_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.i10536_2_lut_3_lut_4_lut_LC_12_30_2 .LUT_INIT=16'b1100110011000100;
    LogicCell40 \c0.i10536_2_lut_3_lut_4_lut_LC_12_30_2  (
            .in0(N__38564),
            .in1(N__38745),
            .in2(N__50742),
            .in3(N__38647),
            .lcout(\c0.n22_adj_2313 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10543_2_lut_3_lut_4_lut_LC_12_30_3 .C_ON=1'b0;
    defparam \c0.i10543_2_lut_3_lut_4_lut_LC_12_30_3 .SEQ_MODE=4'b0000;
    defparam \c0.i10543_2_lut_3_lut_4_lut_LC_12_30_3 .LUT_INIT=16'b1110000011110000;
    LogicCell40 \c0.i10543_2_lut_3_lut_4_lut_LC_12_30_3  (
            .in0(N__50718),
            .in1(N__38638),
            .in2(N__38415),
            .in3(N__38562),
            .lcout(\c0.n27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10539_2_lut_3_lut_4_lut_LC_12_30_4 .C_ON=1'b0;
    defparam \c0.i10539_2_lut_3_lut_4_lut_LC_12_30_4 .SEQ_MODE=4'b0000;
    defparam \c0.i10539_2_lut_3_lut_4_lut_LC_12_30_4 .LUT_INIT=16'b1100110011000100;
    LogicCell40 \c0.i10539_2_lut_3_lut_4_lut_LC_12_30_4  (
            .in0(N__38563),
            .in1(N__38493),
            .in2(N__50741),
            .in3(N__38646),
            .lcout(\c0.n25_adj_2386 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i5_3_lut_LC_12_30_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i5_3_lut_LC_12_30_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i5_3_lut_LC_12_30_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_5_i5_3_lut_LC_12_30_5  (
            .in0(N__43629),
            .in1(N__47653),
            .in2(_gnd_net_),
            .in3(N__48864),
            .lcout(\c0.n5_adj_2163 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10535_2_lut_3_lut_4_lut_LC_12_30_6 .C_ON=1'b0;
    defparam \c0.i10535_2_lut_3_lut_4_lut_LC_12_30_6 .SEQ_MODE=4'b0000;
    defparam \c0.i10535_2_lut_3_lut_4_lut_LC_12_30_6 .LUT_INIT=16'b1100110011000100;
    LogicCell40 \c0.i10535_2_lut_3_lut_4_lut_LC_12_30_6  (
            .in0(N__38565),
            .in1(N__38454),
            .in2(N__50743),
            .in3(N__38648),
            .lcout(\c0.n21_adj_2262 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_2361__i0_LC_12_31_0 .C_ON=1'b1;
    defparam \c0.delay_counter_2361__i0_LC_12_31_0 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_2361__i0_LC_12_31_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_2361__i0_LC_12_31_0  (
            .in0(_gnd_net_),
            .in1(N__38304),
            .in2(N__38289),
            .in3(_gnd_net_),
            .lcout(\c0.delay_counter_0 ),
            .ltout(),
            .carryin(bfn_12_31_0_),
            .carryout(\c0.n16066 ),
            .clk(N__49831),
            .ce(N__36551),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_2361__i1_LC_12_31_1 .C_ON=1'b1;
    defparam \c0.delay_counter_2361__i1_LC_12_31_1 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_2361__i1_LC_12_31_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_2361__i1_LC_12_31_1  (
            .in0(_gnd_net_),
            .in1(N__36495),
            .in2(_gnd_net_),
            .in3(N__36489),
            .lcout(\c0.delay_counter_1 ),
            .ltout(),
            .carryin(\c0.n16066 ),
            .carryout(\c0.n16067 ),
            .clk(N__49831),
            .ce(N__36551),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_2361__i2_LC_12_31_2 .C_ON=1'b1;
    defparam \c0.delay_counter_2361__i2_LC_12_31_2 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_2361__i2_LC_12_31_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_2361__i2_LC_12_31_2  (
            .in0(_gnd_net_),
            .in1(N__38763),
            .in2(_gnd_net_),
            .in3(N__36486),
            .lcout(\c0.delay_counter_2 ),
            .ltout(),
            .carryin(\c0.n16067 ),
            .carryout(\c0.n16068 ),
            .clk(N__49831),
            .ce(N__36551),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_2361__i3_LC_12_31_3 .C_ON=1'b1;
    defparam \c0.delay_counter_2361__i3_LC_12_31_3 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_2361__i3_LC_12_31_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_2361__i3_LC_12_31_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__36483),
            .in3(N__36474),
            .lcout(\c0.delay_counter_3 ),
            .ltout(),
            .carryin(\c0.n16068 ),
            .carryout(\c0.n16069 ),
            .clk(N__49831),
            .ce(N__36551),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_2361__i4_LC_12_31_4 .C_ON=1'b1;
    defparam \c0.delay_counter_2361__i4_LC_12_31_4 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_2361__i4_LC_12_31_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_2361__i4_LC_12_31_4  (
            .in0(_gnd_net_),
            .in1(N__38355),
            .in2(_gnd_net_),
            .in3(N__36471),
            .lcout(\c0.delay_counter_4 ),
            .ltout(),
            .carryin(\c0.n16069 ),
            .carryout(\c0.n16070 ),
            .clk(N__49831),
            .ce(N__36551),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_2361__i5_LC_12_31_5 .C_ON=1'b1;
    defparam \c0.delay_counter_2361__i5_LC_12_31_5 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_2361__i5_LC_12_31_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_2361__i5_LC_12_31_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38298),
            .in3(N__36468),
            .lcout(\c0.delay_counter_5 ),
            .ltout(),
            .carryin(\c0.n16070 ),
            .carryout(\c0.n16071 ),
            .clk(N__49831),
            .ce(N__36551),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_2361__i6_LC_12_31_6 .C_ON=1'b1;
    defparam \c0.delay_counter_2361__i6_LC_12_31_6 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_2361__i6_LC_12_31_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_2361__i6_LC_12_31_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__36591),
            .in3(N__36582),
            .lcout(\c0.delay_counter_6 ),
            .ltout(),
            .carryin(\c0.n16071 ),
            .carryout(\c0.n16072 ),
            .clk(N__49831),
            .ce(N__36551),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_2361__i7_LC_12_31_7 .C_ON=1'b1;
    defparam \c0.delay_counter_2361__i7_LC_12_31_7 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_2361__i7_LC_12_31_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_2361__i7_LC_12_31_7  (
            .in0(_gnd_net_),
            .in1(N__36579),
            .in2(_gnd_net_),
            .in3(N__36573),
            .lcout(\c0.delay_counter_7 ),
            .ltout(),
            .carryin(\c0.n16072 ),
            .carryout(\c0.n16073 ),
            .clk(N__49831),
            .ce(N__36551),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_2361__i8_LC_12_32_0 .C_ON=1'b1;
    defparam \c0.delay_counter_2361__i8_LC_12_32_0 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_2361__i8_LC_12_32_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_2361__i8_LC_12_32_0  (
            .in0(_gnd_net_),
            .in1(N__38460),
            .in2(_gnd_net_),
            .in3(N__36570),
            .lcout(\c0.delay_counter_8 ),
            .ltout(),
            .carryin(bfn_12_32_0_),
            .carryout(\c0.n16074 ),
            .clk(N__49836),
            .ce(N__36552),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_2361__i9_LC_12_32_1 .C_ON=1'b1;
    defparam \c0.delay_counter_2361__i9_LC_12_32_1 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_2361__i9_LC_12_32_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_2361__i9_LC_12_32_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38322),
            .in3(N__36567),
            .lcout(\c0.delay_counter_9 ),
            .ltout(),
            .carryin(\c0.n16074 ),
            .carryout(\c0.n16075 ),
            .clk(N__49836),
            .ce(N__36552),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_2361__i10_LC_12_32_2 .C_ON=1'b1;
    defparam \c0.delay_counter_2361__i10_LC_12_32_2 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_2361__i10_LC_12_32_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_2361__i10_LC_12_32_2  (
            .in0(_gnd_net_),
            .in1(N__38718),
            .in2(_gnd_net_),
            .in3(N__36564),
            .lcout(\c0.delay_counter_10 ),
            .ltout(),
            .carryin(\c0.n16075 ),
            .carryout(\c0.n16076 ),
            .clk(N__49836),
            .ce(N__36552),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_2361__i11_LC_12_32_3 .C_ON=1'b1;
    defparam \c0.delay_counter_2361__i11_LC_12_32_3 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_2361__i11_LC_12_32_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_2361__i11_LC_12_32_3  (
            .in0(_gnd_net_),
            .in1(N__38511),
            .in2(_gnd_net_),
            .in3(N__36561),
            .lcout(\c0.delay_counter_11 ),
            .ltout(),
            .carryin(\c0.n16076 ),
            .carryout(\c0.n16077 ),
            .clk(N__49836),
            .ce(N__36552),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_2361__i12_LC_12_32_4 .C_ON=1'b1;
    defparam \c0.delay_counter_2361__i12_LC_12_32_4 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_2361__i12_LC_12_32_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_2361__i12_LC_12_32_4  (
            .in0(_gnd_net_),
            .in1(N__38778),
            .in2(_gnd_net_),
            .in3(N__36558),
            .lcout(\c0.delay_counter_12 ),
            .ltout(),
            .carryin(\c0.n16077 ),
            .carryout(\c0.n16078 ),
            .clk(N__49836),
            .ce(N__36552),
            .sr(_gnd_net_));
    defparam \c0.delay_counter_2361__i13_LC_12_32_5 .C_ON=1'b0;
    defparam \c0.delay_counter_2361__i13_LC_12_32_5 .SEQ_MODE=4'b1000;
    defparam \c0.delay_counter_2361__i13_LC_12_32_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.delay_counter_2361__i13_LC_12_32_5  (
            .in0(_gnd_net_),
            .in1(N__38700),
            .in2(_gnd_net_),
            .in3(N__36555),
            .lcout(\c0.delay_counter_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49836),
            .ce(N__36552),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_678_LC_13_18_0 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_678_LC_13_18_0 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_678_LC_13_18_0 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \c0.i13_4_lut_adj_678_LC_13_18_0  (
            .in0(N__36528),
            .in1(N__36522),
            .in2(N__36513),
            .in3(N__36501),
            .lcout(\c0.n29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i0_LC_13_18_1 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i0_LC_13_18_1 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i0_LC_13_18_1 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.rx.r_Rx_Byte_i0_LC_13_18_1  (
            .in0(N__37961),
            .in1(N__45216),
            .in2(N__36778),
            .in3(N__45175),
            .lcout(rx_data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49716),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i1_LC_13_18_2 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i1_LC_13_18_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i1_LC_13_18_2 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \c0.data_out_frame2_0___i1_LC_13_18_2  (
            .in0(N__39936),
            .in1(N__39875),
            .in2(N__39846),
            .in3(N__40632),
            .lcout(\c0.data_out_frame2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49716),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Data_50_LC_13_18_3 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Data_50_LC_13_18_3 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Data_50_LC_13_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.rx.r_Rx_Data_50_LC_13_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36738),
            .lcout(r_Rx_Data),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49716),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_561_LC_13_18_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_561_LC_13_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_561_LC_13_18_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i1_2_lut_adj_561_LC_13_18_4  (
            .in0(N__41946),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40243),
            .lcout(\c0.n26_adj_2174 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i7_LC_13_18_5 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i7_LC_13_18_5 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i7_LC_13_18_5 .LUT_INIT=16'b1111010010110000;
    LogicCell40 \c0.rx.r_Rx_Byte_i7_LC_13_18_5  (
            .in0(N__36720),
            .in1(N__39572),
            .in2(N__40501),
            .in3(N__45219),
            .lcout(rx_data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49716),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i1_LC_13_18_6 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i1_LC_13_18_6 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i1_LC_13_18_6 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.rx.r_Rx_Byte_i1_LC_13_18_6  (
            .in0(N__45217),
            .in1(N__37962),
            .in2(N__39446),
            .in3(N__36718),
            .lcout(rx_data_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49716),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i5_LC_13_18_7 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i5_LC_13_18_7 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i5_LC_13_18_7 .LUT_INIT=16'b1100110111001000;
    LogicCell40 \c0.rx.r_Rx_Byte_i5_LC_13_18_7  (
            .in0(N__36719),
            .in1(N__36655),
            .in2(N__45294),
            .in3(N__45218),
            .lcout(rx_data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49716),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_603_LC_13_19_0 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_603_LC_13_19_0 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_603_LC_13_19_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i13_4_lut_adj_603_LC_13_19_0  (
            .in0(N__36618),
            .in1(N__37341),
            .in2(N__36609),
            .in3(N__36597),
            .lcout(\c0.n4494 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15063_3_lut_4_lut_LC_13_19_1 .C_ON=1'b0;
    defparam \c0.i15063_3_lut_4_lut_LC_13_19_1 .SEQ_MODE=4'b0000;
    defparam \c0.i15063_3_lut_4_lut_LC_13_19_1 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \c0.i15063_3_lut_4_lut_LC_13_19_1  (
            .in0(N__37568),
            .in1(N__41957),
            .in2(N__40146),
            .in3(N__40246),
            .lcout(\c0.n17688 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_413_LC_13_19_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_413_LC_13_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_413_LC_13_19_2 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \c0.i1_2_lut_adj_413_LC_13_19_2  (
            .in0(_gnd_net_),
            .in1(N__37191),
            .in2(_gnd_net_),
            .in3(N__37112),
            .lcout(\c0.n15171 ),
            .ltout(\c0.n15171_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i15_LC_13_19_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i15_LC_13_19_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i15_LC_13_19_3 .LUT_INIT=16'b1010101010101100;
    LogicCell40 \c0.data_in_frame_0__i15_LC_13_19_3  (
            .in0(N__37046),
            .in1(N__39519),
            .in2(N__37050),
            .in3(N__40430),
            .lcout(\c0.data_in_frame_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49726),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11_4_lut_adj_676_LC_13_19_5 .C_ON=1'b0;
    defparam \c0.i11_4_lut_adj_676_LC_13_19_5 .SEQ_MODE=4'b0000;
    defparam \c0.i11_4_lut_adj_676_LC_13_19_5 .LUT_INIT=16'b1011111011111111;
    LogicCell40 \c0.i11_4_lut_adj_676_LC_13_19_5  (
            .in0(N__38796),
            .in1(N__37017),
            .in2(N__36999),
            .in3(N__36978),
            .lcout(),
            .ltout(\c0.n27_adj_2381_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_702_LC_13_19_6 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_702_LC_13_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_702_LC_13_19_6 .LUT_INIT=16'b0101010101010100;
    LogicCell40 \c0.i1_4_lut_adj_702_LC_13_19_6  (
            .in0(N__40244),
            .in1(N__36972),
            .in2(N__36966),
            .in3(N__36963),
            .lcout(\c0.n12491 ),
            .ltout(\c0.n12491_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15059_3_lut_4_lut_LC_13_19_7 .C_ON=1'b0;
    defparam \c0.i15059_3_lut_4_lut_LC_13_19_7 .SEQ_MODE=4'b0000;
    defparam \c0.i15059_3_lut_4_lut_LC_13_19_7 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \c0.i15059_3_lut_4_lut_LC_13_19_7  (
            .in0(N__37622),
            .in1(N__41956),
            .in2(N__36957),
            .in3(N__40245),
            .lcout(\c0.n17686 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_458_LC_13_20_0 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_458_LC_13_20_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_458_LC_13_20_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_458_LC_13_20_0  (
            .in0(_gnd_net_),
            .in1(N__41031),
            .in2(_gnd_net_),
            .in3(N__36948),
            .lcout(\c0.n10259 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i18_LC_13_20_1 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i18_LC_13_20_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i18_LC_13_20_1 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \c0.data_in_frame_0__i18_LC_13_20_1  (
            .in0(N__37439),
            .in1(N__37740),
            .in2(N__39480),
            .in3(N__39388),
            .lcout(\c0.data_in_frame_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49736),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i24_LC_13_20_2 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i24_LC_13_20_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i24_LC_13_20_2 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \c0.data_in_frame_0__i24_LC_13_20_2  (
            .in0(N__39387),
            .in1(N__40500),
            .in2(N__37746),
            .in3(N__36902),
            .lcout(\c0.data_in_frame_2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49736),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i19_LC_13_20_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i19_LC_13_20_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i19_LC_13_20_3 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \c0.data_in_frame_0__i19_LC_13_20_3  (
            .in0(N__36840),
            .in1(N__37741),
            .in2(N__37422),
            .in3(N__39389),
            .lcout(\c0.data_in_frame_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49736),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i5_LC_13_20_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i5_LC_13_20_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i5_LC_13_20_4 .LUT_INIT=16'b1111000010101100;
    LogicCell40 \c0.data_out_frame2_0___i5_LC_13_20_4  (
            .in0(N__37644),
            .in1(N__37623),
            .in2(N__39729),
            .in3(N__39946),
            .lcout(\c0.data_out_frame2_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49736),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i4_LC_13_20_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i4_LC_13_20_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i4_LC_13_20_5 .LUT_INIT=16'b1101110010011000;
    LogicCell40 \c0.data_out_frame2_0___i4_LC_13_20_5  (
            .in0(N__39945),
            .in1(N__39725),
            .in2(N__37583),
            .in3(N__37593),
            .lcout(\c0.data_out_frame2_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49736),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_587_LC_13_20_6 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_587_LC_13_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_587_LC_13_20_6 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \c0.i4_4_lut_adj_587_LC_13_20_6  (
            .in0(N__37524),
            .in1(N__37503),
            .in2(N__37491),
            .in3(N__37473),
            .lcout(),
            .ltout(\c0.n18_adj_2316_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9_4_lut_adj_600_LC_13_20_7 .C_ON=1'b0;
    defparam \c0.i9_4_lut_adj_600_LC_13_20_7 .SEQ_MODE=4'b0000;
    defparam \c0.i9_4_lut_adj_600_LC_13_20_7 .LUT_INIT=16'b1111011111111011;
    LogicCell40 \c0.i9_4_lut_adj_600_LC_13_20_7  (
            .in0(N__37438),
            .in1(N__37418),
            .in2(N__37401),
            .in3(N__37389),
            .lcout(\c0.n23_adj_2322 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i23_LC_13_21_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i23_LC_13_21_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i23_LC_13_21_0 .LUT_INIT=16'b1110000011000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i23_LC_13_21_0  (
            .in0(N__44982),
            .in1(N__44714),
            .in2(N__37334),
            .in3(N__44566),
            .lcout(\c0.FRAME_MATCHER_state_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49747),
            .ce(),
            .sr(N__37308));
    defparam \c0.FRAME_MATCHER_state_i11_LC_13_22_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i11_LC_13_22_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i11_LC_13_22_0 .LUT_INIT=16'b1110000011000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i11_LC_13_22_0  (
            .in0(N__44915),
            .in1(N__44676),
            .in2(N__37295),
            .in3(N__44512),
            .lcout(\c0.FRAME_MATCHER_state_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49759),
            .ce(),
            .sr(N__37269));
    defparam \c0.i1_2_lut_adj_754_LC_13_22_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_754_LC_13_22_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_754_LC_13_22_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_754_LC_13_22_1  (
            .in0(_gnd_net_),
            .in1(N__41227),
            .in2(_gnd_net_),
            .in3(N__40718),
            .lcout(\c0.n16658 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_2_lut_LC_13_22_2 .C_ON=1'b0;
    defparam \c0.i3_2_lut_LC_13_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_2_lut_LC_13_22_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i3_2_lut_LC_13_22_2  (
            .in0(_gnd_net_),
            .in1(N__37253),
            .in2(_gnd_net_),
            .in3(N__39263),
            .lcout(\c0.n16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.equal_52_i4_2_lut_LC_13_22_3 .C_ON=1'b0;
    defparam \c0.rx.equal_52_i4_2_lut_LC_13_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.rx.equal_52_i4_2_lut_LC_13_22_3 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \c0.rx.equal_52_i4_2_lut_LC_13_22_3  (
            .in0(N__37917),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37947),
            .lcout(n4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.equal_55_i4_2_lut_LC_13_22_4 .C_ON=1'b0;
    defparam \c0.rx.equal_55_i4_2_lut_LC_13_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.rx.equal_55_i4_2_lut_LC_13_22_4 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \c0.rx.equal_55_i4_2_lut_LC_13_22_4  (
            .in0(N__37948),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37918),
            .lcout(n4_adj_2427),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.equal_56_i4_2_lut_LC_13_22_5 .C_ON=1'b0;
    defparam \c0.rx.equal_56_i4_2_lut_LC_13_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.rx.equal_56_i4_2_lut_LC_13_22_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \c0.rx.equal_56_i4_2_lut_LC_13_22_5  (
            .in0(N__37919),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37949),
            .lcout(n4_adj_2416),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i10445_2_lut_LC_13_22_6 .C_ON=1'b0;
    defparam \c0.rx.i10445_2_lut_LC_13_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i10445_2_lut_LC_13_22_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.rx.i10445_2_lut_LC_13_22_6  (
            .in0(N__37950),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37920),
            .lcout(n13116),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.i1_2_lut_adj_397_LC_13_22_7 .C_ON=1'b0;
    defparam \c0.rx.i1_2_lut_adj_397_LC_13_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.rx.i1_2_lut_adj_397_LC_13_22_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \c0.rx.i1_2_lut_adj_397_LC_13_22_7  (
            .in0(N__37875),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37836),
            .lcout(n9999),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i19_4_lut_LC_13_23_0 .C_ON=1'b0;
    defparam \c0.i19_4_lut_LC_13_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i19_4_lut_LC_13_23_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i19_4_lut_LC_13_23_0  (
            .in0(N__43158),
            .in1(N__37808),
            .in2(N__41192),
            .in3(N__37765),
            .lcout(\c0.n48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i30_LC_13_23_1 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i30_LC_13_23_1 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i30_LC_13_23_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i30_LC_13_23_1  (
            .in0(N__37767),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41545),
            .lcout(\c0.FRAME_MATCHER_state_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49772),
            .ce(),
            .sr(N__37755));
    defparam \c0.i1_2_lut_4_lut_adj_767_LC_13_23_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_767_LC_13_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_767_LC_13_23_2 .LUT_INIT=16'b1011101000000000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_767_LC_13_23_2  (
            .in0(N__41322),
            .in1(N__41400),
            .in2(N__41492),
            .in3(N__37766),
            .lcout(\c0.n16698 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_737_LC_13_23_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_737_LC_13_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_737_LC_13_23_3 .LUT_INIT=16'b1010101000001000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_737_LC_13_23_3  (
            .in0(N__41188),
            .in1(N__41473),
            .in2(N__41417),
            .in3(N__41318),
            .lcout(\c0.n16710 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_746_LC_13_23_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_746_LC_13_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_746_LC_13_23_5 .LUT_INIT=16'b1010101000001000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_746_LC_13_23_5  (
            .in0(N__41263),
            .in1(N__41474),
            .in2(N__41418),
            .in3(N__41319),
            .lcout(\c0.n16704 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_759_LC_13_23_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_759_LC_13_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_759_LC_13_23_6 .LUT_INIT=16'b1011101000000000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_759_LC_13_23_6  (
            .in0(N__41320),
            .in1(N__41396),
            .in2(N__41491),
            .in3(N__43118),
            .lcout(\c0.n16688 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_764_LC_13_23_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_764_LC_13_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_764_LC_13_23_7 .LUT_INIT=16'b1010101000001000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_764_LC_13_23_7  (
            .in0(N__38069),
            .in1(N__41478),
            .in2(N__41419),
            .in3(N__41321),
            .lcout(\c0.n16718 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i18_LC_13_24_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i18_LC_13_24_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i18_LC_13_24_0 .LUT_INIT=16'b1110000011000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i18_LC_13_24_0  (
            .in0(N__44977),
            .in1(N__44677),
            .in2(N__40760),
            .in3(N__44599),
            .lcout(\c0.FRAME_MATCHER_state_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49784),
            .ce(),
            .sr(N__40731));
    defparam \c0.FRAME_MATCHER_state_i27_LC_13_25_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i27_LC_13_25_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i27_LC_13_25_0 .LUT_INIT=16'b1110101000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i27_LC_13_25_0  (
            .in0(N__44718),
            .in1(N__44565),
            .in2(N__45017),
            .in3(N__38065),
            .lcout(\c0.FRAME_MATCHER_state_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49794),
            .ce(),
            .sr(N__38043));
    defparam \c0.data_out_8__0__2192_LC_13_26_0 .C_ON=1'b0;
    defparam \c0.data_out_8__0__2192_LC_13_26_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_8__0__2192_LC_13_26_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.data_out_8__0__2192_LC_13_26_0  (
            .in0(N__38031),
            .in1(N__45406),
            .in2(_gnd_net_),
            .in3(N__49935),
            .lcout(\c0.data_out_8_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49804),
            .ce(),
            .sr(_gnd_net_));
    defparam i53_4_lut_LC_13_26_1.C_ON=1'b0;
    defparam i53_4_lut_LC_13_26_1.SEQ_MODE=4'b0000;
    defparam i53_4_lut_LC_13_26_1.LUT_INIT=16'b1100110011111010;
    LogicCell40 i53_4_lut_LC_13_26_1 (
            .in0(N__47792),
            .in1(N__38001),
            .in2(N__38136),
            .in3(N__47454),
            .lcout(n23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i7_3_lut_LC_13_26_2 .C_ON=1'b0;
    defparam \c0.i7_3_lut_LC_13_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.i7_3_lut_LC_13_26_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.i7_3_lut_LC_13_26_2  (
            .in0(N__49006),
            .in1(N__48827),
            .in2(_gnd_net_),
            .in3(N__47793),
            .lcout(\c0.n3_adj_2193 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_2__0__2240_LC_13_26_3 .C_ON=1'b0;
    defparam \c0.data_out_2__0__2240_LC_13_26_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_2__0__2240_LC_13_26_3 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \c0.data_out_2__0__2240_LC_13_26_3  (
            .in0(N__50541),
            .in1(N__50154),
            .in2(_gnd_net_),
            .in3(N__37995),
            .lcout(data_out_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49804),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_8__7__2185_LC_13_26_4 .C_ON=1'b0;
    defparam \c0.data_out_8__7__2185_LC_13_26_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_8__7__2185_LC_13_26_4 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \c0.data_out_8__7__2185_LC_13_26_4  (
            .in0(N__38157),
            .in1(_gnd_net_),
            .in2(N__45837),
            .in3(N__49934),
            .lcout(data_out_8_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49804),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__0__2256_LC_13_26_5 .C_ON=1'b0;
    defparam \c0.data_out_0__0__2256_LC_13_26_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__0__2256_LC_13_26_5 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \c0.data_out_0__0__2256_LC_13_26_5  (
            .in0(N__38135),
            .in1(N__48150),
            .in2(N__50574),
            .in3(N__50155),
            .lcout(data_out_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49804),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__0__2208_LC_13_26_6 .C_ON=1'b0;
    defparam \c0.data_out_6__0__2208_LC_13_26_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__0__2208_LC_13_26_6 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \c0.data_out_6__0__2208_LC_13_26_6  (
            .in0(N__38124),
            .in1(N__50542),
            .in2(N__43719),
            .in3(N__46817),
            .lcout(\c0.data_out_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49804),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_473_LC_13_26_7 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_473_LC_13_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_473_LC_13_26_7 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_473_LC_13_26_7  (
            .in0(N__45405),
            .in1(N__46507),
            .in2(N__45513),
            .in3(N__46759),
            .lcout(\c0.n17147 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_LC_13_27_0 .C_ON=1'b0;
    defparam \c0.i5_3_lut_LC_13_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_LC_13_27_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.i5_3_lut_LC_13_27_0  (
            .in0(N__47796),
            .in1(N__43308),
            .in2(_gnd_net_),
            .in3(N__48925),
            .lcout(\c0.n1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__7__2193_LC_13_27_1 .C_ON=1'b0;
    defparam \c0.data_out_7__7__2193_LC_13_27_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__7__2193_LC_13_27_1 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \c0.data_out_7__7__2193_LC_13_27_1  (
            .in0(N__43309),
            .in1(N__38103),
            .in2(N__43716),
            .in3(N__46922),
            .lcout(\c0.data_out_7_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49811),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_4_lut_adj_780_LC_13_27_2.C_ON=1'b0;
    defparam i24_4_lut_adj_780_LC_13_27_2.SEQ_MODE=4'b0000;
    defparam i24_4_lut_adj_780_LC_13_27_2.LUT_INIT=16'b0010001011100010;
    LogicCell40 i24_4_lut_adj_780_LC_13_27_2 (
            .in0(N__38166),
            .in1(N__46413),
            .in2(N__38082),
            .in3(N__46298),
            .lcout(),
            .ltout(n10_adj_2411_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i2_LC_13_27_3 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i2_LC_13_27_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i2_LC_13_27_3 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \c0.tx.r_Tx_Data_i2_LC_13_27_3  (
            .in0(N__44103),
            .in1(N__38265),
            .in2(N__38073),
            .in3(N__43815),
            .lcout(r_Tx_Data_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49811),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15044_4_lut_LC_13_27_4 .C_ON=1'b0;
    defparam \c0.i15044_4_lut_LC_13_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.i15044_4_lut_LC_13_27_4 .LUT_INIT=16'b0110000010010000;
    LogicCell40 \c0.i15044_4_lut_LC_13_27_4  (
            .in0(N__46784),
            .in1(N__42518),
            .in2(N__48404),
            .in3(N__44288),
            .lcout(\c0.n17653 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_449_LC_13_27_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_449_LC_13_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_449_LC_13_27_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_449_LC_13_27_7  (
            .in0(_gnd_net_),
            .in1(N__42323),
            .in2(_gnd_net_),
            .in3(N__48465),
            .lcout(\c0.n10392 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_697_LC_13_28_2 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_697_LC_13_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_697_LC_13_28_2 .LUT_INIT=16'b1000110110001000;
    LogicCell40 \c0.i1_4_lut_adj_697_LC_13_28_2  (
            .in0(N__50204),
            .in1(N__38349),
            .in2(N__48144),
            .in3(N__42655),
            .lcout(n4_adj_2414),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.UART_TRANSMITTER_state__i3_LC_13_28_3 .C_ON=1'b0;
    defparam \c0.UART_TRANSMITTER_state__i3_LC_13_28_3 .SEQ_MODE=4'b1000;
    defparam \c0.UART_TRANSMITTER_state__i3_LC_13_28_3 .LUT_INIT=16'b0010001001110010;
    LogicCell40 \c0.UART_TRANSMITTER_state__i3_LC_13_28_3  (
            .in0(N__48302),
            .in1(N__38220),
            .in2(N__43715),
            .in3(N__38280),
            .lcout(UART_TRANSMITTER_state_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49819),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_2_i5_3_lut_LC_13_28_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_2_i5_3_lut_LC_13_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_2_i5_3_lut_LC_13_28_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_2_i5_3_lut_LC_13_28_4  (
            .in0(N__43465),
            .in1(N__46997),
            .in2(_gnd_net_),
            .in3(N__47671),
            .lcout(\c0.n5_adj_2141 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam r_Bit_Index_2__bdd_4_lut_LC_13_28_5.C_ON=1'b0;
    defparam r_Bit_Index_2__bdd_4_lut_LC_13_28_5.SEQ_MODE=4'b0000;
    defparam r_Bit_Index_2__bdd_4_lut_LC_13_28_5.LUT_INIT=16'b1010111111000000;
    LogicCell40 r_Bit_Index_2__bdd_4_lut_LC_13_28_5 (
            .in0(N__43758),
            .in1(N__38264),
            .in2(N__42636),
            .in3(N__42555),
            .lcout(),
            .ltout(n18196_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n18196_bdd_4_lut_LC_13_28_6.C_ON=1'b0;
    defparam n18196_bdd_4_lut_LC_13_28_6.SEQ_MODE=4'b0000;
    defparam n18196_bdd_4_lut_LC_13_28_6.LUT_INIT=16'b1111000011001010;
    LogicCell40 n18196_bdd_4_lut_LC_13_28_6 (
            .in0(N__43515),
            .in1(N__38253),
            .in2(N__38235),
            .in3(N__42624),
            .lcout(n18199),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i26_3_lut_LC_13_28_7 .C_ON=1'b0;
    defparam \c0.tx.i26_3_lut_LC_13_28_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i26_3_lut_LC_13_28_7 .LUT_INIT=16'b0100010001100110;
    LogicCell40 \c0.tx.i26_3_lut_LC_13_28_7  (
            .in0(N__44208),
            .in1(N__44015),
            .in2(_gnd_net_),
            .in3(N__38226),
            .lcout(\c0.tx.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15178_4_lut_LC_13_29_0.C_ON=1'b0;
    defparam i15178_4_lut_LC_13_29_0.SEQ_MODE=4'b0000;
    defparam i15178_4_lut_LC_13_29_0.LUT_INIT=16'b0000001100000010;
    LogicCell40 i15178_4_lut_LC_13_29_0 (
            .in0(N__50270),
            .in1(N__38341),
            .in2(N__48100),
            .in3(N__42656),
            .lcout(n17759),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15020_4_lut_LC_13_29_1.C_ON=1'b0;
    defparam i15020_4_lut_LC_13_29_1.SEQ_MODE=4'b0000;
    defparam i15020_4_lut_LC_13_29_1.LUT_INIT=16'b1111000111110011;
    LogicCell40 i15020_4_lut_LC_13_29_1 (
            .in0(N__38424),
            .in1(N__42671),
            .in2(N__50721),
            .in3(N__43040),
            .lcout(n17664),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18166_bdd_4_lut_LC_13_29_2 .C_ON=1'b0;
    defparam \c0.n18166_bdd_4_lut_LC_13_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.n18166_bdd_4_lut_LC_13_29_2 .LUT_INIT=16'b1010101011011000;
    LogicCell40 \c0.n18166_bdd_4_lut_LC_13_29_2  (
            .in0(N__38205),
            .in1(N__38196),
            .in2(N__38184),
            .in3(N__46254),
            .lcout(n18169),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i149_3_lut_LC_13_29_3 .C_ON=1'b0;
    defparam \c0.i149_3_lut_LC_13_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.i149_3_lut_LC_13_29_3 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \c0.i149_3_lut_LC_13_29_3  (
            .in0(N__50688),
            .in1(N__42670),
            .in2(_gnd_net_),
            .in3(N__43039),
            .lcout(\c0.n453 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i14639_4_lut_LC_13_29_4.C_ON=1'b0;
    defparam i14639_4_lut_LC_13_29_4.SEQ_MODE=4'b0000;
    defparam i14639_4_lut_LC_13_29_4.LUT_INIT=16'b1111101011101010;
    LogicCell40 i14639_4_lut_LC_13_29_4 (
            .in0(N__50271),
            .in1(N__38342),
            .in2(N__48410),
            .in3(N__42657),
            .lcout(n17416),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i7_LC_13_29_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i7_LC_13_29_5 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i7_LC_13_29_5 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \c0.byte_transmit_counter__i7_LC_13_29_5  (
            .in0(N__42699),
            .in1(N__42351),
            .in2(N__42462),
            .in3(N__43076),
            .lcout(byte_transmit_counter_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49826),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10532_2_lut_3_lut_4_lut_LC_13_29_6 .C_ON=1'b0;
    defparam \c0.i10532_2_lut_3_lut_4_lut_LC_13_29_6 .SEQ_MODE=4'b0000;
    defparam \c0.i10532_2_lut_3_lut_4_lut_LC_13_29_6 .LUT_INIT=16'b1111000010110000;
    LogicCell40 \c0.i10532_2_lut_3_lut_4_lut_LC_13_29_6  (
            .in0(N__50733),
            .in1(N__38570),
            .in2(N__38397),
            .in3(N__38662),
            .lcout(\c0.n19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_733_LC_13_30_0 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_733_LC_13_30_0 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_733_LC_13_30_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i3_4_lut_adj_733_LC_13_30_0  (
            .in0(N__42961),
            .in1(N__42934),
            .in2(N__42989),
            .in3(N__43075),
            .lcout(n9524),
            .ltout(n9524_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_4_lut_adj_736_LC_13_30_1 .C_ON=1'b0;
    defparam \c0.i2_4_lut_adj_736_LC_13_30_1 .SEQ_MODE=4'b0000;
    defparam \c0.i2_4_lut_adj_736_LC_13_30_1 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \c0.i2_4_lut_adj_736_LC_13_30_1  (
            .in0(N__43038),
            .in1(N__42844),
            .in2(N__38310),
            .in3(N__42876),
            .lcout(\c0.n16267 ),
            .ltout(\c0.n16267_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15186_2_lut_3_lut_LC_13_30_2 .C_ON=1'b0;
    defparam \c0.i15186_2_lut_3_lut_LC_13_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.i15186_2_lut_3_lut_LC_13_30_2 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \c0.i15186_2_lut_3_lut_LC_13_30_2  (
            .in0(N__50780),
            .in1(_gnd_net_),
            .in2(N__38307),
            .in3(N__50817),
            .lcout(\c0.n445 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10537_2_lut_3_lut_4_lut_LC_13_30_3 .C_ON=1'b0;
    defparam \c0.i10537_2_lut_3_lut_4_lut_LC_13_30_3 .SEQ_MODE=4'b0000;
    defparam \c0.i10537_2_lut_3_lut_4_lut_LC_13_30_3 .LUT_INIT=16'b1111000011010000;
    LogicCell40 \c0.i10537_2_lut_3_lut_4_lut_LC_13_30_3  (
            .in0(N__38560),
            .in1(N__50698),
            .in2(N__38442),
            .in3(N__38636),
            .lcout(\c0.n23_adj_2314 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10454_2_lut_3_lut_4_lut_LC_13_30_4 .C_ON=1'b0;
    defparam \c0.i10454_2_lut_3_lut_4_lut_LC_13_30_4 .SEQ_MODE=4'b0000;
    defparam \c0.i10454_2_lut_3_lut_4_lut_LC_13_30_4 .LUT_INIT=16'b1100100011001100;
    LogicCell40 \c0.i10454_2_lut_3_lut_4_lut_LC_13_30_4  (
            .in0(N__38635),
            .in1(N__38757),
            .in2(N__50723),
            .in3(N__38559),
            .lcout(\c0.n28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14615_2_lut_4_lut_LC_13_30_5 .C_ON=1'b0;
    defparam \c0.i14615_2_lut_4_lut_LC_13_30_5 .SEQ_MODE=4'b0000;
    defparam \c0.i14615_2_lut_4_lut_LC_13_30_5 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \c0.i14615_2_lut_4_lut_LC_13_30_5  (
            .in0(N__38561),
            .in1(N__50699),
            .in2(N__48411),
            .in3(N__38637),
            .lcout(),
            .ltout(n17392_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.UART_TRANSMITTER_state__i1_LC_13_30_6 .C_ON=1'b0;
    defparam \c0.UART_TRANSMITTER_state__i1_LC_13_30_6 .SEQ_MODE=4'b1000;
    defparam \c0.UART_TRANSMITTER_state__i1_LC_13_30_6 .LUT_INIT=16'b1000101110111011;
    LogicCell40 \c0.UART_TRANSMITTER_state__i1_LC_13_30_6  (
            .in0(N__38475),
            .in1(N__48032),
            .in2(N__38469),
            .in3(N__38466),
            .lcout(UART_TRANSMITTER_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49832),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10566_2_lut_LC_13_30_7 .C_ON=1'b0;
    defparam \c0.i10566_2_lut_LC_13_30_7 .SEQ_MODE=4'b0000;
    defparam \c0.i10566_2_lut_LC_13_30_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i10566_2_lut_LC_13_30_7  (
            .in0(_gnd_net_),
            .in1(N__48021),
            .in2(_gnd_net_),
            .in3(N__50259),
            .lcout(n2594),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10533_2_lut_3_lut_4_lut_LC_13_31_0 .C_ON=1'b0;
    defparam \c0.i10533_2_lut_3_lut_4_lut_LC_13_31_0 .SEQ_MODE=4'b0000;
    defparam \c0.i10533_2_lut_3_lut_4_lut_LC_13_31_0 .LUT_INIT=16'b1111110100000000;
    LogicCell40 \c0.i10533_2_lut_3_lut_4_lut_LC_13_31_0  (
            .in0(N__38568),
            .in1(N__50676),
            .in2(N__38660),
            .in3(N__38505),
            .lcout(\c0.n20_adj_2255 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10_4_lut_adj_741_LC_13_31_1 .C_ON=1'b0;
    defparam \c0.i10_4_lut_adj_741_LC_13_31_1 .SEQ_MODE=4'b0000;
    defparam \c0.i10_4_lut_adj_741_LC_13_31_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i10_4_lut_adj_741_LC_13_31_1  (
            .in0(N__38675),
            .in1(N__38789),
            .in2(N__38370),
            .in3(N__38453),
            .lcout(),
            .ltout(\c0.n24_adj_2389_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i12_4_lut_adj_744_LC_13_31_2 .C_ON=1'b0;
    defparam \c0.i12_4_lut_adj_744_LC_13_31_2 .SEQ_MODE=4'b0000;
    defparam \c0.i12_4_lut_adj_744_LC_13_31_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i12_4_lut_adj_744_LC_13_31_2  (
            .in0(N__38438),
            .in1(N__38771),
            .in2(N__38427),
            .in3(N__38481),
            .lcout(\c0.n26_adj_2391 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14552_2_lut_3_lut_LC_13_31_3 .C_ON=1'b0;
    defparam \c0.i14552_2_lut_3_lut_LC_13_31_3 .SEQ_MODE=4'b0000;
    defparam \c0.i14552_2_lut_3_lut_LC_13_31_3 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \c0.i14552_2_lut_3_lut_LC_13_31_3  (
            .in0(N__50248),
            .in1(N__42845),
            .in2(_gnd_net_),
            .in3(N__42874),
            .lcout(n17327),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i13_4_lut_adj_748_LC_13_31_4 .C_ON=1'b0;
    defparam \c0.i13_4_lut_adj_748_LC_13_31_4 .SEQ_MODE=4'b0000;
    defparam \c0.i13_4_lut_adj_748_LC_13_31_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i13_4_lut_adj_748_LC_13_31_4  (
            .in0(N__38414),
            .in1(N__38733),
            .in2(N__38393),
            .in3(N__38376),
            .lcout(\c0.n9453 ),
            .ltout(\c0.n9453_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10538_2_lut_3_lut_4_lut_LC_13_31_5 .C_ON=1'b0;
    defparam \c0.i10538_2_lut_3_lut_4_lut_LC_13_31_5 .SEQ_MODE=4'b0000;
    defparam \c0.i10538_2_lut_3_lut_4_lut_LC_13_31_5 .LUT_INIT=16'b1010100010101010;
    LogicCell40 \c0.i10538_2_lut_3_lut_4_lut_LC_13_31_5  (
            .in0(N__38369),
            .in1(N__50684),
            .in2(N__38358),
            .in3(N__38567),
            .lcout(\c0.n24_adj_2342 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10527_2_lut_3_lut_4_lut_LC_13_31_6 .C_ON=1'b0;
    defparam \c0.i10527_2_lut_3_lut_4_lut_LC_13_31_6 .SEQ_MODE=4'b0000;
    defparam \c0.i10527_2_lut_3_lut_4_lut_LC_13_31_6 .LUT_INIT=16'b1111110100000000;
    LogicCell40 \c0.i10527_2_lut_3_lut_4_lut_LC_13_31_6  (
            .in0(N__38569),
            .in1(N__50677),
            .in2(N__38661),
            .in3(N__38790),
            .lcout(\c0.n16_adj_2212 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10541_2_lut_3_lut_4_lut_LC_13_31_7 .C_ON=1'b0;
    defparam \c0.i10541_2_lut_3_lut_4_lut_LC_13_31_7 .SEQ_MODE=4'b0000;
    defparam \c0.i10541_2_lut_3_lut_4_lut_LC_13_31_7 .LUT_INIT=16'b1010100010101010;
    LogicCell40 \c0.i10541_2_lut_3_lut_4_lut_LC_13_31_7  (
            .in0(N__38772),
            .in1(N__38639),
            .in2(N__50717),
            .in3(N__38566),
            .lcout(\c0.n26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_743_LC_13_32_0 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_743_LC_13_32_0 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_743_LC_13_32_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i8_4_lut_adj_743_LC_13_32_0  (
            .in0(N__38726),
            .in1(N__38756),
            .in2(N__38712),
            .in3(N__38744),
            .lcout(\c0.n22_adj_2390 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10531_2_lut_3_lut_4_lut_LC_13_32_2 .C_ON=1'b0;
    defparam \c0.i10531_2_lut_3_lut_4_lut_LC_13_32_2 .SEQ_MODE=4'b0000;
    defparam \c0.i10531_2_lut_3_lut_4_lut_LC_13_32_2 .LUT_INIT=16'b1010100010101010;
    LogicCell40 \c0.i10531_2_lut_3_lut_4_lut_LC_13_32_2  (
            .in0(N__38727),
            .in1(N__38652),
            .in2(N__50744),
            .in3(N__38578),
            .lcout(\c0.n18_adj_2220 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10522_2_lut_3_lut_4_lut_LC_13_32_3 .C_ON=1'b0;
    defparam \c0.i10522_2_lut_3_lut_4_lut_LC_13_32_3 .SEQ_MODE=4'b0000;
    defparam \c0.i10522_2_lut_3_lut_4_lut_LC_13_32_3 .LUT_INIT=16'b1111110100000000;
    LogicCell40 \c0.i10522_2_lut_3_lut_4_lut_LC_13_32_3  (
            .in0(N__38580),
            .in1(N__50740),
            .in2(N__38663),
            .in3(N__38711),
            .lcout(\c0.n15_adj_2211 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i5_LC_13_32_5 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i5_LC_13_32_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i5_LC_13_32_5 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \c0.tx.r_Tx_Data_i5_LC_13_32_5  (
            .in0(N__38690),
            .in1(N__43290),
            .in2(N__44106),
            .in3(N__43845),
            .lcout(r_Tx_Data_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49838),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10528_2_lut_3_lut_4_lut_LC_13_32_6 .C_ON=1'b0;
    defparam \c0.i10528_2_lut_3_lut_4_lut_LC_13_32_6 .SEQ_MODE=4'b0000;
    defparam \c0.i10528_2_lut_3_lut_4_lut_LC_13_32_6 .LUT_INIT=16'b1010100010101010;
    LogicCell40 \c0.i10528_2_lut_3_lut_4_lut_LC_13_32_6  (
            .in0(N__38676),
            .in1(N__38653),
            .in2(N__50745),
            .in3(N__38579),
            .lcout(\c0.n17_adj_2219 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_2_lut_LC_13_32_7 .C_ON=1'b0;
    defparam \c0.i4_2_lut_LC_13_32_7 .SEQ_MODE=4'b0000;
    defparam \c0.i4_2_lut_LC_13_32_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.i4_2_lut_LC_13_32_7  (
            .in0(_gnd_net_),
            .in1(N__38504),
            .in2(_gnd_net_),
            .in3(N__38492),
            .lcout(\c0.n18_adj_2388 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter2_i5_LC_14_17_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter2_i5_LC_14_17_0 .SEQ_MODE=4'b1001;
    defparam \c0.byte_transmit_counter2_i5_LC_14_17_0 .LUT_INIT=16'b1100101000000000;
    LogicCell40 \c0.byte_transmit_counter2_i5_LC_14_17_0  (
            .in0(N__39711),
            .in1(N__39612),
            .in2(N__39697),
            .in3(N__42094),
            .lcout(\c0.byte_transmit_counter2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49711),
            .ce(),
            .sr(N__39588));
    defparam \c0.rx.r_Rx_Byte_i6_LC_14_18_1 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i6_LC_14_18_1 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i6_LC_14_18_1 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \c0.rx.r_Rx_Byte_i6_LC_14_18_1  (
            .in0(N__45220),
            .in1(N__39576),
            .in2(N__39523),
            .in3(N__45177),
            .lcout(rx_data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49727),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i1_3_lut_LC_14_18_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i1_3_lut_LC_14_18_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i1_3_lut_LC_14_18_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_6_i1_3_lut_LC_14_18_2  (
            .in0(N__45054),
            .in1(N__45315),
            .in2(_gnd_net_),
            .in3(N__47846),
            .lcout(\c0.n1_adj_2160 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i26_LC_14_18_3 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i26_LC_14_18_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i26_LC_14_18_3 .LUT_INIT=16'b1100110011011000;
    LogicCell40 \c0.data_in_frame_0__i26_LC_14_18_3  (
            .in0(N__40567),
            .in1(N__39281),
            .in2(N__39462),
            .in3(N__39395),
            .lcout(\c0.data_in_frame_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49727),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14695_4_lut_LC_14_18_4 .C_ON=1'b0;
    defparam \c0.i14695_4_lut_LC_14_18_4 .SEQ_MODE=4'b0000;
    defparam \c0.i14695_4_lut_LC_14_18_4 .LUT_INIT=16'b1111101011010000;
    LogicCell40 \c0.i14695_4_lut_LC_14_18_4  (
            .in0(N__39835),
            .in1(N__40317),
            .in2(N__39258),
            .in3(N__40145),
            .lcout(),
            .ltout(\c0.n17472_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i7_LC_14_18_5 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i7_LC_14_18_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i7_LC_14_18_5 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \c0.data_out_frame2_0___i7_LC_14_18_5  (
            .in0(N__39837),
            .in1(N__39951),
            .in2(N__39267),
            .in3(N__39879),
            .lcout(\c0.data_out_frame2_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49727),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_2__2__2275_LC_14_19_0 .C_ON=1'b0;
    defparam \c0.data_in_2__2__2275_LC_14_19_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_2__2__2275_LC_14_19_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_in_2__2__2275_LC_14_19_0  (
            .in0(N__39222),
            .in1(N__38985),
            .in2(_gnd_net_),
            .in3(N__38922),
            .lcout(data_in_2_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49737),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_633_LC_14_19_2 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_633_LC_14_19_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_633_LC_14_19_2 .LUT_INIT=16'b1110101110111110;
    LogicCell40 \c0.i5_4_lut_adj_633_LC_14_19_2  (
            .in0(N__39957),
            .in1(N__38901),
            .in2(N__38853),
            .in3(N__38832),
            .lcout(\c0.n21_adj_2357 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14713_4_lut_LC_14_19_3 .C_ON=1'b0;
    defparam \c0.i14713_4_lut_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \c0.i14713_4_lut_LC_14_19_3 .LUT_INIT=16'b1111110010110000;
    LogicCell40 \c0.i14713_4_lut_LC_14_19_3  (
            .in0(N__40313),
            .in1(N__39831),
            .in2(N__40663),
            .in3(N__40140),
            .lcout(\c0.n17490 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_in_frame_0__i16_LC_14_19_5 .C_ON=1'b0;
    defparam \c0.data_in_frame_0__i16_LC_14_19_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_in_frame_0__i16_LC_14_19_5 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.data_in_frame_0__i16_LC_14_19_5  (
            .in0(N__40598),
            .in1(N__40499),
            .in2(N__40984),
            .in3(N__40431),
            .lcout(\c0.data_in_frame_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49737),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14710_4_lut_LC_14_19_6 .C_ON=1'b0;
    defparam \c0.i14710_4_lut_LC_14_19_6 .SEQ_MODE=4'b0000;
    defparam \c0.i14710_4_lut_LC_14_19_6 .LUT_INIT=16'b1110110010101100;
    LogicCell40 \c0.i14710_4_lut_LC_14_19_6  (
            .in0(N__40141),
            .in1(N__40272),
            .in2(N__39844),
            .in3(N__40314),
            .lcout(),
            .ltout(\c0.n17487_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i2_LC_14_19_7 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i2_LC_14_19_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i2_LC_14_19_7 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \c0.data_out_frame2_0___i2_LC_14_19_7  (
            .in0(N__39836),
            .in1(N__39876),
            .in2(N__40293),
            .in3(N__39947),
            .lcout(\c0.data_out_frame2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49737),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15061_3_lut_4_lut_LC_14_20_3 .C_ON=1'b0;
    defparam \c0.i15061_3_lut_4_lut_LC_14_20_3 .SEQ_MODE=4'b0000;
    defparam \c0.i15061_3_lut_4_lut_LC_14_20_3 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \c0.i15061_3_lut_4_lut_LC_14_20_3  (
            .in0(N__41968),
            .in1(N__40247),
            .in2(N__40089),
            .in3(N__40142),
            .lcout(),
            .ltout(\c0.n17690_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_frame2_0___i3_LC_14_20_4 .C_ON=1'b0;
    defparam \c0.data_out_frame2_0___i3_LC_14_20_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_frame2_0___i3_LC_14_20_4 .LUT_INIT=16'b1111101001000100;
    LogicCell40 \c0.data_out_frame2_0___i3_LC_14_20_4  (
            .in0(N__39944),
            .in1(N__40079),
            .in2(N__40107),
            .in3(N__39724),
            .lcout(\c0.data_out_frame2_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49748),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_adj_622_LC_14_20_5 .C_ON=1'b0;
    defparam \c0.i1_3_lut_adj_622_LC_14_20_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_adj_622_LC_14_20_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_3_lut_adj_622_LC_14_20_5  (
            .in0(N__40049),
            .in1(N__40026),
            .in2(_gnd_net_),
            .in3(N__39999),
            .lcout(\c0.n17102 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n5817_bdd_4_lut_15430_4_lut_LC_14_20_6 .C_ON=1'b0;
    defparam \c0.n5817_bdd_4_lut_15430_4_lut_LC_14_20_6 .SEQ_MODE=4'b0000;
    defparam \c0.n5817_bdd_4_lut_15430_4_lut_LC_14_20_6 .LUT_INIT=16'b0101100011111000;
    LogicCell40 \c0.n5817_bdd_4_lut_15430_4_lut_LC_14_20_6  (
            .in0(N__39943),
            .in1(N__39874),
            .in2(N__39845),
            .in3(N__39759),
            .lcout(\c0.n18202 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i29_LC_14_21_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i29_LC_14_21_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i29_LC_14_21_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i29_LC_14_21_0  (
            .in0(_gnd_net_),
            .in1(N__41228),
            .in2(_gnd_net_),
            .in3(N__41552),
            .lcout(\c0.FRAME_MATCHER_state_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49760),
            .ce(),
            .sr(N__41208));
    defparam \c0.FRAME_MATCHER_state_i10_LC_14_22_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i10_LC_14_22_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i10_LC_14_22_0 .LUT_INIT=16'b1110000011000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i10_LC_14_22_0  (
            .in0(N__44975),
            .in1(N__44673),
            .in2(N__41193),
            .in3(N__44510),
            .lcout(\c0.FRAME_MATCHER_state_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49773),
            .ce(),
            .sr(N__41169));
    defparam \c0.i1_2_lut_adj_488_LC_14_22_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_488_LC_14_22_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_488_LC_14_22_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_488_LC_14_22_2  (
            .in0(N__41145),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41109),
            .lcout(\c0.n17315 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_543_LC_14_22_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_543_LC_14_22_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_543_LC_14_22_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_543_LC_14_22_3  (
            .in0(N__41032),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40978),
            .lcout(\c0.n17213 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_551_LC_14_22_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_551_LC_14_22_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_551_LC_14_22_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_551_LC_14_22_4  (
            .in0(_gnd_net_),
            .in1(N__40933),
            .in2(_gnd_net_),
            .in3(N__40891),
            .lcout(\c0.n10472 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_715_LC_14_22_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_715_LC_14_22_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_715_LC_14_22_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i1_2_lut_adj_715_LC_14_22_5  (
            .in0(N__43183),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40820),
            .lcout(\c0.n8_adj_2330 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_719_LC_14_22_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_719_LC_14_22_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_719_LC_14_22_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i1_2_lut_adj_719_LC_14_22_6  (
            .in0(N__40821),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40759),
            .lcout(\c0.n8_adj_2329 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_728_LC_14_22_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_728_LC_14_22_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_728_LC_14_22_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i1_2_lut_adj_728_LC_14_22_7  (
            .in0(_gnd_net_),
            .in1(N__43150),
            .in2(_gnd_net_),
            .in3(N__40719),
            .lcout(\c0.n16686 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i17_4_lut_LC_14_23_0 .C_ON=1'b0;
    defparam \c0.i17_4_lut_LC_14_23_0 .SEQ_MODE=4'b0000;
    defparam \c0.i17_4_lut_LC_14_23_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i17_4_lut_LC_14_23_0  (
            .in0(N__41524),
            .in1(N__43264),
            .in2(N__43230),
            .in3(N__44372),
            .lcout(\c0.n46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_732_LC_14_23_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_732_LC_14_23_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_732_LC_14_23_1 .LUT_INIT=16'b1010101000001000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_732_LC_14_23_1  (
            .in0(N__41525),
            .in1(N__41493),
            .in2(N__41420),
            .in3(N__41334),
            .lcout(\c0.n16700 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i260_2_lut_3_lut_LC_14_23_2 .C_ON=1'b0;
    defparam \c0.i260_2_lut_3_lut_LC_14_23_2 .SEQ_MODE=4'b0000;
    defparam \c0.i260_2_lut_3_lut_LC_14_23_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.i260_2_lut_3_lut_LC_14_23_2  (
            .in0(N__42040),
            .in1(N__41972),
            .in2(_gnd_net_),
            .in3(N__41858),
            .lcout(\c0.n276 ),
            .ltout(\c0.n276_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_404_LC_14_23_3 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_404_LC_14_23_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_404_LC_14_23_3 .LUT_INIT=16'b1111001011110000;
    LogicCell40 \c0.i1_4_lut_adj_404_LC_14_23_3  (
            .in0(N__41859),
            .in1(N__41605),
            .in2(N__41559),
            .in3(N__44513),
            .lcout(\c0.n4_adj_2135 ),
            .ltout(\c0.n4_adj_2135_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i31_LC_14_23_4 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i31_LC_14_23_4 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i31_LC_14_23_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i31_LC_14_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__41529),
            .in3(N__41526),
            .lcout(\c0.FRAME_MATCHER_state_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49785),
            .ce(),
            .sr(N__41511));
    defparam \c0.i1_2_lut_4_lut_adj_755_LC_14_23_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_755_LC_14_23_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_755_LC_14_23_5 .LUT_INIT=16'b1010101000001000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_755_LC_14_23_5  (
            .in0(N__44373),
            .in1(N__41494),
            .in2(N__41421),
            .in3(N__41335),
            .lcout(\c0.n16714 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_760_LC_14_23_6 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_760_LC_14_23_6 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_760_LC_14_23_6 .LUT_INIT=16'b1011101000000000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_760_LC_14_23_6  (
            .in0(N__41336),
            .in1(N__41407),
            .in2(N__41499),
            .in3(N__43265),
            .lcout(\c0.n16690 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_761_LC_14_23_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_761_LC_14_23_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_761_LC_14_23_7 .LUT_INIT=16'b1010101000001000;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_761_LC_14_23_7  (
            .in0(N__43229),
            .in1(N__41498),
            .in2(N__41422),
            .in3(N__41337),
            .lcout(\c0.n16702 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i17_LC_14_24_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i17_LC_14_24_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i17_LC_14_24_0 .LUT_INIT=16'b1110000011000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i17_LC_14_24_0  (
            .in0(N__44978),
            .in1(N__44674),
            .in2(N__41264),
            .in3(N__44600),
            .lcout(\c0.FRAME_MATCHER_state_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49795),
            .ce(),
            .sr(N__42222));
    defparam \c0.data_out_9__3__2181_LC_14_25_0 .C_ON=1'b0;
    defparam \c0.data_out_9__3__2181_LC_14_25_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_9__3__2181_LC_14_25_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_9__3__2181_LC_14_25_0  (
            .in0(N__43407),
            .in1(N__45620),
            .in2(N__46599),
            .in3(N__43533),
            .lcout(\c0.data_out_9_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49805),
            .ce(N__49970),
            .sr(_gnd_net_));
    defparam \c0.i8_4_lut_adj_463_LC_14_25_2 .C_ON=1'b0;
    defparam \c0.i8_4_lut_adj_463_LC_14_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.i8_4_lut_adj_463_LC_14_25_2 .LUT_INIT=16'b0010111000100010;
    LogicCell40 \c0.i8_4_lut_adj_463_LC_14_25_2  (
            .in0(N__42216),
            .in1(N__47488),
            .in2(N__47847),
            .in3(N__45671),
            .lcout(n10_adj_2431),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_10__3__2173_LC_14_25_3 .C_ON=1'b0;
    defparam \c0.data_out_10__3__2173_LC_14_25_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_10__3__2173_LC_14_25_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_out_10__3__2173_LC_14_25_3  (
            .in0(N__49005),
            .in1(N__42177),
            .in2(_gnd_net_),
            .in3(N__46626),
            .lcout(\c0.data_out_10_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49805),
            .ce(N__49970),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_512_LC_14_25_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_512_LC_14_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_512_LC_14_25_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_512_LC_14_25_4  (
            .in0(_gnd_net_),
            .in1(N__45670),
            .in2(_gnd_net_),
            .in3(N__46696),
            .lcout(\c0.n6_adj_2221 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i6_4_lut_adj_437_LC_14_25_6 .C_ON=1'b0;
    defparam \c0.i6_4_lut_adj_437_LC_14_25_6 .SEQ_MODE=4'b0000;
    defparam \c0.i6_4_lut_adj_437_LC_14_25_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i6_4_lut_adj_437_LC_14_25_6  (
            .in0(N__42176),
            .in1(N__43431),
            .in2(N__45696),
            .in3(N__48500),
            .lcout(\c0.n15_adj_2177 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__0__2200_LC_14_26_1 .C_ON=1'b0;
    defparam \c0.data_out_7__0__2200_LC_14_26_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__0__2200_LC_14_26_1 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \c0.data_out_7__0__2200_LC_14_26_1  (
            .in0(N__48156),
            .in1(N__42168),
            .in2(N__50314),
            .in3(N__42150),
            .lcout(\c0.data_out_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49812),
            .ce(N__46934),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_489_LC_14_26_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_489_LC_14_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_489_LC_14_26_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_489_LC_14_26_3  (
            .in0(N__45398),
            .in1(N__42144),
            .in2(_gnd_net_),
            .in3(N__43313),
            .lcout(\c0.n10183 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_LC_14_26_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_LC_14_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_LC_14_26_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_LC_14_26_4  (
            .in0(N__46506),
            .in1(N__47124),
            .in2(_gnd_net_),
            .in3(N__49111),
            .lcout(\c0.n17129 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15405_LC_14_27_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15405_LC_14_27_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15405_LC_14_27_0 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \c0.byte_transmit_counter_1__bdd_4_lut_15405_LC_14_27_0  (
            .in0(N__42276),
            .in1(N__46295),
            .in2(N__42309),
            .in3(N__47486),
            .lcout(),
            .ltout(\c0.n18184_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18184_bdd_4_lut_LC_14_27_1 .C_ON=1'b0;
    defparam \c0.n18184_bdd_4_lut_LC_14_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.n18184_bdd_4_lut_LC_14_27_1 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \c0.n18184_bdd_4_lut_LC_14_27_1  (
            .in0(N__46296),
            .in1(N__42108),
            .in2(N__42099),
            .in3(N__42270),
            .lcout(),
            .ltout(n18187_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_4_lut_adj_773_LC_14_27_2.C_ON=1'b0;
    defparam i24_4_lut_adj_773_LC_14_27_2.SEQ_MODE=4'b0000;
    defparam i24_4_lut_adj_773_LC_14_27_2.LUT_INIT=16'b0101000011011000;
    LogicCell40 i24_4_lut_adj_773_LC_14_27_2 (
            .in0(N__46402),
            .in1(N__43908),
            .in2(N__42327),
            .in3(N__46297),
            .lcout(n10_adj_2443),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i5_3_lut_LC_14_27_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i5_3_lut_LC_14_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i5_3_lut_LC_14_27_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_6_i5_3_lut_LC_14_27_4  (
            .in0(N__47256),
            .in1(N__42324),
            .in2(_gnd_net_),
            .in3(N__47812),
            .lcout(\c0.n5_adj_2159 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_5__6__2210_LC_14_27_5 .C_ON=1'b0;
    defparam \c0.data_out_5__6__2210_LC_14_27_5 .SEQ_MODE=4'b1001;
    defparam \c0.data_out_5__6__2210_LC_14_27_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.data_out_5__6__2210_LC_14_27_5  (
            .in0(_gnd_net_),
            .in1(N__48164),
            .in2(_gnd_net_),
            .in3(N__42300),
            .lcout(\c0.data_out_7__2__N_447 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49820),
            .ce(N__50567),
            .sr(N__42793));
    defparam \c0.i15149_2_lut_LC_14_27_6 .C_ON=1'b0;
    defparam \c0.i15149_2_lut_LC_14_27_6 .SEQ_MODE=4'b0000;
    defparam \c0.i15149_2_lut_LC_14_27_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i15149_2_lut_LC_14_27_6  (
            .in0(_gnd_net_),
            .in1(N__47300),
            .in2(_gnd_net_),
            .in3(N__47811),
            .lcout(\c0.n17698 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15119_2_lut_LC_14_27_7 .C_ON=1'b0;
    defparam \c0.i15119_2_lut_LC_14_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.i15119_2_lut_LC_14_27_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i15119_2_lut_LC_14_27_7  (
            .in0(N__47813),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43284),
            .lcout(\c0.n17612 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_452_LC_14_28_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_452_LC_14_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_452_LC_14_28_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_452_LC_14_28_1  (
            .in0(_gnd_net_),
            .in1(N__45836),
            .in2(_gnd_net_),
            .in3(N__47873),
            .lcout(\c0.n10395 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_6__1__2207_LC_14_28_2 .C_ON=1'b0;
    defparam \c0.data_out_6__1__2207_LC_14_28_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_6__1__2207_LC_14_28_2 .LUT_INIT=16'b1111000010111011;
    LogicCell40 \c0.data_out_6__1__2207_LC_14_28_2  (
            .in0(N__43360),
            .in1(N__48303),
            .in2(N__42264),
            .in3(N__50290),
            .lcout(\c0.data_out_6_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49827),
            .ce(N__50548),
            .sr(_gnd_net_));
    defparam i51_4_lut_adj_778_LC_14_28_4.C_ON=1'b0;
    defparam i51_4_lut_adj_778_LC_14_28_4.SEQ_MODE=4'b0000;
    defparam i51_4_lut_adj_778_LC_14_28_4.LUT_INIT=16'b0111001101000000;
    LogicCell40 i51_4_lut_adj_778_LC_14_28_4 (
            .in0(N__46294),
            .in1(N__46403),
            .in2(N__42246),
            .in3(N__42678),
            .lcout(n28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9889_3_lut_LC_14_28_5 .C_ON=1'b0;
    defparam \c0.i9889_3_lut_LC_14_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.i9889_3_lut_LC_14_28_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.i9889_3_lut_LC_14_28_5  (
            .in0(N__48652),
            .in1(N__46750),
            .in2(_gnd_net_),
            .in3(N__47820),
            .lcout(),
            .ltout(n5_adj_2448_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i53_4_lut_adj_776_LC_14_28_6.C_ON=1'b0;
    defparam i53_4_lut_adj_776_LC_14_28_6.SEQ_MODE=4'b0000;
    defparam i53_4_lut_adj_776_LC_14_28_6.LUT_INIT=16'b1111000010001000;
    LogicCell40 i53_4_lut_adj_776_LC_14_28_6 (
            .in0(N__47874),
            .in1(N__47821),
            .in2(N__42684),
            .in3(N__47484),
            .lcout(),
            .ltout(n31_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i49_4_lut_adj_777_LC_14_28_7.C_ON=1'b0;
    defparam i49_4_lut_adj_777_LC_14_28_7.SEQ_MODE=4'b0000;
    defparam i49_4_lut_adj_777_LC_14_28_7.LUT_INIT=16'b1111000000100010;
    LogicCell40 i49_4_lut_adj_777_LC_14_28_7 (
            .in0(N__43563),
            .in1(N__47485),
            .in2(N__42681),
            .in3(N__46293),
            .lcout(n22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i146_4_lut_LC_14_29_1 .C_ON=1'b0;
    defparam \c0.i146_4_lut_LC_14_29_1 .SEQ_MODE=4'b0000;
    defparam \c0.i146_4_lut_LC_14_29_1 .LUT_INIT=16'b1111000011110111;
    LogicCell40 \c0.i146_4_lut_LC_14_29_1  (
            .in0(N__42816),
            .in1(N__43041),
            .in2(N__50722),
            .in3(N__42672),
            .lcout(n450),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i15099_4_lut_LC_14_29_2 .C_ON=1'b0;
    defparam \c0.tx.i15099_4_lut_LC_14_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i15099_4_lut_LC_14_29_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.tx.i15099_4_lut_LC_14_29_2  (
            .in0(N__42642),
            .in1(N__43938),
            .in2(N__42591),
            .in3(N__42554),
            .lcout(),
            .ltout(\c0.tx.n17673_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i29_3_lut_LC_14_29_3 .C_ON=1'b0;
    defparam \c0.tx.i29_3_lut_LC_14_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i29_3_lut_LC_14_29_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \c0.tx.i29_3_lut_LC_14_29_3  (
            .in0(N__44179),
            .in1(_gnd_net_),
            .in2(N__42522),
            .in3(N__50823),
            .lcout(\c0.tx.n12_adj_2134 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_LC_14_29_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_LC_14_29_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_LC_14_29_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_LC_14_29_5  (
            .in0(N__47106),
            .in1(N__49084),
            .in2(N__42519),
            .in3(N__47313),
            .lcout(\c0.n17126 ),
            .ltout(\c0.n17126_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15003_3_lut_LC_14_29_6 .C_ON=1'b0;
    defparam \c0.i15003_3_lut_LC_14_29_6 .SEQ_MODE=4'b0000;
    defparam \c0.i15003_3_lut_LC_14_29_6 .LUT_INIT=16'b1010000000001010;
    LogicCell40 \c0.i15003_3_lut_LC_14_29_6  (
            .in0(N__48313),
            .in1(_gnd_net_),
            .in2(N__42477),
            .in3(N__46509),
            .lcout(\c0.n17651 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter__i5_LC_14_29_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter__i5_LC_14_29_7 .SEQ_MODE=4'b1000;
    defparam \c0.byte_transmit_counter__i5_LC_14_29_7 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \c0.byte_transmit_counter__i5_LC_14_29_7  (
            .in0(N__42735),
            .in1(N__42460),
            .in2(N__42966),
            .in3(N__42365),
            .lcout(byte_transmit_counter_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49833),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2506_2_lut_LC_14_30_0 .C_ON=1'b1;
    defparam \c0.add_2506_2_lut_LC_14_30_0 .SEQ_MODE=4'b0000;
    defparam \c0.add_2506_2_lut_LC_14_30_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_2506_2_lut_LC_14_30_0  (
            .in0(_gnd_net_),
            .in1(N__44022),
            .in2(N__47825),
            .in3(_gnd_net_),
            .lcout(tx_transmit_N_1947_0),
            .ltout(),
            .carryin(bfn_14_30_0_),
            .carryout(\c0.n16110 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2506_3_lut_LC_14_30_1 .C_ON=1'b1;
    defparam \c0.add_2506_3_lut_LC_14_30_1 .SEQ_MODE=4'b0000;
    defparam \c0.add_2506_3_lut_LC_14_30_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_2506_3_lut_LC_14_30_1  (
            .in0(_gnd_net_),
            .in1(N__47483),
            .in2(_gnd_net_),
            .in3(N__42747),
            .lcout(tx_transmit_N_1947_1),
            .ltout(),
            .carryin(\c0.n16110 ),
            .carryout(\c0.n16111 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2506_4_lut_LC_14_30_2 .C_ON=1'b1;
    defparam \c0.add_2506_4_lut_LC_14_30_2 .SEQ_MODE=4'b0000;
    defparam \c0.add_2506_4_lut_LC_14_30_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_2506_4_lut_LC_14_30_2  (
            .in0(_gnd_net_),
            .in1(N__46291),
            .in2(_gnd_net_),
            .in3(N__42744),
            .lcout(tx_transmit_N_1947_2),
            .ltout(),
            .carryin(\c0.n16111 ),
            .carryout(\c0.n16112 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2506_5_lut_LC_14_30_3 .C_ON=1'b1;
    defparam \c0.add_2506_5_lut_LC_14_30_3 .SEQ_MODE=4'b0000;
    defparam \c0.add_2506_5_lut_LC_14_30_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_2506_5_lut_LC_14_30_3  (
            .in0(_gnd_net_),
            .in1(N__46401),
            .in2(_gnd_net_),
            .in3(N__42741),
            .lcout(tx_transmit_N_1947_3),
            .ltout(),
            .carryin(\c0.n16112 ),
            .carryout(\c0.n16113 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2506_6_lut_LC_14_30_4 .C_ON=1'b1;
    defparam \c0.add_2506_6_lut_LC_14_30_4 .SEQ_MODE=4'b0000;
    defparam \c0.add_2506_6_lut_LC_14_30_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_2506_6_lut_LC_14_30_4  (
            .in0(_gnd_net_),
            .in1(N__43836),
            .in2(_gnd_net_),
            .in3(N__42738),
            .lcout(tx_transmit_N_1947_4),
            .ltout(),
            .carryin(\c0.n16113 ),
            .carryout(\c0.n16114 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2506_7_lut_LC_14_30_5 .C_ON=1'b1;
    defparam \c0.add_2506_7_lut_LC_14_30_5 .SEQ_MODE=4'b0000;
    defparam \c0.add_2506_7_lut_LC_14_30_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_2506_7_lut_LC_14_30_5  (
            .in0(_gnd_net_),
            .in1(N__42734),
            .in2(_gnd_net_),
            .in3(N__42723),
            .lcout(tx_transmit_N_1947_5),
            .ltout(),
            .carryin(\c0.n16114 ),
            .carryout(\c0.n16115 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2506_8_lut_LC_14_30_6 .C_ON=1'b1;
    defparam \c0.add_2506_8_lut_LC_14_30_6 .SEQ_MODE=4'b0000;
    defparam \c0.add_2506_8_lut_LC_14_30_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_2506_8_lut_LC_14_30_6  (
            .in0(_gnd_net_),
            .in1(N__42720),
            .in2(_gnd_net_),
            .in3(N__42702),
            .lcout(tx_transmit_N_1947_6),
            .ltout(),
            .carryin(\c0.n16115 ),
            .carryout(\c0.n16116 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.add_2506_9_lut_LC_14_30_7 .C_ON=1'b0;
    defparam \c0.add_2506_9_lut_LC_14_30_7 .SEQ_MODE=4'b0000;
    defparam \c0.add_2506_9_lut_LC_14_30_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.add_2506_9_lut_LC_14_30_7  (
            .in0(_gnd_net_),
            .in1(N__42698),
            .in2(_gnd_net_),
            .in3(N__42687),
            .lcout(tx_transmit_N_1947_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_LC_14_31_0 .C_ON=1'b0;
    defparam \c0.i1_4_lut_LC_14_31_0 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_LC_14_31_0 .LUT_INIT=16'b0101000011011100;
    LogicCell40 \c0.i1_4_lut_LC_14_31_0  (
            .in0(N__43043),
            .in1(N__43008),
            .in2(N__43002),
            .in3(N__42875),
            .lcout(),
            .ltout(\c0.n68_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_transmit_2168_LC_14_31_1 .C_ON=1'b0;
    defparam \c0.tx_transmit_2168_LC_14_31_1 .SEQ_MODE=4'b1000;
    defparam \c0.tx_transmit_2168_LC_14_31_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \c0.tx_transmit_2168_LC_14_31_1  (
            .in0(N__48110),
            .in1(N__42918),
            .in2(N__43080),
            .in3(N__43077),
            .lcout(\c0.r_SM_Main_2_N_2034_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49839),
            .ce(),
            .sr(N__43059));
    defparam \c0.i2_3_lut_adj_766_LC_14_31_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_766_LC_14_31_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_766_LC_14_31_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.i2_3_lut_adj_766_LC_14_31_2  (
            .in0(N__48022),
            .in1(N__48314),
            .in2(_gnd_net_),
            .in3(N__50276),
            .lcout(\c0.n4650 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i90_4_lut_LC_14_31_3 .C_ON=1'b0;
    defparam \c0.i90_4_lut_LC_14_31_3 .SEQ_MODE=4'b0000;
    defparam \c0.i90_4_lut_LC_14_31_3 .LUT_INIT=16'b0010001001110010;
    LogicCell40 \c0.i90_4_lut_LC_14_31_3  (
            .in0(N__50275),
            .in1(N__43042),
            .in2(N__48379),
            .in3(N__42842),
            .lcout(\c0.n59 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_3_lut_adj_768_LC_14_31_4 .C_ON=1'b0;
    defparam \c0.i1_3_lut_adj_768_LC_14_31_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_3_lut_adj_768_LC_14_31_4 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \c0.i1_3_lut_adj_768_LC_14_31_4  (
            .in0(N__42843),
            .in1(N__48315),
            .in2(_gnd_net_),
            .in3(N__50277),
            .lcout(\c0.n65 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i14627_4_lut_LC_14_31_5 .C_ON=1'b0;
    defparam \c0.i14627_4_lut_LC_14_31_5 .SEQ_MODE=4'b0000;
    defparam \c0.i14627_4_lut_LC_14_31_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.i14627_4_lut_LC_14_31_5  (
            .in0(N__42985),
            .in1(N__42962),
            .in2(N__50720),
            .in3(N__42935),
            .lcout(\c0.n17404 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i10986_2_lut_LC_14_31_6 .C_ON=1'b0;
    defparam \c0.i10986_2_lut_LC_14_31_6 .SEQ_MODE=4'b0000;
    defparam \c0.i10986_2_lut_LC_14_31_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i10986_2_lut_LC_14_31_6  (
            .in0(_gnd_net_),
            .in1(N__42905),
            .in2(_gnd_net_),
            .in3(N__42887),
            .lcout(\c0.n13662 ),
            .ltout(\c0.n13662_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i11047_2_lut_LC_14_31_7 .C_ON=1'b0;
    defparam \c0.i11047_2_lut_LC_14_31_7 .SEQ_MODE=4'b0000;
    defparam \c0.i11047_2_lut_LC_14_31_7 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \c0.i11047_2_lut_LC_14_31_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42855),
            .in3(N__42841),
            .lcout(\c0.n13726 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15194_2_lut_LC_14_32_1 .C_ON=1'b0;
    defparam \c0.i15194_2_lut_LC_14_32_1 .SEQ_MODE=4'b0000;
    defparam \c0.i15194_2_lut_LC_14_32_1 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \c0.i15194_2_lut_LC_14_32_1  (
            .in0(N__50322),
            .in1(N__50492),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\c0.n10815 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__3__2253_LC_14_32_2 .C_ON=1'b0;
    defparam \c0.data_out_0__3__2253_LC_14_32_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__3__2253_LC_14_32_2 .LUT_INIT=16'b0011111100110000;
    LogicCell40 \c0.data_out_0__3__2253_LC_14_32_2  (
            .in0(_gnd_net_),
            .in1(N__50323),
            .in2(N__50546),
            .in3(N__42761),
            .lcout(data_out_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49844),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_4_lut_adj_790_LC_14_32_4.C_ON=1'b0;
    defparam i24_4_lut_adj_790_LC_14_32_4.SEQ_MODE=4'b0000;
    defparam i24_4_lut_adj_790_LC_14_32_4.LUT_INIT=16'b0010001011100010;
    LogicCell40 i24_4_lut_adj_790_LC_14_32_4 (
            .in0(N__45330),
            .in1(N__46414),
            .in2(N__44223),
            .in3(N__46292),
            .lcout(n10_adj_2483),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_3__6__2226_LC_14_32_6 .C_ON=1'b0;
    defparam \c0.data_out_3__6__2226_LC_14_32_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_3__6__2226_LC_14_32_6 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \c0.data_out_3__6__2226_LC_14_32_6  (
            .in0(N__50319),
            .in1(N__48416),
            .in2(N__50547),
            .in3(N__43280),
            .lcout(\c0.data_out_3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49844),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i25_LC_15_19_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i25_LC_15_19_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i25_LC_15_19_0 .LUT_INIT=16'b1110000011000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i25_LC_15_19_0  (
            .in0(N__45030),
            .in1(N__44737),
            .in2(N__43266),
            .in3(N__44605),
            .lcout(\c0.FRAME_MATCHER_state_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49749),
            .ce(),
            .sr(N__43242));
    defparam \c0.FRAME_MATCHER_state_i26_LC_15_20_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i26_LC_15_20_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i26_LC_15_20_0 .LUT_INIT=16'b1100110010000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i26_LC_15_20_0  (
            .in0(N__45029),
            .in1(N__43225),
            .in2(N__44604),
            .in3(N__44738),
            .lcout(\c0.FRAME_MATCHER_state_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49761),
            .ce(),
            .sr(N__43203));
    defparam \c0.FRAME_MATCHER_state_i15_LC_15_21_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i15_LC_15_21_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i15_LC_15_21_0 .LUT_INIT=16'b1110000011000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i15_LC_15_21_0  (
            .in0(N__45018),
            .in1(N__44702),
            .in2(N__43190),
            .in3(N__44573),
            .lcout(\c0.FRAME_MATCHER_state_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49774),
            .ce(),
            .sr(N__43164));
    defparam \c0.FRAME_MATCHER_state_i21_LC_15_22_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i21_LC_15_22_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i21_LC_15_22_0 .LUT_INIT=16'b1110000011000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i21_LC_15_22_0  (
            .in0(N__44976),
            .in1(N__44678),
            .in2(N__43157),
            .in3(N__44511),
            .lcout(\c0.FRAME_MATCHER_state_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49786),
            .ce(),
            .sr(N__43131));
    defparam \c0.FRAME_MATCHER_state_i24_LC_15_23_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i24_LC_15_23_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i24_LC_15_23_0 .LUT_INIT=16'b1110000011000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i24_LC_15_23_0  (
            .in0(N__45028),
            .in1(N__44675),
            .in2(N__43114),
            .in3(N__44583),
            .lcout(\c0.FRAME_MATCHER_state_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49796),
            .ce(),
            .sr(N__43089));
    defparam \c0.data_out_10__4__2172_LC_15_25_1 .C_ON=1'b0;
    defparam \c0.data_out_10__4__2172_LC_15_25_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_10__4__2172_LC_15_25_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_out_10__4__2172_LC_15_25_1  (
            .in0(N__43415),
            .in1(N__46726),
            .in2(_gnd_net_),
            .in3(N__47265),
            .lcout(\c0.data_out_10_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49813),
            .ce(N__49980),
            .sr(_gnd_net_));
    defparam \c0.i3_4_lut_adj_421_LC_15_25_2 .C_ON=1'b0;
    defparam \c0.i3_4_lut_adj_421_LC_15_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.i3_4_lut_adj_421_LC_15_25_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i3_4_lut_adj_421_LC_15_25_2  (
            .in0(N__43406),
            .in1(N__47132),
            .in2(N__45843),
            .in3(N__45420),
            .lcout(\c0.n17201 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_9__7__2177_LC_15_25_3 .C_ON=1'b0;
    defparam \c0.data_out_9__7__2177_LC_15_25_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_9__7__2177_LC_15_25_3 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_9__7__2177_LC_15_25_3  (
            .in0(N__43416),
            .in1(N__43491),
            .in2(N__43485),
            .in3(N__47277),
            .lcout(\c0.data_out_9_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49813),
            .ce(N__49980),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_435_LC_15_25_5 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_435_LC_15_25_5 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_435_LC_15_25_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_435_LC_15_25_5  (
            .in0(_gnd_net_),
            .in1(N__47536),
            .in2(_gnd_net_),
            .in3(N__43470),
            .lcout(\c0.n10316 ),
            .ltout(\c0.n10316_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_9__4__2180_LC_15_25_6 .C_ON=1'b0;
    defparam \c0.data_out_9__4__2180_LC_15_25_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_9__4__2180_LC_15_25_6 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_9__4__2180_LC_15_25_6  (
            .in0(N__43425),
            .in1(N__43551),
            .in2(N__43419),
            .in3(N__45743),
            .lcout(\c0.data_out_9_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49813),
            .ce(N__49980),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_731_LC_15_26_0 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_731_LC_15_26_0 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_731_LC_15_26_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_731_LC_15_26_0  (
            .in0(N__47038),
            .in1(N__46825),
            .in2(N__47199),
            .in3(N__47014),
            .lcout(\c0.n17177 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i8_3_lut_LC_15_26_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i8_3_lut_LC_15_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i8_3_lut_LC_15_26_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_6_i8_3_lut_LC_15_26_1  (
            .in0(N__43399),
            .in1(N__45435),
            .in2(_gnd_net_),
            .in3(N__47791),
            .lcout(\c0.n8_adj_2157 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_3_lut_adj_694_LC_15_26_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_3_lut_adj_694_LC_15_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_3_lut_adj_694_LC_15_26_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i1_2_lut_3_lut_adj_694_LC_15_26_2  (
            .in0(N__43359),
            .in1(N__43398),
            .in2(_gnd_net_),
            .in3(N__45614),
            .lcout(\c0.n26_adj_2165 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9952_3_lut_LC_15_26_3 .C_ON=1'b0;
    defparam \c0.i9952_3_lut_LC_15_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.i9952_3_lut_LC_15_26_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.i9952_3_lut_LC_15_26_3  (
            .in0(N__43549),
            .in1(N__43358),
            .in2(_gnd_net_),
            .in3(N__47487),
            .lcout(\c0.n12630 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_471_LC_15_26_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_471_LC_15_26_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_471_LC_15_26_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_471_LC_15_26_4  (
            .in0(N__43320),
            .in1(N__47264),
            .in2(_gnd_net_),
            .in3(N__43624),
            .lcout(\c0.n10179 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__1__2255_LC_15_26_5 .C_ON=1'b0;
    defparam \c0.data_out_0__1__2255_LC_15_26_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__1__2255_LC_15_26_5 .LUT_INIT=16'b0111011101000100;
    LogicCell40 \c0.data_out_0__1__2255_LC_15_26_5  (
            .in0(N__50262),
            .in1(N__50537),
            .in2(_gnd_net_),
            .in3(N__43575),
            .lcout(data_out_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49821),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_8__5__2187_LC_15_26_6 .C_ON=1'b0;
    defparam \c0.data_out_8__5__2187_LC_15_26_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_8__5__2187_LC_15_26_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.data_out_8__5__2187_LC_15_26_6  (
            .in0(N__49977),
            .in1(N__43743),
            .in2(_gnd_net_),
            .in3(N__45615),
            .lcout(data_out_8_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49821),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_7__5__2195_LC_15_26_7 .C_ON=1'b0;
    defparam \c0.data_out_7__5__2195_LC_15_26_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_7__5__2195_LC_15_26_7 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \c0.data_out_7__5__2195_LC_15_26_7  (
            .in0(N__43625),
            .in1(N__43717),
            .in2(N__43650),
            .in3(N__46898),
            .lcout(\c0.data_out_7_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49821),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i7_LC_15_27_0 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i7_LC_15_27_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i7_LC_15_27_0 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \c0.tx.r_Tx_Data_i7_LC_15_27_0  (
            .in0(N__46176),
            .in1(N__43601),
            .in2(N__44098),
            .in3(N__43844),
            .lcout(r_Tx_Data_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49828),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_1_i1_3_lut_LC_15_27_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_1_i1_3_lut_LC_15_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_1_i1_3_lut_LC_15_27_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_1_i1_3_lut_LC_15_27_2  (
            .in0(N__43587),
            .in1(N__43574),
            .in2(_gnd_net_),
            .in3(N__47803),
            .lcout(n1_adj_2449),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9953_4_lut_LC_15_27_3 .C_ON=1'b0;
    defparam \c0.i9953_4_lut_LC_15_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.i9953_4_lut_LC_15_27_3 .LUT_INIT=16'b1101100010001000;
    LogicCell40 \c0.i9953_4_lut_LC_15_27_3  (
            .in0(N__47804),
            .in1(N__43557),
            .in2(N__46832),
            .in3(N__47495),
            .lcout(n6_adj_2446),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_453_LC_15_27_4 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_453_LC_15_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_453_LC_15_27_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_453_LC_15_27_4  (
            .in0(N__43550),
            .in1(N__45590),
            .in2(N__45464),
            .in3(N__43529),
            .lcout(),
            .ltout(\c0.n10_adj_2189_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_454_LC_15_27_5 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_454_LC_15_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_454_LC_15_27_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.i5_3_lut_adj_454_LC_15_27_5  (
            .in0(N__49033),
            .in1(_gnd_net_),
            .in2(N__43518),
            .in3(N__48896),
            .lcout(data_out_9__2__N_367),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i0_LC_15_27_6 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i0_LC_15_27_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i0_LC_15_27_6 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \c0.tx.r_Tx_Data_i0_LC_15_27_6  (
            .in0(N__43511),
            .in1(N__45750),
            .in2(N__44097),
            .in3(N__43843),
            .lcout(r_Tx_Data_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49828),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i10_4_lut_LC_15_27_7 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i10_4_lut_LC_15_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_6_i10_4_lut_LC_15_27_7 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_6_i10_4_lut_LC_15_27_7  (
            .in0(N__47805),
            .in1(N__43497),
            .in2(N__49040),
            .in3(N__47496),
            .lcout(n10_adj_2422),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i5_3_lut_LC_15_28_0 .C_ON=1'b0;
    defparam \c0.tx.i5_3_lut_LC_15_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i5_3_lut_LC_15_28_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \c0.tx.i5_3_lut_LC_15_28_0  (
            .in0(N__46051),
            .in1(N__45784),
            .in2(_gnd_net_),
            .in3(N__43851),
            .lcout(),
            .ltout(\c0.tx.n77_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i101_4_lut_LC_15_28_1 .C_ON=1'b0;
    defparam \c0.tx.i101_4_lut_LC_15_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i101_4_lut_LC_15_28_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \c0.tx.i101_4_lut_LC_15_28_1  (
            .in0(N__45990),
            .in1(N__46021),
            .in2(N__43899),
            .in3(N__46546),
            .lcout(\c0.tx.n83 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i3_LC_15_28_2 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i3_LC_15_28_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i3_LC_15_28_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.tx.r_Clock_Count__i3_LC_15_28_2  (
            .in0(_gnd_net_),
            .in1(N__45522),
            .in2(_gnd_net_),
            .in3(N__46123),
            .lcout(\c0.tx.r_Clock_Count_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49834),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.o_Tx_Serial_45_LC_15_28_3 .C_ON=1'b0;
    defparam \c0.tx.o_Tx_Serial_45_LC_15_28_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.o_Tx_Serial_45_LC_15_28_3 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \c0.tx.o_Tx_Serial_45_LC_15_28_3  (
            .in0(N__45945),
            .in1(N__43862),
            .in2(_gnd_net_),
            .in3(N__43896),
            .lcout(tx_o),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49834),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i4_4_lut_LC_15_28_4 .C_ON=1'b0;
    defparam \c0.tx.i4_4_lut_LC_15_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i4_4_lut_LC_15_28_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \c0.tx.i4_4_lut_LC_15_28_4  (
            .in0(N__46153),
            .in1(N__46084),
            .in2(N__45543),
            .in3(N__45568),
            .lcout(\c0.tx.n10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i6_LC_15_28_5 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i6_LC_15_28_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i6_LC_15_28_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \c0.tx.r_Clock_Count__i6_LC_15_28_5  (
            .in0(N__46125),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46005),
            .lcout(\c0.tx.r_Clock_Count_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49834),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Data_i6_LC_15_28_6 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Data_i6_LC_15_28_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Data_i6_LC_15_28_6 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \c0.tx.r_Tx_Data_i6_LC_15_28_6  (
            .in0(N__43840),
            .in1(N__43764),
            .in2(N__44075),
            .in3(N__43757),
            .lcout(r_Tx_Data_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49834),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i5_LC_15_28_7 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i5_LC_15_28_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i5_LC_15_28_7 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \c0.tx.r_Clock_Count__i5_LC_15_28_7  (
            .in0(N__46124),
            .in1(_gnd_net_),
            .in2(N__46035),
            .in3(_gnd_net_),
            .lcout(\c0.tx.r_Clock_Count_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49834),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_2_lut_adj_402_LC_15_29_1 .C_ON=1'b0;
    defparam \c0.tx.i1_2_lut_adj_402_LC_15_29_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_2_lut_adj_402_LC_15_29_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.tx.i1_2_lut_adj_402_LC_15_29_1  (
            .in0(_gnd_net_),
            .in1(N__43986),
            .in2(_gnd_net_),
            .in3(N__43936),
            .lcout(\c0.tx.n13702 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_i0_LC_15_29_2 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_i0_LC_15_29_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_SM_Main_i0_LC_15_29_2 .LUT_INIT=16'b0001001100010000;
    LogicCell40 \c0.tx.r_SM_Main_i0_LC_15_29_2  (
            .in0(N__43937),
            .in1(N__45941),
            .in2(N__44004),
            .in3(N__44115),
            .lcout(\c0.tx.r_SM_Main_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49837),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i2_LC_15_29_3 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i2_LC_15_29_3 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i2_LC_15_29_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.tx.r_Clock_Count__i2_LC_15_29_3  (
            .in0(_gnd_net_),
            .in1(N__45552),
            .in2(_gnd_net_),
            .in3(N__46111),
            .lcout(\c0.tx.r_Clock_Count_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49837),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i8_3_lut_LC_15_29_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i8_3_lut_LC_15_29_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i8_3_lut_LC_15_29_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_7_i8_3_lut_LC_15_29_4  (
            .in0(N__46627),
            .in1(N__45838),
            .in2(_gnd_net_),
            .in3(N__47833),
            .lcout(),
            .ltout(\c0.n8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i10_4_lut_LC_15_29_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i10_4_lut_LC_15_29_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i10_4_lut_LC_15_29_5 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_7_i10_4_lut_LC_15_29_5  (
            .in0(N__47834),
            .in1(N__48446),
            .in2(N__44109),
            .in3(N__47494),
            .lcout(n10_adj_2413),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_2_lut_3_lut_4_lut_LC_15_29_6 .C_ON=1'b0;
    defparam \c0.tx.i1_2_lut_3_lut_4_lut_LC_15_29_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_2_lut_3_lut_4_lut_LC_15_29_6 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \c0.tx.i1_2_lut_3_lut_4_lut_LC_15_29_6  (
            .in0(N__50819),
            .in1(N__44178),
            .in2(N__44003),
            .in3(N__45940),
            .lcout(n9257),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_2_lut_LC_15_29_7 .C_ON=1'b0;
    defparam \c0.tx.i1_2_lut_LC_15_29_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_2_lut_LC_15_29_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \c0.tx.i1_2_lut_LC_15_29_7  (
            .in0(_gnd_net_),
            .in1(N__43985),
            .in2(_gnd_net_),
            .in3(N__50818),
            .lcout(\c0.tx.n6759 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_SM_Main_i1_LC_15_30_0 .C_ON=1'b0;
    defparam \c0.tx.r_SM_Main_i1_LC_15_30_0 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_SM_Main_i1_LC_15_30_0 .LUT_INIT=16'b0001001000110000;
    LogicCell40 \c0.tx.r_SM_Main_i1_LC_15_30_0  (
            .in0(N__43999),
            .in1(N__45926),
            .in2(N__44193),
            .in3(N__43952),
            .lcout(\c0.tx.r_SM_Main_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49840),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_2_lut_adj_401_LC_15_30_1 .C_ON=1'b0;
    defparam \c0.tx.i1_2_lut_adj_401_LC_15_30_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_2_lut_adj_401_LC_15_30_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.tx.i1_2_lut_adj_401_LC_15_30_1  (
            .in0(_gnd_net_),
            .in1(N__44295),
            .in2(_gnd_net_),
            .in3(N__50762),
            .lcout(\c0.n65_adj_2192 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_3_lut_4_lut_4_lut_LC_15_30_4 .C_ON=1'b0;
    defparam \c0.tx.i1_3_lut_4_lut_4_lut_LC_15_30_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_3_lut_4_lut_4_lut_LC_15_30_4 .LUT_INIT=16'b0011001100000001;
    LogicCell40 \c0.tx.i1_3_lut_4_lut_4_lut_LC_15_30_4  (
            .in0(N__43998),
            .in1(N__45924),
            .in2(N__44191),
            .in3(N__43951),
            .lcout(n5142),
            .ltout(n5142_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i8_LC_15_30_5 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i8_LC_15_30_5 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i8_LC_15_30_5 .LUT_INIT=16'b0000110000001100;
    LogicCell40 \c0.tx.r_Clock_Count__i8_LC_15_30_5  (
            .in0(_gnd_net_),
            .in1(N__45849),
            .in2(N__44313),
            .in3(_gnd_net_),
            .lcout(\c0.tx.r_Clock_Count_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49840),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_4_lut_adj_399_LC_15_30_6 .C_ON=1'b0;
    defparam \c0.tx.i1_4_lut_adj_399_LC_15_30_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_4_lut_adj_399_LC_15_30_6 .LUT_INIT=16'b0000000011001010;
    LogicCell40 \c0.tx.i1_4_lut_adj_399_LC_15_30_6  (
            .in0(N__44310),
            .in1(N__44301),
            .in2(N__44192),
            .in3(N__45925),
            .lcout(\c0.tx.n10613 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx_active_prev_2167_LC_15_30_7 .C_ON=1'b0;
    defparam \c0.tx_active_prev_2167_LC_15_30_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx_active_prev_2167_LC_15_30_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \c0.tx_active_prev_2167_LC_15_30_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50763),
            .lcout(\c0.tx_active_prev ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49840),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15104_2_lut_LC_15_31_0 .C_ON=1'b0;
    defparam \c0.i15104_2_lut_LC_15_31_0 .SEQ_MODE=4'b0000;
    defparam \c0.i15104_2_lut_LC_15_31_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \c0.i15104_2_lut_LC_15_31_0  (
            .in0(N__47826),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44289),
            .lcout(),
            .ltout(\c0.n17581_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15361_LC_15_31_1 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15361_LC_15_31_1 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15361_LC_15_31_1 .LUT_INIT=16'b1011101111000000;
    LogicCell40 \c0.byte_transmit_counter_1__bdd_4_lut_15361_LC_15_31_1  (
            .in0(N__44238),
            .in1(N__46299),
            .in2(N__44226),
            .in3(N__47507),
            .lcout(\c0.n18088 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_3__7__2225_LC_15_31_4 .C_ON=1'b0;
    defparam \c0.data_out_3__7__2225_LC_15_31_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_3__7__2225_LC_15_31_4 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \c0.data_out_3__7__2225_LC_15_31_4  (
            .in0(N__48112),
            .in1(N__50317),
            .in2(N__50529),
            .in3(N__46530),
            .lcout(data_out_3_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49845),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i10_4_lut_LC_15_31_5 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i10_4_lut_LC_15_31_5 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i10_4_lut_LC_15_31_5 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_5_i10_4_lut_LC_15_31_5  (
            .in0(N__44325),
            .in1(N__47508),
            .in2(N__48687),
            .in3(N__47827),
            .lcout(n10_adj_2432),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Tx_Active_47_LC_15_31_6 .C_ON=1'b0;
    defparam \c0.tx.r_Tx_Active_47_LC_15_31_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Tx_Active_47_LC_15_31_6 .LUT_INIT=16'b0111010001110100;
    LogicCell40 \c0.tx.r_Tx_Active_47_LC_15_31_6  (
            .in0(N__44180),
            .in1(N__44121),
            .in2(N__50781),
            .in3(_gnd_net_),
            .lcout(\c0.tx_active ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49845),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i2_3_lut_LC_15_32_2 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i2_3_lut_LC_15_32_2 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i2_3_lut_LC_15_32_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_5_i2_3_lut_LC_15_32_2  (
            .in0(N__45323),
            .in1(N__50007),
            .in2(_gnd_net_),
            .in3(N__47828),
            .lcout(),
            .ltout(\c0.n2_adj_2164_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18088_bdd_4_lut_LC_15_32_3 .C_ON=1'b0;
    defparam \c0.n18088_bdd_4_lut_LC_15_32_3 .SEQ_MODE=4'b0000;
    defparam \c0.n18088_bdd_4_lut_LC_15_32_3 .LUT_INIT=16'b1100110011100010;
    LogicCell40 \c0.n18088_bdd_4_lut_LC_15_32_3  (
            .in0(N__45354),
            .in1(N__45339),
            .in2(N__45333),
            .in3(N__46321),
            .lcout(n18091),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_3__5__2227_LC_15_32_4 .C_ON=1'b0;
    defparam \c0.data_out_3__5__2227_LC_15_32_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_3__5__2227_LC_15_32_4 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \c0.data_out_3__5__2227_LC_15_32_4  (
            .in0(N__45324),
            .in1(N__48113),
            .in2(N__50333),
            .in3(N__50418),
            .lcout(data_out_3_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49848),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_0__6__2250_LC_15_32_7 .C_ON=1'b0;
    defparam \c0.data_out_0__6__2250_LC_15_32_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_0__6__2250_LC_15_32_7 .LUT_INIT=16'b0001111100010000;
    LogicCell40 \c0.data_out_0__6__2250_LC_15_32_7  (
            .in0(N__48383),
            .in1(N__50324),
            .in2(N__50471),
            .in3(N__45308),
            .lcout(\c0.data_out_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49848),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.rx.r_Rx_Byte_i4_LC_16_20_4 .C_ON=1'b0;
    defparam \c0.rx.r_Rx_Byte_i4_LC_16_20_4 .SEQ_MODE=4'b1000;
    defparam \c0.rx.r_Rx_Byte_i4_LC_16_20_4 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \c0.rx.r_Rx_Byte_i4_LC_16_20_4  (
            .in0(N__45293),
            .in1(N__45259),
            .in2(N__45097),
            .in3(N__45176),
            .lcout(rx_data_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49775),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_1__6__2242_LC_16_22_5 .C_ON=1'b0;
    defparam \c0.data_out_1__6__2242_LC_16_22_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_1__6__2242_LC_16_22_5 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \c0.data_out_1__6__2242_LC_16_22_5  (
            .in0(N__48168),
            .in1(N__50291),
            .in2(N__50583),
            .in3(N__45050),
            .lcout(data_out_1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49797),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.FRAME_MATCHER_state_i22_LC_16_24_0 .C_ON=1'b0;
    defparam \c0.FRAME_MATCHER_state_i22_LC_16_24_0 .SEQ_MODE=4'b1001;
    defparam \c0.FRAME_MATCHER_state_i22_LC_16_24_0 .LUT_INIT=16'b1110000011000000;
    LogicCell40 \c0.FRAME_MATCHER_state_i22_LC_16_24_0  (
            .in0(N__45031),
            .in1(N__44724),
            .in2(N__44371),
            .in3(N__44617),
            .lcout(\c0.FRAME_MATCHER_state_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49814),
            .ce(),
            .sr(N__44349));
    defparam \c0.data_out_1__7__2241_LC_16_25_1 .C_ON=1'b0;
    defparam \c0.data_out_1__7__2241_LC_16_25_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_1__7__2241_LC_16_25_1 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \c0.data_out_1__7__2241_LC_16_25_1  (
            .in0(N__50533),
            .in1(N__50292),
            .in2(_gnd_net_),
            .in3(N__44334),
            .lcout(data_out_1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49822),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15018_2_lut_LC_16_25_3 .C_ON=1'b0;
    defparam \c0.i15018_2_lut_LC_16_25_3 .SEQ_MODE=4'b0000;
    defparam \c0.i15018_2_lut_LC_16_25_3 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \c0.i15018_2_lut_LC_16_25_3  (
            .in0(N__47839),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44333),
            .lcout(\c0.n17607 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i8_3_lut_LC_16_25_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i8_3_lut_LC_16_25_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_5_i8_3_lut_LC_16_25_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_5_i8_3_lut_LC_16_25_4  (
            .in0(N__48533),
            .in1(N__45616),
            .in2(_gnd_net_),
            .in3(N__47838),
            .lcout(\c0.n8_adj_2352 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_10__2__2174_LC_16_26_0 .C_ON=1'b0;
    defparam \c0.data_out_10__2__2174_LC_16_26_0 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_10__2__2174_LC_16_26_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_10__2__2174_LC_16_26_0  (
            .in0(N__45434),
            .in1(N__45509),
            .in2(N__46965),
            .in3(N__49168),
            .lcout(\c0.data_out_10_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49829),
            .ce(N__49988),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_497_LC_16_26_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_497_LC_16_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_497_LC_16_26_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_497_LC_16_26_1  (
            .in0(_gnd_net_),
            .in1(N__45433),
            .in2(_gnd_net_),
            .in3(N__45656),
            .lcout(\c0.n17209 ),
            .ltout(\c0.n17209_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_10__6__2170_LC_16_26_2 .C_ON=1'b0;
    defparam \c0.data_out_10__6__2170_LC_16_26_2 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_10__6__2170_LC_16_26_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_10__6__2170_LC_16_26_2  (
            .in0(N__45441),
            .in1(N__45494),
            .in2(N__45468),
            .in3(N__47015),
            .lcout(\c0.data_out_10_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49829),
            .ce(N__49988),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_501_LC_16_26_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_501_LC_16_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_501_LC_16_26_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_501_LC_16_26_3  (
            .in0(_gnd_net_),
            .in1(N__45414),
            .in2(_gnd_net_),
            .in3(N__45463),
            .lcout(\c0.n6_adj_2216 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_9__6__2178_LC_16_26_4 .C_ON=1'b0;
    defparam \c0.data_out_9__6__2178_LC_16_26_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_9__6__2178_LC_16_26_4 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \c0.data_out_9__6__2178_LC_16_26_4  (
            .in0(N__48616),
            .in1(N__46574),
            .in2(N__48948),
            .in3(N__48572),
            .lcout(\c0.data_out_9_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49829),
            .ce(N__49988),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_425_LC_16_26_7 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_425_LC_16_26_7 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_425_LC_16_26_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_425_LC_16_26_7  (
            .in0(N__48571),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48615),
            .lcout(\c0.n17200 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i51_4_lut_LC_16_27_0.C_ON=1'b0;
    defparam i51_4_lut_LC_16_27_0.SEQ_MODE=4'b0000;
    defparam i51_4_lut_LC_16_27_0.LUT_INIT=16'b0101000011001100;
    LogicCell40 i51_4_lut_LC_16_27_0 (
            .in0(N__47832),
            .in1(N__45378),
            .in2(N__47195),
            .in3(N__47513),
            .lcout(n32),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i9896_3_lut_LC_16_27_1 .C_ON=1'b0;
    defparam \c0.i9896_3_lut_LC_16_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.i9896_3_lut_LC_16_27_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \c0.i9896_3_lut_LC_16_27_1  (
            .in0(N__45413),
            .in1(N__48614),
            .in2(_gnd_net_),
            .in3(N__47831),
            .lcout(n8_adj_2445),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i52_3_lut_LC_16_27_2.C_ON=1'b0;
    defparam i52_3_lut_LC_16_27_2.SEQ_MODE=4'b0000;
    defparam i52_3_lut_LC_16_27_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 i52_3_lut_LC_16_27_2 (
            .in0(N__45372),
            .in1(N__45366),
            .in2(_gnd_net_),
            .in3(N__46322),
            .lcout(),
            .ltout(n29_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i49_4_lut_LC_16_27_3.C_ON=1'b0;
    defparam i49_4_lut_LC_16_27_3.SEQ_MODE=4'b0000;
    defparam i49_4_lut_LC_16_27_3.LUT_INIT=16'b0100010011110000;
    LogicCell40 i49_4_lut_LC_16_27_3 (
            .in0(N__46323),
            .in1(N__45759),
            .in2(N__45753),
            .in3(N__46415),
            .lcout(n26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_742_LC_16_27_4 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_742_LC_16_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_742_LC_16_27_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_742_LC_16_27_4  (
            .in0(N__48659),
            .in1(N__48926),
            .in2(N__48620),
            .in3(N__45744),
            .lcout(\c0.n10196 ),
            .ltout(\c0.n10196_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_448_LC_16_27_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_448_LC_16_27_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_448_LC_16_27_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i2_3_lut_adj_448_LC_16_27_5  (
            .in0(_gnd_net_),
            .in1(N__48447),
            .in2(N__45681),
            .in3(N__45678),
            .lcout(\c0.n17243 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_9__0__2184_LC_16_27_6 .C_ON=1'b0;
    defparam \c0.data_out_9__0__2184_LC_16_27_6 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_9__0__2184_LC_16_27_6 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_9__0__2184_LC_16_27_6  (
            .in0(N__45657),
            .in1(N__45621),
            .in2(N__46662),
            .in3(N__45591),
            .lcout(\c0.data_out_9_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49835),
            .ce(N__49979),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_2_lut_LC_16_28_0 .C_ON=1'b1;
    defparam \c0.tx.add_59_2_lut_LC_16_28_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_2_lut_LC_16_28_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.tx.add_59_2_lut_LC_16_28_0  (
            .in0(N__46086),
            .in1(N__46085),
            .in2(N__45958),
            .in3(N__45576),
            .lcout(n10994),
            .ltout(),
            .carryin(bfn_16_28_0_),
            .carryout(\c0.tx.n16117 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_3_lut_LC_16_28_1 .C_ON=1'b1;
    defparam \c0.tx.add_59_3_lut_LC_16_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_3_lut_LC_16_28_1 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.tx.add_59_3_lut_LC_16_28_1  (
            .in0(N__45786),
            .in1(N__45785),
            .in2(N__45963),
            .in3(N__45573),
            .lcout(n10951),
            .ltout(),
            .carryin(\c0.tx.n16117 ),
            .carryout(\c0.tx.n16118 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_4_lut_LC_16_28_2 .C_ON=1'b1;
    defparam \c0.tx.add_59_4_lut_LC_16_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_4_lut_LC_16_28_2 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.tx.add_59_4_lut_LC_16_28_2  (
            .in0(N__45570),
            .in1(N__45569),
            .in2(N__45959),
            .in3(N__45546),
            .lcout(n10954),
            .ltout(),
            .carryin(\c0.tx.n16118 ),
            .carryout(\c0.tx.n16119 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_5_lut_LC_16_28_3 .C_ON=1'b1;
    defparam \c0.tx.add_59_5_lut_LC_16_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_5_lut_LC_16_28_3 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.tx.add_59_5_lut_LC_16_28_3  (
            .in0(N__45542),
            .in1(N__45541),
            .in2(N__45964),
            .in3(N__45516),
            .lcout(n10957),
            .ltout(),
            .carryin(\c0.tx.n16119 ),
            .carryout(\c0.tx.n16120 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_6_lut_LC_16_28_4 .C_ON=1'b1;
    defparam \c0.tx.add_59_6_lut_LC_16_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_6_lut_LC_16_28_4 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.tx.add_59_6_lut_LC_16_28_4  (
            .in0(N__46155),
            .in1(N__46154),
            .in2(N__45960),
            .in3(N__46059),
            .lcout(n10960),
            .ltout(),
            .carryin(\c0.tx.n16120 ),
            .carryout(\c0.tx.n16121 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_7_lut_LC_16_28_5 .C_ON=1'b1;
    defparam \c0.tx.add_59_7_lut_LC_16_28_5 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_7_lut_LC_16_28_5 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.tx.add_59_7_lut_LC_16_28_5  (
            .in0(N__46055),
            .in1(N__46056),
            .in2(N__45965),
            .in3(N__46026),
            .lcout(n10963),
            .ltout(),
            .carryin(\c0.tx.n16121 ),
            .carryout(\c0.tx.n16122 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_8_lut_LC_16_28_6 .C_ON=1'b1;
    defparam \c0.tx.add_59_8_lut_LC_16_28_6 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_8_lut_LC_16_28_6 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.tx.add_59_8_lut_LC_16_28_6  (
            .in0(N__46023),
            .in1(N__46022),
            .in2(N__45961),
            .in3(N__45996),
            .lcout(n10966),
            .ltout(),
            .carryin(\c0.tx.n16122 ),
            .carryout(\c0.tx.n16123 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_9_lut_LC_16_28_7 .C_ON=1'b1;
    defparam \c0.tx.add_59_9_lut_LC_16_28_7 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_9_lut_LC_16_28_7 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.tx.add_59_9_lut_LC_16_28_7  (
            .in0(N__46551),
            .in1(N__46547),
            .in2(N__45966),
            .in3(N__45993),
            .lcout(n10969),
            .ltout(),
            .carryin(\c0.tx.n16123 ),
            .carryout(\c0.tx.n16124 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.add_59_10_lut_LC_16_29_0 .C_ON=1'b0;
    defparam \c0.tx.add_59_10_lut_LC_16_29_0 .SEQ_MODE=4'b0000;
    defparam \c0.tx.add_59_10_lut_LC_16_29_0 .LUT_INIT=16'b1010001110101100;
    LogicCell40 \c0.tx.add_59_10_lut_LC_16_29_0  (
            .in0(N__45985),
            .in1(N__45986),
            .in2(N__45962),
            .in3(N__45852),
            .lcout(n10972),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_468_LC_16_29_2 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_468_LC_16_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_468_LC_16_29_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_468_LC_16_29_2  (
            .in0(N__46833),
            .in1(N__48971),
            .in2(_gnd_net_),
            .in3(N__47322),
            .lcout(\c0.n17197 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_423_LC_16_29_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_423_LC_16_29_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_423_LC_16_29_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_423_LC_16_29_3  (
            .in0(_gnd_net_),
            .in1(N__48683),
            .in2(_gnd_net_),
            .in3(N__45839),
            .lcout(\c0.n6_adj_2169 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i1_LC_16_29_6 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i1_LC_16_29_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i1_LC_16_29_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.tx.r_Clock_Count__i1_LC_16_29_6  (
            .in0(_gnd_net_),
            .in1(N__45792),
            .in2(_gnd_net_),
            .in3(N__46121),
            .lcout(\c0.tx.r_Clock_Count_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49841),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i7_LC_16_29_7 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i7_LC_16_29_7 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i7_LC_16_29_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \c0.tx.r_Clock_Count__i7_LC_16_29_7  (
            .in0(N__46122),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45768),
            .lcout(\c0.tx.r_Clock_Count_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49841),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i2_3_lut_LC_16_30_0 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i2_3_lut_LC_16_30_0 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_7_i2_3_lut_LC_16_30_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_7_i2_3_lut_LC_16_30_0  (
            .in0(N__47829),
            .in1(N__46529),
            .in2(_gnd_net_),
            .in3(N__46517),
            .lcout(\c0.n2_adj_2156 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_2__7__2233_LC_16_30_1 .C_ON=1'b0;
    defparam \c0.data_out_2__7__2233_LC_16_30_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_2__7__2233_LC_16_30_1 .LUT_INIT=16'b0000101011111010;
    LogicCell40 \c0.data_out_2__7__2233_LC_16_30_1  (
            .in0(N__46518),
            .in1(_gnd_net_),
            .in2(N__50470),
            .in3(N__50244),
            .lcout(data_out_2_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49846),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15148_2_lut_LC_16_30_3 .C_ON=1'b0;
    defparam \c0.i15148_2_lut_LC_16_30_3 .SEQ_MODE=4'b0000;
    defparam \c0.i15148_2_lut_LC_16_30_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \c0.i15148_2_lut_LC_16_30_3  (
            .in0(_gnd_net_),
            .in1(N__46508),
            .in2(_gnd_net_),
            .in3(N__47830),
            .lcout(),
            .ltout(\c0.n17747_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15445_LC_16_30_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15445_LC_16_30_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_1__bdd_4_lut_15445_LC_16_30_4 .LUT_INIT=16'b1011101111000000;
    LogicCell40 \c0.byte_transmit_counter_1__bdd_4_lut_15445_LC_16_30_4  (
            .in0(N__46449),
            .in1(N__46313),
            .in2(N__46437),
            .in3(N__47509),
            .lcout(),
            .ltout(\c0.n18220_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.n18220_bdd_4_lut_LC_16_30_5 .C_ON=1'b0;
    defparam \c0.n18220_bdd_4_lut_LC_16_30_5 .SEQ_MODE=4'b0000;
    defparam \c0.n18220_bdd_4_lut_LC_16_30_5 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \c0.n18220_bdd_4_lut_LC_16_30_5  (
            .in0(N__46314),
            .in1(N__46434),
            .in2(N__46428),
            .in3(N__46425),
            .lcout(),
            .ltout(n18223_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_4_lut_LC_16_30_6.C_ON=1'b0;
    defparam i24_4_lut_LC_16_30_6.SEQ_MODE=4'b0000;
    defparam i24_4_lut_LC_16_30_6.LUT_INIT=16'b0101000011011000;
    LogicCell40 i24_4_lut_LC_16_30_6 (
            .in0(N__46416),
            .in1(N__46332),
            .in2(N__46326),
            .in3(N__46315),
            .lcout(n10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i4_LC_16_31_2 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i4_LC_16_31_2 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i4_LC_16_31_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.tx.r_Clock_Count__i4_LC_16_31_2  (
            .in0(_gnd_net_),
            .in1(N__46164),
            .in2(_gnd_net_),
            .in3(N__46120),
            .lcout(\c0.tx.r_Clock_Count_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49849),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.tx.r_Clock_Count__i0_LC_16_31_6 .C_ON=1'b0;
    defparam \c0.tx.r_Clock_Count__i0_LC_16_31_6 .SEQ_MODE=4'b1000;
    defparam \c0.tx.r_Clock_Count__i0_LC_16_31_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \c0.tx.r_Clock_Count__i0_LC_16_31_6  (
            .in0(_gnd_net_),
            .in1(N__46134),
            .in2(_gnd_net_),
            .in3(N__46119),
            .lcout(\c0.tx.r_Clock_Count_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49849),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15208_4_lut_2_lut_3_lut_LC_16_31_7 .C_ON=1'b0;
    defparam \c0.i15208_4_lut_2_lut_3_lut_LC_16_31_7 .SEQ_MODE=4'b0000;
    defparam \c0.i15208_4_lut_2_lut_3_lut_LC_16_31_7 .LUT_INIT=16'b0100010011001100;
    LogicCell40 \c0.i15208_4_lut_2_lut_3_lut_LC_16_31_7  (
            .in0(N__48372),
            .in1(N__48111),
            .in2(_gnd_net_),
            .in3(N__50236),
            .lcout(n10596),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i15202_2_lut_3_lut_LC_16_32_1 .C_ON=1'b0;
    defparam \c0.i15202_2_lut_3_lut_LC_16_32_1 .SEQ_MODE=4'b0000;
    defparam \c0.i15202_2_lut_3_lut_LC_16_32_1 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \c0.i15202_2_lut_3_lut_LC_16_32_1  (
            .in0(N__50390),
            .in1(N__48382),
            .in2(_gnd_net_),
            .in3(N__50237),
            .lcout(\c0.n10595 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_727_LC_17_25_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_727_LC_17_25_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_727_LC_17_25_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_727_LC_17_25_2  (
            .in0(N__46704),
            .in1(N__48534),
            .in2(N__46734),
            .in3(N__46766),
            .lcout(\c0.n17252 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_479_LC_17_26_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_479_LC_17_26_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_479_LC_17_26_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_479_LC_17_26_1  (
            .in0(_gnd_net_),
            .in1(N__46824),
            .in2(_gnd_net_),
            .in3(N__47016),
            .lcout(),
            .ltout(\c0.n10447_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_4_lut_adj_440_LC_17_26_2 .C_ON=1'b0;
    defparam \c0.i5_4_lut_adj_440_LC_17_26_2 .SEQ_MODE=4'b0000;
    defparam \c0.i5_4_lut_adj_440_LC_17_26_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i5_4_lut_adj_440_LC_17_26_2  (
            .in0(N__46788),
            .in1(N__48770),
            .in2(N__46773),
            .in3(N__49014),
            .lcout(\c0.n12_adj_2180 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_490_LC_17_26_3 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_490_LC_17_26_3 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_490_LC_17_26_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_490_LC_17_26_3  (
            .in0(N__46770),
            .in1(N__46727),
            .in2(_gnd_net_),
            .in3(N__46703),
            .lcout(\c0.n17180 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_4_lut_adj_688_LC_17_26_5 .C_ON=1'b0;
    defparam \c0.i2_3_lut_4_lut_adj_688_LC_17_26_5 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_4_lut_adj_688_LC_17_26_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i2_3_lut_4_lut_adj_688_LC_17_26_5  (
            .in0(N__47546),
            .in1(N__48826),
            .in2(N__47194),
            .in3(N__48728),
            .lcout(\c0.n17222 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_461_LC_17_27_1 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_461_LC_17_27_1 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_461_LC_17_27_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_461_LC_17_27_1  (
            .in0(N__46658),
            .in1(N__48570),
            .in2(N__46646),
            .in3(N__46589),
            .lcout(),
            .ltout(\c0.n10_adj_2191_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_4_lut_adj_462_LC_17_27_2 .C_ON=1'b0;
    defparam \c0.i1_4_lut_adj_462_LC_17_27_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_4_lut_adj_462_LC_17_27_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_4_lut_adj_462_LC_17_27_2  (
            .in0(N__46578),
            .in1(N__48884),
            .in2(N__46554),
            .in3(N__47331),
            .lcout(\c0.n17261 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i8_3_lut_LC_17_27_3 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i8_3_lut_LC_17_27_3 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i8_3_lut_LC_17_27_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_4_i8_3_lut_LC_17_27_3  (
            .in0(N__47048),
            .in1(N__48473),
            .in2(_gnd_net_),
            .in3(N__47840),
            .lcout(),
            .ltout(\c0.n8_adj_2198_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i10_4_lut_LC_17_27_4 .C_ON=1'b0;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i10_4_lut_LC_17_27_4 .SEQ_MODE=4'b0000;
    defparam \c0.byte_transmit_counter_4__I_0_Mux_4_i10_4_lut_LC_17_27_4 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \c0.byte_transmit_counter_4__I_0_Mux_4_i10_4_lut_LC_17_27_4  (
            .in0(N__47841),
            .in1(N__47547),
            .in2(N__47517),
            .in3(N__47514),
            .lcout(n10_adj_2430),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i2_3_lut_adj_457_LC_17_27_6 .C_ON=1'b0;
    defparam \c0.i2_3_lut_adj_457_LC_17_27_6 .SEQ_MODE=4'b0000;
    defparam \c0.i2_3_lut_adj_457_LC_17_27_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.i2_3_lut_adj_457_LC_17_27_6  (
            .in0(N__48791),
            .in1(N__47337),
            .in2(_gnd_net_),
            .in3(N__49865),
            .lcout(\c0.n17297 ),
            .ltout(\c0.n17297_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i5_3_lut_adj_436_LC_17_27_7 .C_ON=1'b0;
    defparam \c0.i5_3_lut_adj_436_LC_17_27_7 .SEQ_MODE=4'b0000;
    defparam \c0.i5_3_lut_adj_436_LC_17_27_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.i5_3_lut_adj_436_LC_17_27_7  (
            .in0(_gnd_net_),
            .in1(N__48532),
            .in2(N__47325),
            .in3(N__47320),
            .lcout(\c0.n14_adj_2176 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_10__0__2176_LC_17_28_1 .C_ON=1'b0;
    defparam \c0.data_out_10__0__2176_LC_17_28_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_10__0__2176_LC_17_28_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_10__0__2176_LC_17_28_1  (
            .in0(N__47163),
            .in1(N__47263),
            .in2(N__47211),
            .in3(N__46943),
            .lcout(data_out_10_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49842),
            .ce(N__49984),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_4_lut_adj_738_LC_17_28_3 .C_ON=1'b0;
    defparam \c0.i1_2_lut_4_lut_adj_738_LC_17_28_3 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_4_lut_adj_738_LC_17_28_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i1_2_lut_4_lut_adj_738_LC_17_28_3  (
            .in0(N__47162),
            .in1(N__47131),
            .in2(N__49161),
            .in3(N__49113),
            .lcout(\c0.n17162 ),
            .ltout(\c0.n17162_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_466_LC_17_28_4 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_466_LC_17_28_4 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_466_LC_17_28_4 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_466_LC_17_28_4  (
            .in0(N__47058),
            .in1(N__47049),
            .in2(N__47019),
            .in3(N__47013),
            .lcout(),
            .ltout(\c0.n10_adj_2196_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_10__1__2175_LC_17_28_5 .C_ON=1'b0;
    defparam \c0.data_out_10__1__2175_LC_17_28_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_10__1__2175_LC_17_28_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \c0.data_out_10__1__2175_LC_17_28_5  (
            .in0(_gnd_net_),
            .in1(N__46958),
            .in2(N__46947),
            .in3(N__46944),
            .lcout(data_out_10_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49842),
            .ce(N__49984),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_LC_17_29_0 .C_ON=1'b0;
    defparam \c0.i4_4_lut_LC_17_29_0 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_LC_17_29_0 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_LC_17_29_0  (
            .in0(N__48933),
            .in1(N__48903),
            .in2(N__48792),
            .in3(N__48885),
            .lcout(),
            .ltout(\c0.n10_adj_2166_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_9__1__2183_LC_17_29_1 .C_ON=1'b0;
    defparam \c0.data_out_9__1__2183_LC_17_29_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_9__1__2183_LC_17_29_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \c0.data_out_9__1__2183_LC_17_29_1  (
            .in0(N__48834),
            .in1(_gnd_net_),
            .in2(N__48795),
            .in3(N__48483),
            .lcout(\c0.data_out_9_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49847),
            .ce(N__49989),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_455_LC_17_29_2 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_455_LC_17_29_2 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_455_LC_17_29_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \c0.i1_2_lut_adj_455_LC_17_29_2  (
            .in0(N__48745),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48673),
            .lcout(\c0.n10170 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_10__5__2171_LC_17_29_3 .C_ON=1'b0;
    defparam \c0.data_out_10__5__2171_LC_17_29_3 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_10__5__2171_LC_17_29_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \c0.data_out_10__5__2171_LC_17_29_3  (
            .in0(N__48774),
            .in1(N__48746),
            .in2(_gnd_net_),
            .in3(N__48732),
            .lcout(\c0.data_out_10_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49847),
            .ce(N__49989),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_444_LC_17_29_4 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_444_LC_17_29_4 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_444_LC_17_29_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_444_LC_17_29_4  (
            .in0(_gnd_net_),
            .in1(N__48660),
            .in2(_gnd_net_),
            .in3(N__48621),
            .lcout(),
            .ltout(\c0.n17150_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_9__5__2179_LC_17_29_5 .C_ON=1'b0;
    defparam \c0.data_out_9__5__2179_LC_17_29_5 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_9__5__2179_LC_17_29_5 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.data_out_9__5__2179_LC_17_29_5  (
            .in0(N__48591),
            .in1(N__48582),
            .in2(N__48576),
            .in3(N__48566),
            .lcout(\c0.data_out_9_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49847),
            .ce(N__49989),
            .sr(_gnd_net_));
    defparam \c0.data_out_10__7__2169_LC_17_29_7 .C_ON=1'b0;
    defparam \c0.data_out_10__7__2169_LC_17_29_7 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_10__7__2169_LC_17_29_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.data_out_10__7__2169_LC_17_29_7  (
            .in0(_gnd_net_),
            .in1(N__48510),
            .in2(_gnd_net_),
            .in3(N__48482),
            .lcout(\c0.data_out_10_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49847),
            .ce(N__49989),
            .sr(_gnd_net_));
    defparam \c0.data_out_5__1__2215_LC_17_30_1 .C_ON=1'b0;
    defparam \c0.data_out_5__1__2215_LC_17_30_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_5__1__2215_LC_17_30_1 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \c0.data_out_5__1__2215_LC_17_30_1  (
            .in0(N__48412),
            .in1(N__48134),
            .in2(N__47901),
            .in3(N__50316),
            .lcout(data_out_5_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49850),
            .ce(N__50491),
            .sr(_gnd_net_));
    defparam \c0.tx.i1_2_lut_adj_403_LC_17_31_2 .C_ON=1'b0;
    defparam \c0.tx.i1_2_lut_adj_403_LC_17_31_2 .SEQ_MODE=4'b0000;
    defparam \c0.tx.i1_2_lut_adj_403_LC_17_31_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \c0.tx.i1_2_lut_adj_403_LC_17_31_2  (
            .in0(_gnd_net_),
            .in1(N__50816),
            .in2(_gnd_net_),
            .in3(N__50773),
            .lcout(n444),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_2__5__2235_LC_17_31_4 .C_ON=1'b0;
    defparam \c0.data_out_2__5__2235_LC_17_31_4 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_2__5__2235_LC_17_31_4 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \c0.data_out_2__5__2235_LC_17_31_4  (
            .in0(N__50411),
            .in1(N__50318),
            .in2(_gnd_net_),
            .in3(N__50003),
            .lcout(data_out_2_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49851),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.data_out_9__2__2182_LC_18_27_1 .C_ON=1'b0;
    defparam \c0.data_out_9__2__2182_LC_18_27_1 .SEQ_MODE=4'b1000;
    defparam \c0.data_out_9__2__2182_LC_18_27_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \c0.data_out_9__2__2182_LC_18_27_1  (
            .in0(N__49978),
            .in1(N__49151),
            .in2(_gnd_net_),
            .in3(N__49866),
            .lcout(data_out_9_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__49843),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i1_2_lut_adj_443_LC_18_28_1 .C_ON=1'b0;
    defparam \c0.i1_2_lut_adj_443_LC_18_28_1 .SEQ_MODE=4'b0000;
    defparam \c0.i1_2_lut_adj_443_LC_18_28_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \c0.i1_2_lut_adj_443_LC_18_28_1  (
            .in0(_gnd_net_),
            .in1(N__49147),
            .in2(_gnd_net_),
            .in3(N__49112),
            .lcout(),
            .ltout(\c0.n10204_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \c0.i4_4_lut_adj_426_LC_18_28_2 .C_ON=1'b0;
    defparam \c0.i4_4_lut_adj_426_LC_18_28_2 .SEQ_MODE=4'b0000;
    defparam \c0.i4_4_lut_adj_426_LC_18_28_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \c0.i4_4_lut_adj_426_LC_18_28_2  (
            .in0(N__49041),
            .in1(N__49013),
            .in2(N__48981),
            .in3(N__48978),
            .lcout(\c0.n10_adj_2172 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // TinyFPGA_B
